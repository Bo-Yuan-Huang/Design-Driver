
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire [15:0] _26874_;
  wire [7:0] _26875_;
  wire [7:0] _26876_;
  wire [7:0] _26877_;
  wire [7:0] _26878_;
  wire [7:0] _26879_;
  wire [7:0] _26880_;
  wire [7:0] _26881_;
  wire [7:0] _26882_;
  wire [7:0] _26883_;
  wire [7:0] _26884_;
  wire [7:0] _26885_;
  wire [7:0] _26886_;
  wire [7:0] _26887_;
  wire [7:0] _26888_;
  wire [7:0] _26889_;
  wire [7:0] _26890_;
  wire _26891_;
  wire [7:0] _26892_;
  wire [2:0] _26893_;
  wire [2:0] _26894_;
  wire [1:0] _26895_;
  wire [7:0] _26896_;
  wire _26897_;
  wire [1:0] _26898_;
  wire [1:0] _26899_;
  wire [2:0] _26900_;
  wire [2:0] _26901_;
  wire [1:0] _26902_;
  wire [3:0] _26903_;
  wire [1:0] _26904_;
  wire _26905_;
  wire [7:0] _26906_;
  wire [7:0] _26907_;
  wire [7:0] _26908_;
  wire [7:0] _26909_;
  wire [7:0] _26910_;
  wire [7:0] _26911_;
  wire [7:0] _26912_;
  wire [7:0] _26913_;
  wire [15:0] _26914_;
  wire [15:0] _26915_;
  wire _26916_;
  wire [4:0] _26917_;
  wire [7:0] _26918_;
  wire _26919_;
  wire _26920_;
  wire [15:0] _26921_;
  wire [15:0] _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire [7:0] _26926_;
  wire [2:0] _26927_;
  wire [7:0] _26928_;
  wire [7:0] _26929_;
  wire _26930_;
  wire [7:0] _26931_;
  wire _26932_;
  wire _26933_;
  wire [3:0] _26934_;
  wire [31:0] _26935_;
  wire [31:0] _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire [15:0] _26940_;
  wire _26941_;
  wire _26942_;
  wire [7:0] _26943_;
  wire _26944_;
  wire [2:0] _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire [7:0] _27326_;
  wire _27327_;
  wire [3:0] _27328_;
  wire _27329_;
  wire _27330_;
  wire [7:0] _27331_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  and (_22732_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_22733_, _22732_);
  not (_22734_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_22735_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_22736_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_22737_, _22736_, _22735_);
  nor (_22738_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_22739_, _22738_, _22734_);
  and (_22740_, _22739_, _22737_);
  not (_22741_, _22740_);
  not (_22742_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_22743_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_22744_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand (_22745_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_22746_, _22745_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_22747_, _22746_, _22744_);
  not (_22748_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_22749_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_22750_, _22749_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_22751_, _22750_, _22748_);
  not (_22752_, _22751_);
  nand (_22753_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_22754_, _22753_, _22747_);
  or (_22755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_22756_, _22755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_22757_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  not (_22758_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_22759_, _22755_, _22748_);
  or (_22760_, _22759_, _22758_);
  and (_22761_, _22760_, _22757_);
  nor (_22762_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_22763_, _22762_, _22748_);
  nand (_22764_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not (_22765_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_22766_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_22767_, _22766_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_22768_, _22767_, _22765_);
  and (_22769_, _22768_, _22764_);
  and (_22770_, _22769_, _22761_);
  nand (_22772_, _22770_, _22754_);
  nand (_22773_, _22772_, _22743_);
  nand (_22774_, _22773_, _22742_);
  nor (_22775_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _22742_);
  not (_22776_, _22775_);
  and (_22777_, _22776_, _22774_);
  or (_22778_, _22777_, _22741_);
  not (_22779_, _22737_);
  nor (_22780_, _22739_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_22781_, _22780_, _22779_);
  and (_22782_, _22781_, _22778_);
  not (_22783_, _22782_);
  nand (_22784_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  not (_22785_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_22786_, _22746_, _22785_);
  and (_22787_, _22786_, _22784_);
  not (_22788_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_22789_, _22767_, _22788_);
  nand (_22790_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_22791_, _22790_, _22789_);
  nand (_22793_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not (_22794_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_22796_, _22759_, _22794_);
  and (_22797_, _22796_, _22793_);
  and (_22798_, _22797_, _22791_);
  nand (_22799_, _22798_, _22787_);
  nand (_22800_, _22799_, _22743_);
  nand (_22801_, _22800_, _22742_);
  nor (_22802_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _22742_);
  not (_22803_, _22802_);
  and (_22804_, _22803_, _22801_);
  or (_22805_, _22804_, _22741_);
  nor (_22806_, _22739_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_22807_, _22806_, _22779_);
  nand (_22808_, _22807_, _22805_);
  and (_22809_, _22808_, _22783_);
  nand (_22810_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not (_22811_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_22812_, _22767_, _22811_);
  and (_22813_, _22812_, _22810_);
  nand (_22814_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  not (_22815_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_22816_, _22759_, _22815_);
  and (_22817_, _22816_, _22814_);
  nand (_22818_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_22819_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_22820_, _22746_, _22819_);
  and (_22821_, _22820_, _22818_);
  and (_22822_, _22821_, _22817_);
  and (_22823_, _22822_, _22813_);
  or (_22824_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_22825_, _22824_, _22823_);
  and (_22827_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not (_22828_, _22827_);
  and (_22830_, _22828_, _22825_);
  nand (_22831_, _22830_, _22740_);
  nor (_22832_, _22739_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_22833_, _22832_, _22779_);
  and (_22835_, _22833_, _22831_);
  not (_22836_, _22835_);
  not (_22837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_22838_, _22759_, _22837_);
  not (_22839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_22840_, _22746_, _22839_);
  and (_22841_, _22840_, _22838_);
  not (_22842_, _22767_);
  and (_22843_, _22842_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_22844_, _22843_);
  and (_22845_, _22844_, _22841_);
  nand (_22846_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_22847_, _22846_, _22743_);
  nand (_22848_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_22849_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_22850_, _22849_, _22848_);
  and (_22851_, _22850_, _22847_);
  and (_22852_, _22851_, _22845_);
  and (_22853_, _22852_, _22742_);
  nor (_22854_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _22742_);
  or (_22855_, _22854_, _22853_);
  and (_22856_, _22855_, _22740_);
  not (_22857_, _22856_);
  nor (_22858_, _22739_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_22859_, _22858_, _22779_);
  nand (_22860_, _22859_, _22857_);
  and (_22861_, _22860_, _22836_);
  and (_22862_, _22861_, _22809_);
  nor (_22863_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_22864_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_22865_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_22866_, _22865_, _22864_);
  not (_22868_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_22869_, _22746_, _22868_);
  not (_22871_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_22872_, _22767_, _22871_);
  and (_22873_, _22872_, _22869_);
  nand (_22874_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_22875_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_22876_, _22759_, _22875_);
  and (_22877_, _22876_, _22874_);
  and (_22878_, _22877_, _22873_);
  nand (_22879_, _22878_, _22866_);
  nand (_22880_, _22879_, _22863_);
  and (_22881_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_22882_, _22881_);
  and (_22883_, _22882_, _22880_);
  nand (_22885_, _22883_, _22740_);
  nor (_22886_, _22739_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_22888_, _22886_, _22779_);
  and (_22889_, _22888_, _22885_);
  nand (_22891_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_22892_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_22894_, _22892_, _22891_);
  not (_22895_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_22896_, _22746_, _22895_);
  not (_22897_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_22898_, _22767_, _22897_);
  and (_22899_, _22898_, _22896_);
  nand (_22900_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not (_22901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_22902_, _22759_, _22901_);
  and (_22903_, _22902_, _22900_);
  and (_22904_, _22903_, _22899_);
  and (_22905_, _22904_, _22894_);
  or (_22906_, _22905_, _22824_);
  and (_22907_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_22908_, _22907_);
  nand (_22909_, _22908_, _22906_);
  or (_22910_, _22909_, _22741_);
  nor (_22911_, _22739_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_22912_, _22911_, _22779_);
  and (_22913_, _22912_, _22910_);
  not (_22914_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_22915_, _22759_, _22914_);
  not (_22916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_22917_, _22751_, _22916_);
  and (_22918_, _22917_, _22915_);
  not (_22919_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_22920_, _22746_, _22919_);
  not (_22921_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_22922_, _22767_, _22921_);
  and (_22923_, _22922_, _22920_);
  and (_22924_, _22923_, _22918_);
  nand (_22925_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_22926_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_22927_, _22926_, _22925_);
  and (_22928_, _22927_, _22924_);
  or (_22929_, _22928_, _22824_);
  and (_22931_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_22932_, _22931_);
  nand (_22934_, _22932_, _22929_);
  or (_22935_, _22934_, _22741_);
  nor (_22936_, _22739_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_22937_, _22936_, _22779_);
  nand (_22938_, _22937_, _22935_);
  nor (_22939_, _22938_, _22913_);
  and (_22940_, _22939_, _22889_);
  not (_22942_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_22943_, \oc8051_top_1.oc8051_decoder1.state [1], _22734_);
  and (_22944_, _22943_, _22942_);
  and (_22945_, _22944_, _22940_);
  and (_22946_, _22945_, _22862_);
  not (_22947_, _22860_);
  and (_22948_, _22947_, _22809_);
  and (_22949_, _22948_, _22835_);
  and (_22950_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_22951_, _22746_);
  and (_22952_, _22951_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_22953_, _22842_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_22954_, _22953_, _22952_);
  or (_22956_, _22954_, _22950_);
  and (_22957_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_22958_, _22957_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_22959_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  not (_22960_, _22759_);
  and (_22961_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_22962_, _22961_, _22959_);
  or (_22963_, _22962_, _22958_);
  or (_22964_, _22963_, _22956_);
  or (_22965_, _22964_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_22966_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _22742_);
  not (_22967_, _22966_);
  and (_22968_, _22967_, _22965_);
  or (_22969_, _22968_, _22741_);
  nor (_22970_, _22739_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_22971_, _22970_, _22779_);
  and (_22972_, _22971_, _22969_);
  not (_22973_, _22972_);
  and (_22974_, _22938_, _22913_);
  and (_22975_, _22974_, _22889_);
  and (_22976_, _22975_, _22973_);
  and (_22977_, _22976_, _22949_);
  not (_22979_, _22977_);
  not (_22980_, _22889_);
  and (_22981_, _22972_, _22980_);
  and (_22982_, _22981_, _22974_);
  and (_22983_, _22982_, _22949_);
  and (_22984_, _22972_, _22940_);
  and (_22985_, _22984_, _22949_);
  nor (_22986_, _22985_, _22983_);
  and (_22987_, _22986_, _22979_);
  nor (_22988_, _22860_, _22783_);
  and (_22989_, _22988_, _22808_);
  not (_22990_, _22913_);
  and (_22991_, _22938_, _22990_);
  and (_22992_, _22991_, _22889_);
  and (_22993_, _22939_, _22980_);
  and (_22994_, _22993_, _22972_);
  or (_22995_, _22994_, _22992_);
  and (_22996_, _22995_, _22989_);
  and (_22997_, _22991_, _22980_);
  and (_22998_, _22997_, _22989_);
  and (_22999_, _22972_, _22808_);
  and (_23000_, _22999_, _22988_);
  and (_23001_, _23000_, _22975_);
  nor (_23002_, _23001_, _22998_);
  not (_23004_, _23002_);
  nor (_23005_, _23004_, _22996_);
  not (_23006_, _22938_);
  and (_23007_, _23006_, _22889_);
  and (_23008_, _23007_, _22913_);
  and (_23009_, _23008_, _22973_);
  and (_23010_, _22993_, _22973_);
  or (_23011_, _23010_, _23009_);
  and (_23012_, _23011_, _22989_);
  not (_23013_, _23012_);
  and (_23015_, _23013_, _23005_);
  nor (_23016_, _22938_, _22889_);
  and (_23017_, _23016_, _22913_);
  and (_23018_, _23017_, _22972_);
  and (_23019_, _23018_, _22862_);
  and (_23021_, _23017_, _22989_);
  and (_23022_, _22974_, _22980_);
  and (_23023_, _23000_, _23022_);
  nor (_23024_, _23023_, _23021_);
  not (_23025_, _23024_);
  nor (_23026_, _23025_, _23019_);
  and (_23027_, _22948_, _22836_);
  and (_23028_, _23027_, _22992_);
  not (_23029_, _23028_);
  and (_23030_, _23022_, _22973_);
  and (_23031_, _23030_, _22989_);
  and (_23032_, _22973_, _22940_);
  and (_23034_, _23032_, _22989_);
  nor (_23035_, _23034_, _23031_);
  and (_23036_, _23035_, _23029_);
  and (_23037_, _23036_, _23026_);
  and (_23038_, _23037_, _23015_);
  and (_23039_, _23038_, _22987_);
  or (_23040_, _22738_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23041_, \oc8051_top_1.oc8051_decoder1.state [0], _22734_);
  and (_23042_, _23041_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_23043_, _23042_, _23028_);
  nor (_23044_, _23043_, _23040_);
  nor (_23045_, _23044_, _23039_);
  or (_23046_, _23045_, _22946_);
  nand (_23047_, _23046_, _22734_);
  and (_23048_, _23047_, _22733_);
  not (_23049_, rst);
  and (_23050_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23051_, _22808_, _22782_);
  and (_23052_, _23051_, _22861_);
  and (_23053_, _23052_, _23030_);
  and (_23054_, _23052_, _22976_);
  nor (_23055_, _23054_, _23053_);
  and (_23056_, _22939_, _22862_);
  and (_23057_, _23056_, _22944_);
  not (_23058_, _23057_);
  and (_23059_, _23058_, _23055_);
  not (_23061_, _23040_);
  or (_23062_, _23061_, _22987_);
  and (_23063_, _23062_, _23059_);
  nor (_23064_, _23063_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_23065_, _23064_, _23050_);
  nand (_23066_, _23065_, _23049_);
  nor (_26941_, _23066_, _23048_);
  and (_23067_, \oc8051_top_1.oc8051_decoder1.wr , _22734_);
  not (_23068_, _23067_);
  not (_23069_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23070_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22734_);
  and (_23071_, _23070_, _23069_);
  and (_23072_, _23071_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23074_, _23073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_23075_, _23074_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_23076_, _23075_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_23077_, _23076_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_23078_, _23077_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_23079_, _23078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_23080_, _23078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_23081_, _23080_, _23079_);
  and (_23082_, _23081_, _23072_);
  not (_23083_, _23082_);
  and (_23084_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23085_, _23084_, _23070_);
  nor (_23086_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23087_, _23086_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23088_, _23087_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23089_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_23090_, _23089_, _23085_);
  and (_23091_, _23087_, _23069_);
  and (_23092_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_23093_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23094_, _23093_, _23070_);
  and (_23095_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor (_23096_, _23095_, _23092_);
  and (_23097_, _23096_, _23090_);
  and (_23098_, _23097_, _23083_);
  nor (_23099_, _23098_, _23071_);
  nor (_23100_, _23099_, _23068_);
  not (_23101_, _23100_);
  and (_23102_, _23098_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23103_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  not (_23104_, _23103_);
  and (_23105_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_23106_, _23105_, _23085_);
  and (_23108_, _23106_, _23104_);
  nor (_23109_, _23075_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_23110_, _23109_);
  not (_23111_, _23072_);
  nor (_23112_, _23111_, _23076_);
  and (_23113_, _23112_, _23110_);
  nor (_23114_, _23093_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_23115_, _23114_, _23070_);
  not (_23116_, _23115_);
  and (_23117_, _23116_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_23118_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_23119_, _23118_, _23117_);
  not (_23120_, _23119_);
  nor (_23121_, _23120_, _23113_);
  and (_23122_, _23121_, _23108_);
  not (_23123_, _23122_);
  and (_23124_, _23123_, _23102_);
  nor (_23125_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_23126_, _23125_, _23073_);
  and (_23127_, _23126_, _23072_);
  and (_23129_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_23130_, _23129_, _23127_);
  and (_23131_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_23132_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_23133_, _23116_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_23134_, _23133_, _23132_);
  nor (_23136_, _23134_, _23131_);
  and (_23137_, _23136_, _23130_);
  nor (_23138_, _23137_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23139_, _23138_, _23124_);
  nor (_23140_, _23139_, _23101_);
  nor (_23142_, _23074_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_23143_, _23142_, _23075_);
  and (_23144_, _23143_, _23072_);
  not (_23145_, _23144_);
  and (_23146_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_23147_, _23116_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_23148_, _23147_, _23146_);
  and (_23149_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_23150_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_23151_, _23150_, _23149_);
  and (_23152_, _23151_, _23148_);
  and (_23153_, _23152_, _23145_);
  not (_23154_, _23153_);
  and (_23155_, _23154_, _23102_);
  and (_23156_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_23157_, _23116_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_23158_, _23157_, _23156_);
  not (_23159_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23160_, _23072_, _23159_);
  not (_23161_, _23160_);
  and (_23162_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_23163_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_23165_, _23163_, _23162_);
  and (_23166_, _23165_, _23161_);
  and (_23167_, _23166_, _23158_);
  nor (_23168_, _23167_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23169_, _23168_, _23155_);
  and (_23170_, _23169_, _23140_);
  nor (_23171_, _23077_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_23173_, _23171_);
  nor (_23174_, _23111_, _23078_);
  and (_23175_, _23174_, _23173_);
  not (_23176_, _23175_);
  and (_23177_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_23178_, _23177_, _23085_);
  and (_23179_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23180_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor (_23181_, _23180_, _23179_);
  and (_23182_, _23181_, _23178_);
  and (_23183_, _23182_, _23176_);
  not (_23184_, _23183_);
  and (_23185_, _23184_, _23102_);
  nor (_23186_, _23153_, _23102_);
  nor (_23187_, _23186_, _23185_);
  nor (_23189_, _23187_, _23101_);
  nor (_23190_, _23076_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_23191_, _23190_);
  nor (_23192_, _23111_, _23077_);
  and (_23193_, _23192_, _23191_);
  not (_23194_, _23193_);
  and (_23195_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_23196_, _23195_, _23085_);
  and (_23197_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_23198_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_23199_, _23198_, _23197_);
  and (_23200_, _23199_, _23196_);
  and (_23201_, _23200_, _23194_);
  not (_23202_, _23201_);
  and (_23203_, _23202_, _23102_);
  nor (_23204_, _23073_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_23205_, _23204_, _23074_);
  and (_23207_, _23205_, _23072_);
  and (_23208_, _23094_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_23209_, _23208_, _23207_);
  and (_23210_, _23088_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_23211_, _23091_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_23212_, _23116_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_23213_, _23212_, _23211_);
  nor (_23214_, _23213_, _23210_);
  and (_23215_, _23214_, _23209_);
  nor (_23216_, _23215_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23217_, _23216_, _23203_);
  nor (_23218_, _23217_, _23101_);
  and (_23219_, _23218_, _23189_);
  and (_23220_, _23219_, _23170_);
  nor (_23221_, _23122_, _23102_);
  and (_23222_, _23221_, _23100_);
  and (_23223_, _23222_, _23201_);
  nor (_23224_, _23183_, _23102_);
  and (_23225_, _23224_, _23100_);
  not (_23226_, _23098_);
  and (_23227_, _23100_, _23226_);
  nor (_23229_, _23227_, _23225_);
  and (_23230_, _23229_, _23223_);
  and (_23231_, _23230_, _23220_);
  and (_23232_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22734_);
  and (_23233_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22734_);
  nor (_23234_, _23233_, _23232_);
  not (_23235_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_23236_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _22734_);
  and (_23237_, _23236_, _23235_);
  and (_23238_, _23237_, _23234_);
  not (_23239_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_23240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_23242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23243_, _23242_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_23244_, _23243_, _23240_);
  or (_23245_, _23244_, _23239_);
  nor (_23246_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_23247_, _23246_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23248_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_23249_, _23248_, _23245_);
  not (_23250_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_23251_, _23243_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23252_, _23251_, _23250_);
  not (_23253_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_23255_, _23240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23256_, _23255_, _23242_);
  or (_23257_, _23256_, _23253_);
  and (_23258_, _23257_, _23252_);
  and (_23259_, _23258_, _23249_);
  nand (_23260_, _23246_, _23240_);
  or (_23261_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_23262_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23263_, _23262_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23264_, _23263_, _23261_);
  not (_23265_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_23266_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23265_);
  or (_23267_, _23266_, _23264_);
  nand (_23268_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _23265_);
  or (_23269_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23270_, _23269_, _23267_);
  or (_23271_, _23270_, _23260_);
  and (_23272_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_23273_, _23272_, _23240_);
  nand (_23274_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_23275_, _23272_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23276_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_23277_, _23276_, _23274_);
  and (_23278_, _23277_, _23271_);
  and (_23279_, _23278_, _23259_);
  or (_23280_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23281_, _23280_, _23270_);
  and (_23282_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_23283_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23284_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_23285_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23286_, _23285_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor (_23287_, _23286_, _23284_);
  nor (_23288_, _23287_, _23283_);
  and (_23289_, _23288_, _23281_);
  nor (_23290_, _23289_, _23279_);
  not (_23291_, _23290_);
  not (_23292_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23293_, _23251_, _23292_);
  not (_23294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or (_23295_, _23256_, _23294_);
  and (_23296_, _23295_, _23293_);
  nand (_23297_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_23298_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23299_, _23244_, _23298_);
  and (_23300_, _23299_, _23297_);
  and (_23302_, _23300_, _23296_);
  or (_23303_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_23304_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23262_);
  and (_23305_, _23304_, _23303_);
  or (_23306_, _23305_, _23266_);
  or (_23307_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23308_, _23307_, _23306_);
  or (_23309_, _23308_, _23260_);
  nand (_23311_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand (_23312_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_23313_, _23312_, _23311_);
  and (_23315_, _23313_, _23309_);
  nand (_23316_, _23315_, _23302_);
  or (_23317_, _23308_, _23280_);
  nand (_23318_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_23319_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_23320_, _23286_, _23319_);
  and (_23321_, _23320_, _23318_);
  nand (_23322_, _23321_, _23317_);
  and (_23323_, _23322_, _23316_);
  nor (_23324_, _23322_, _23316_);
  nor (_23325_, _23324_, _23323_);
  not (_23326_, _23244_);
  nand (_23327_, _23326_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_23328_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_23329_, _23328_, _23327_);
  not (_23331_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or (_23332_, _23256_, _23331_);
  not (_23333_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23334_, _23251_, _23333_);
  and (_23335_, _23334_, _23332_);
  and (_23336_, _23335_, _23329_);
  or (_23337_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_23338_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23262_);
  and (_23339_, _23338_, _23337_);
  or (_23340_, _23339_, _23266_);
  or (_23341_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_23342_, _23341_, _23340_);
  or (_23343_, _23342_, _23260_);
  nand (_23344_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nand (_23345_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_23346_, _23345_, _23344_);
  and (_23347_, _23346_, _23343_);
  and (_23348_, _23347_, _23336_);
  or (_23349_, _23342_, _23280_);
  nand (_23350_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_23351_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_23352_, _23286_, _23351_);
  and (_23353_, _23352_, _23350_);
  and (_23354_, _23353_, _23349_);
  nor (_23355_, _23354_, _23348_);
  and (_23356_, _23354_, _23348_);
  nor (_23357_, _23356_, _23355_);
  nand (_23358_, _23326_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_23359_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_23360_, _23359_, _23358_);
  not (_23361_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23362_, _23251_, _23361_);
  not (_23363_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_23364_, _23256_, _23363_);
  and (_23365_, _23364_, _23362_);
  and (_23366_, _23365_, _23360_);
  or (_23367_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_23368_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23262_);
  and (_23369_, _23368_, _23367_);
  or (_23370_, _23369_, _23266_);
  or (_23371_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_23372_, _23371_, _23370_);
  or (_23373_, _23372_, _23260_);
  nand (_23374_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nand (_23375_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_23376_, _23375_, _23374_);
  and (_23377_, _23376_, _23373_);
  and (_23378_, _23377_, _23366_);
  or (_23379_, _23372_, _23280_);
  nand (_23380_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_23381_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_23382_, _23286_, _23381_);
  and (_23383_, _23382_, _23380_);
  and (_23384_, _23383_, _23379_);
  nor (_23385_, _23384_, _23378_);
  and (_23386_, _23384_, _23378_);
  nor (_23387_, _23386_, _23385_);
  nand (_23388_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_23389_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_23390_, _23389_, _23388_);
  not (_23391_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23392_, _23244_, _23391_);
  nand (_23393_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_23394_, _23393_, _23392_);
  and (_23395_, _23394_, _23390_);
  or (_23397_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_23398_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23262_);
  and (_23400_, _23398_, _23397_);
  or (_23401_, _23400_, _23266_);
  or (_23402_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_23403_, _23402_, _23401_);
  or (_23404_, _23403_, _23260_);
  not (_23405_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23406_, _23251_, _23405_);
  not (_23407_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or (_23408_, _23256_, _23407_);
  and (_23410_, _23408_, _23406_);
  and (_23411_, _23410_, _23404_);
  nand (_23412_, _23411_, _23395_);
  or (_23414_, _23403_, _23280_);
  nand (_23415_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_23416_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_23417_, _23286_, _23416_);
  and (_23418_, _23417_, _23415_);
  nand (_23419_, _23418_, _23414_);
  and (_23420_, _23419_, _23412_);
  nor (_23421_, _23419_, _23412_);
  nor (_23422_, _23421_, _23420_);
  not (_23423_, _23422_);
  not (_23424_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_23425_, _23244_, _23424_);
  nand (_23426_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_23427_, _23426_, _23425_);
  not (_23428_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_23429_, _23256_, _23428_);
  not (_23430_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23432_, _23251_, _23430_);
  and (_23433_, _23432_, _23429_);
  and (_23435_, _23433_, _23427_);
  or (_23436_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_23437_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23262_);
  and (_23438_, _23437_, _23436_);
  or (_23439_, _23438_, _23266_);
  or (_23440_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_23441_, _23440_, _23439_);
  or (_23443_, _23441_, _23260_);
  nand (_23444_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand (_23445_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_23446_, _23445_, _23444_);
  and (_23447_, _23446_, _23443_);
  nand (_23448_, _23447_, _23435_);
  or (_23449_, _23441_, _23280_);
  nand (_23450_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_23451_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_23452_, _23286_, _23451_);
  and (_23453_, _23452_, _23450_);
  nand (_23454_, _23453_, _23449_);
  and (_23455_, _23454_, _23448_);
  and (_23456_, _23326_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_23457_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_23458_, _23457_, _23456_);
  not (_23459_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_23460_, _23256_, _23459_);
  not (_23461_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_23462_, _23251_, _23461_);
  nor (_23463_, _23462_, _23460_);
  and (_23464_, _23463_, _23458_);
  or (_23465_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_23466_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23262_);
  and (_23467_, _23466_, _23465_);
  or (_23468_, _23467_, _23266_);
  or (_23469_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_23470_, _23469_, _23468_);
  or (_23471_, _23470_, _23260_);
  and (_23472_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_23473_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_23474_, _23473_, _23472_);
  and (_23475_, _23474_, _23471_);
  and (_23476_, _23475_, _23464_);
  or (_23478_, _23470_, _23280_);
  nand (_23479_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_23480_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_23481_, _23286_, _23480_);
  and (_23482_, _23481_, _23479_);
  nand (_23483_, _23482_, _23478_);
  not (_23484_, _23483_);
  nor (_23485_, _23484_, _23476_);
  nor (_23486_, _23454_, _23448_);
  nor (_23487_, _23486_, _23455_);
  and (_23488_, _23487_, _23485_);
  nor (_23489_, _23488_, _23455_);
  nor (_23490_, _23489_, _23423_);
  nor (_23491_, _23490_, _23420_);
  nor (_23492_, _23491_, _23387_);
  and (_23493_, _23491_, _23387_);
  nor (_23494_, _23493_, _23492_);
  not (_23495_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or (_23496_, _23305_, _23495_);
  not (_23497_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23498_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _23497_);
  or (_23499_, _23438_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_23500_, _23499_, _23498_);
  nand (_23501_, _23500_, _23496_);
  not (_23502_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_23503_, _23502_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  or (_23504_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_23505_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23262_);
  and (_23506_, _23505_, _23504_);
  nand (_23507_, _23506_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23509_, _23400_, _23495_);
  nand (_23510_, _23509_, _23507_);
  nand (_23511_, _23510_, _23503_);
  and (_23512_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23513_, _23512_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23514_, _23513_, _23264_);
  nor (_23515_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23516_, _23515_, _23495_);
  nand (_23517_, _23516_, _23467_);
  and (_23518_, _23517_, _23514_);
  and (_23519_, _23512_, _23495_);
  nand (_23520_, _23519_, _23369_);
  and (_23521_, _23515_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23522_, _23521_, _23339_);
  and (_23523_, _23522_, _23520_);
  and (_23524_, _23523_, _23518_);
  and (_23525_, _23524_, _23511_);
  nand (_23526_, _23525_, _23501_);
  nand (_23527_, _23526_, _23268_);
  and (_23528_, _23266_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_23529_, _23528_);
  and (_23530_, _23529_, _23527_);
  and (_23531_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_23532_, _23531_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor (_23533_, _23532_, _23530_);
  not (_23534_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23535_, _23532_, _23534_);
  nor (_23536_, _23535_, _23533_);
  and (_23538_, _23484_, _23476_);
  nor (_23539_, _23538_, _23485_);
  not (_23540_, _23539_);
  nor (_23541_, _23540_, _23536_);
  and (_23542_, _23541_, _23487_);
  and (_23543_, _23489_, _23423_);
  nor (_23544_, _23543_, _23490_);
  and (_23545_, _23544_, _23542_);
  not (_23546_, _23545_);
  nor (_23547_, _23546_, _23494_);
  nor (_23548_, _23491_, _23386_);
  or (_23549_, _23548_, _23385_);
  or (_23550_, _23549_, _23547_);
  and (_23551_, _23550_, _23357_);
  and (_23552_, _23551_, _23325_);
  not (_23553_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23554_, _23251_, _23553_);
  not (_23555_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_23556_, _23256_, _23555_);
  and (_23557_, _23556_, _23554_);
  nand (_23558_, _23247_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_23559_, _23326_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_23560_, _23559_, _23558_);
  and (_23561_, _23560_, _23557_);
  or (_23562_, _23506_, _23266_);
  or (_23563_, _23268_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_23564_, _23563_, _23562_);
  or (_23565_, _23564_, _23260_);
  nand (_23566_, _23275_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nand (_23567_, _23273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_23568_, _23567_, _23566_);
  and (_23569_, _23568_, _23565_);
  and (_23570_, _23569_, _23561_);
  or (_23571_, _23564_, _23280_);
  nand (_23572_, _23282_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_23573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_23574_, _23286_, _23573_);
  and (_23575_, _23574_, _23572_);
  nand (_23576_, _23575_, _23571_);
  not (_23577_, _23576_);
  nor (_23578_, _23577_, _23570_);
  and (_23579_, _23577_, _23570_);
  nor (_23580_, _23579_, _23578_);
  not (_23581_, _23580_);
  and (_23582_, _23355_, _23325_);
  nor (_23583_, _23582_, _23323_);
  nor (_23584_, _23583_, _23581_);
  and (_23585_, _23583_, _23581_);
  nor (_23586_, _23585_, _23584_);
  and (_23587_, _23586_, _23552_);
  nor (_23588_, _23584_, _23578_);
  not (_23589_, _23588_);
  nor (_23590_, _23589_, _23587_);
  and (_23591_, _23289_, _23279_);
  or (_23592_, _23591_, _23590_);
  nand (_23594_, _23592_, _23291_);
  and (_23595_, _23594_, _23238_);
  not (_23597_, _23595_);
  not (_23598_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23599_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22734_);
  and (_23600_, _23599_, _23598_);
  and (_23601_, _23600_, _23234_);
  not (_23602_, _23601_);
  not (_23603_, _23289_);
  and (_23604_, _23603_, _23279_);
  nor (_23605_, _23591_, _23290_);
  nor (_23606_, _23576_, _23570_);
  and (_23607_, _23321_, _23317_);
  and (_23608_, _23607_, _23316_);
  nand (_23609_, _23353_, _23349_);
  and (_23610_, _23609_, _23348_);
  nor (_23611_, _23610_, _23325_);
  nor (_23612_, _23611_, _23608_);
  nor (_23613_, _23612_, _23580_);
  nor (_23614_, _23613_, _23606_);
  and (_23615_, _23612_, _23580_);
  nor (_23616_, _23615_, _23613_);
  not (_23617_, _23616_);
  and (_23618_, _23610_, _23325_);
  nor (_23619_, _23618_, _23611_);
  not (_23620_, _23619_);
  not (_23621_, _23357_);
  and (_23622_, _23483_, _23476_);
  nor (_23623_, _23622_, _23487_);
  not (_23624_, _23454_);
  and (_23625_, _23624_, _23448_);
  nor (_23626_, _23625_, _23623_);
  nor (_23627_, _23626_, _23422_);
  and (_23628_, _23418_, _23414_);
  and (_23629_, _23628_, _23412_);
  nor (_23630_, _23629_, _23627_);
  nor (_23631_, _23630_, _23387_);
  and (_23632_, _23630_, _23387_);
  nor (_23633_, _23632_, _23631_);
  and (_23634_, _23626_, _23422_);
  nor (_23635_, _23634_, _23627_);
  not (_23636_, _23635_);
  and (_23637_, _23622_, _23487_);
  nor (_23639_, _23637_, _23623_);
  not (_23640_, _23639_);
  nor (_23642_, _23539_, _23536_);
  and (_23643_, _23642_, _23640_);
  and (_23644_, _23643_, _23636_);
  not (_23645_, _23644_);
  nor (_23646_, _23645_, _23633_);
  nand (_23647_, _23383_, _23379_);
  or (_23648_, _23647_, _23378_);
  and (_23649_, _23647_, _23378_);
  or (_23650_, _23630_, _23649_);
  and (_23651_, _23650_, _23648_);
  or (_23652_, _23651_, _23646_);
  and (_23653_, _23652_, _23621_);
  and (_23654_, _23653_, _23620_);
  and (_23655_, _23654_, _23617_);
  nor (_23656_, _23655_, _23614_);
  nor (_23657_, _23656_, _23605_);
  nor (_23659_, _23657_, _23604_);
  nor (_23660_, _23659_, _23602_);
  not (_23661_, _23348_);
  not (_23662_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23663_, _23233_, _23662_);
  and (_23664_, _23663_, _23237_);
  nor (_23665_, _23448_, _23412_);
  nor (_23666_, _23665_, _23378_);
  and (_23667_, _23666_, _23664_);
  and (_23668_, _23667_, _23661_);
  not (_23669_, _23316_);
  and (_23670_, _23570_, _23669_);
  not (_23671_, _23670_);
  nor (_23672_, _23671_, _23668_);
  not (_23673_, _23672_);
  nor (_23674_, _23536_, _23279_);
  and (_23675_, _23674_, _23673_);
  nor (_23676_, _23668_, _23316_);
  and (_23677_, _23570_, _23536_);
  and (_23678_, _23677_, _23676_);
  not (_23679_, _23664_);
  and (_23680_, _23536_, _23279_);
  or (_23681_, _23680_, _23679_);
  or (_23682_, _23681_, _23678_);
  nor (_23683_, _23682_, _23675_);
  not (_23684_, _23683_);
  not (_23685_, _23530_);
  and (_23686_, _23532_, _23685_);
  not (_23687_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23688_, _23232_, _23687_);
  and (_23689_, _23688_, _23600_);
  and (_23690_, _23599_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23691_, _23690_, _23663_);
  and (_23692_, _23691_, _23685_);
  nor (_23693_, _23692_, _23689_);
  nor (_23694_, _23693_, _23686_);
  nor (_23695_, _23599_, _23236_);
  and (_23696_, _23232_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23697_, _23696_, _23695_);
  and (_23698_, _23697_, _23535_);
  and (_23699_, _23698_, _23530_);
  and (_23700_, _23663_, _23600_);
  and (_23701_, _23700_, _23536_);
  or (_23702_, _23701_, _23699_);
  nor (_23703_, _23535_, _23685_);
  and (_23704_, _23688_, _23237_);
  and (_23705_, _23695_, _23688_);
  not (_23706_, _23705_);
  nor (_23707_, _23706_, _23533_);
  nor (_23708_, _23707_, _23704_);
  nor (_23709_, _23708_, _23703_);
  not (_23710_, _23536_);
  and (_23711_, _23695_, _23234_);
  and (_23712_, _23711_, _23710_);
  not (_23713_, _23712_);
  not (_23714_, _23279_);
  and (_23715_, _23690_, _23688_);
  and (_23716_, _23715_, _23714_);
  not (_23717_, _23476_);
  and (_23718_, _23696_, _23237_);
  and (_23719_, _23718_, _23717_);
  or (_23720_, _23719_, _23667_);
  nor (_23721_, _23720_, _23716_);
  nand (_23722_, _23721_, _23713_);
  or (_23723_, _23722_, _23709_);
  or (_23724_, _23723_, _23702_);
  nor (_23725_, _23724_, _23694_);
  and (_23726_, _23725_, _23684_);
  not (_23727_, _23726_);
  nor (_23728_, _23727_, _23660_);
  and (_23729_, _23728_, _23597_);
  not (_23730_, _23729_);
  and (_23731_, _23495_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23732_, _23731_, _23515_);
  and (_23733_, _23732_, _23730_);
  and (_23734_, _23705_, _23539_);
  and (_23735_, _23691_, _23485_);
  not (_23736_, _23704_);
  nor (_23737_, _23736_, _23538_);
  and (_23738_, _23700_, _23476_);
  or (_23739_, _23738_, _23737_);
  or (_23740_, _23739_, _23735_);
  nor (_23741_, _23740_, _23734_);
  and (_23742_, _23696_, _23690_);
  and (_23743_, _23742_, _23483_);
  and (_23744_, _23696_, _23600_);
  and (_23745_, _23744_, _23476_);
  nor (_23746_, _23745_, _23743_);
  and (_23747_, _23688_, _23599_);
  not (_23748_, _23747_);
  and (_23749_, _23236_, _23234_);
  nor (_23750_, _23664_, _23749_);
  and (_23751_, _23750_, _23748_);
  and (_23752_, _23695_, _23663_);
  nor (_23753_, _23752_, _23697_);
  and (_23754_, _23753_, _23751_);
  nor (_23755_, _23754_, _23476_);
  not (_23756_, _23755_);
  and (_23757_, _23711_, _23717_);
  nor (_23758_, _23757_, _23719_);
  and (_23759_, _23758_, _23756_);
  and (_23760_, _23759_, _23746_);
  and (_23761_, _23760_, _23741_);
  nor (_23762_, _23761_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_23763_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23764_, _23732_, _23763_);
  and (_23765_, _23764_, _23467_);
  or (_23766_, _23765_, _23762_);
  or (_23767_, _23766_, _23733_);
  and (_23768_, _23767_, _23100_);
  and (_23769_, _23768_, _23231_);
  not (_23770_, _23231_);
  and (_23771_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_00877_, _23771_, _23769_);
  nor (_23772_, _23169_, _23101_);
  and (_23773_, _23772_, _23140_);
  nor (_23774_, _23218_, _23189_);
  and (_23775_, _23774_, _23773_);
  and (_23776_, _23222_, _23202_);
  nor (_23777_, _23184_, _23098_);
  and (_23779_, _23777_, _23776_);
  and (_23780_, _23779_, _23775_);
  not (_23782_, _23780_);
  and (_23783_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_23784_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23786_, _23784_, _23515_);
  nor (_23787_, _23786_, _23729_);
  and (_23788_, _23536_, _23661_);
  nor (_23789_, _23536_, _23354_);
  or (_23790_, _23789_, _23788_);
  and (_23791_, _23790_, _23742_);
  and (_23792_, _23665_, _23476_);
  and (_23793_, _23792_, _23378_);
  or (_23794_, _23793_, _23536_);
  not (_23795_, _23378_);
  and (_23796_, _23717_, _23448_);
  and (_23797_, _23796_, _23412_);
  and (_23798_, _23797_, _23795_);
  or (_23799_, _23798_, _23710_);
  and (_23800_, _23799_, _23794_);
  or (_23801_, _23800_, _23661_);
  nand (_23802_, _23800_, _23661_);
  and (_23803_, _23802_, _23801_);
  and (_23804_, _23803_, _23744_);
  nor (_23805_, _23804_, _23791_);
  nor (_23806_, _23711_, _23749_);
  and (_23807_, _23696_, _23235_);
  and (_23808_, _23663_, _23235_);
  nor (_23809_, _23808_, _23807_);
  and (_23810_, _23809_, _23748_);
  and (_23811_, _23810_, _23806_);
  nor (_23812_, _23811_, _23348_);
  not (_23813_, _23812_);
  and (_23814_, _23705_, _23357_);
  not (_23815_, _23814_);
  nor (_23816_, _23736_, _23356_);
  not (_23817_, _23816_);
  and (_23818_, _23691_, _23355_);
  and (_23819_, _23700_, _23348_);
  nor (_23820_, _23819_, _23818_);
  and (_23821_, _23820_, _23817_);
  and (_23822_, _23821_, _23815_);
  and (_23823_, _23822_, _23813_);
  and (_23824_, _23823_, _23805_);
  nor (_23825_, _23824_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23826_, _23339_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23827_, _23826_, _23521_);
  or (_23828_, _23827_, _23825_);
  or (_23829_, _23828_, _23787_);
  and (_23830_, _23829_, _23100_);
  and (_23831_, _23830_, _23780_);
  or (_02939_, _23831_, _23783_);
  not (_23832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  not (_23833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_23834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_23835_, _23834_, _23833_);
  nor (_23836_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_23837_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_23838_, _23837_, _23836_);
  and (_23839_, _23838_, _23835_);
  and (_23840_, _23839_, _23832_);
  not (_23841_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand (_23842_, _22739_, _23841_);
  nand (_23843_, _23842_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_23844_, _23843_, _23840_);
  and (_26925_, _23844_, _23049_);
  and (_26924_, _23049_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_23845_, rst, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_26923_, _23845_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_23846_, _23218_, _23187_);
  and (_23847_, _23846_, _23170_);
  and (_23848_, _23776_, _23229_);
  and (_23849_, _23848_, _23847_);
  and (_23850_, _23849_, _23830_);
  not (_23851_, _23849_);
  and (_23852_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_09853_, _23852_, _23850_);
  and (_23853_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _23049_);
  and (_23854_, _23853_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_23855_, _22739_, _22743_);
  not (_23856_, _23855_);
  not (_23857_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_23858_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_23859_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_23860_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_23861_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_23862_, _23861_, _23859_);
  and (_23863_, _23862_, _23860_);
  nor (_23864_, _23863_, _23859_);
  nor (_23865_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_23866_, _23865_, _23858_);
  not (_23867_, _23866_);
  nor (_23868_, _23867_, _23864_);
  nor (_23869_, _23868_, _23858_);
  not (_23870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_23871_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_23872_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_23873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_23874_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_23875_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_23876_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_23877_, _23876_, _23875_);
  and (_23878_, _23877_, _23874_);
  and (_23879_, _23878_, _23873_);
  nor (_23880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_23882_, _23880_, _23879_);
  and (_23883_, _23882_, _23872_);
  and (_23884_, _23883_, _23871_);
  and (_23885_, _23884_, _23870_);
  and (_23886_, _23885_, _23869_);
  nor (_23887_, _23886_, _23857_);
  and (_23888_, _23885_, _23857_);
  and (_23889_, _23888_, _23869_);
  nor (_23890_, _23889_, _23887_);
  not (_23891_, _23890_);
  and (_23892_, _23882_, _23869_);
  and (_23893_, _23892_, _23872_);
  nor (_23894_, _23893_, _23871_);
  and (_23895_, _23884_, _23869_);
  nor (_23896_, _23895_, _23894_);
  not (_23897_, _23896_);
  nor (_23898_, _23892_, _23872_);
  or (_23899_, _23898_, _23893_);
  not (_23900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_23901_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_23902_, _23879_, _23869_);
  and (_23903_, _23902_, _23901_);
  nor (_23904_, _23903_, _23900_);
  or (_23905_, _23904_, _23892_);
  and (_23906_, _23878_, _23869_);
  nor (_23907_, _23906_, _23873_);
  or (_23908_, _23907_, _23902_);
  and (_23909_, _23877_, _23869_);
  nor (_23910_, _23909_, _23874_);
  or (_23911_, _23910_, _23906_);
  and (_23912_, _23876_, _23869_);
  nor (_23913_, _23912_, _23875_);
  or (_23914_, _23913_, _23909_);
  not (_23915_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_23916_, _23869_, _23915_);
  nor (_23918_, _23869_, _23915_);
  nor (_23919_, _23918_, _23916_);
  not (_23920_, _23919_);
  nor (_23921_, _22804_, _22777_);
  and (_23922_, _22855_, _22830_);
  and (_23923_, _23922_, _23921_);
  not (_23925_, _22909_);
  and (_23926_, _22934_, _23925_);
  not (_23928_, _22883_);
  nor (_23929_, _22968_, _23928_);
  and (_23930_, _23929_, _23926_);
  and (_23931_, _23930_, _23923_);
  not (_23932_, _22830_);
  not (_23933_, _22804_);
  and (_23934_, _22855_, _22777_);
  and (_23935_, _23934_, _23933_);
  and (_23936_, _23935_, _23932_);
  nor (_23937_, _22968_, _22883_);
  and (_23938_, _22934_, _22909_);
  and (_23939_, _23938_, _23937_);
  and (_23940_, _23939_, _23936_);
  nor (_23941_, _22855_, _22777_);
  nor (_23942_, _23932_, _22804_);
  and (_23943_, _23942_, _23941_);
  and (_23944_, _22968_, _22883_);
  and (_23945_, _23944_, _23938_);
  not (_23946_, _22934_);
  and (_23947_, _23946_, _22909_);
  and (_23948_, _22968_, _23928_);
  nor (_23949_, _23948_, _23929_);
  and (_23950_, _23949_, _23947_);
  or (_23951_, _23950_, _23945_);
  and (_23952_, _23951_, _23943_);
  or (_23953_, _23952_, _23940_);
  or (_23954_, _23953_, _23931_);
  not (_23955_, _23936_);
  and (_23956_, _23947_, _23944_);
  and (_23957_, _23938_, _23929_);
  nor (_23958_, _23957_, _23956_);
  nor (_23959_, _23958_, _23955_);
  not (_23960_, _23943_);
  and (_23961_, _23948_, _23947_);
  nor (_23962_, _23961_, _23957_);
  nor (_23963_, _23962_, _23960_);
  or (_23964_, _23963_, _23959_);
  not (_23965_, _23923_);
  and (_23966_, _22883_, _22909_);
  and (_23967_, _23966_, _22934_);
  and (_23968_, _23947_, _23937_);
  nor (_23969_, _23968_, _23967_);
  nor (_23970_, _23969_, _23965_);
  nor (_23971_, _22934_, _22909_);
  and (_23972_, _23971_, _22883_);
  and (_23973_, _23972_, _23936_);
  or (_23974_, _23973_, _23970_);
  or (_23975_, _23974_, _23964_);
  or (_23976_, _23975_, _23954_);
  and (_23977_, _23942_, _23934_);
  and (_23978_, _23977_, _23961_);
  not (_23979_, _23978_);
  and (_23980_, _23945_, _23936_);
  and (_23982_, _23971_, _23949_);
  and (_23983_, _23982_, _23923_);
  nor (_23985_, _23983_, _23980_);
  and (_23986_, _23985_, _23979_);
  nor (_23987_, _23943_, _23935_);
  and (_23988_, _23948_, _23938_);
  and (_23989_, _23988_, _23936_);
  nor (_23990_, _23989_, _23930_);
  nor (_23991_, _23990_, _23987_);
  not (_23992_, _23991_);
  nand (_23993_, _23992_, _23986_);
  or (_23994_, _23993_, _23976_);
  and (_23995_, _23944_, _23926_);
  not (_23996_, _23995_);
  nor (_23997_, _23996_, _23987_);
  and (_23998_, _23948_, _23926_);
  or (_23999_, _23943_, _22804_);
  and (_24000_, _23999_, _23998_);
  or (_24001_, _24000_, _23997_);
  and (_24002_, _23961_, _23936_);
  not (_24003_, _22855_);
  and (_24004_, _23921_, _24003_);
  and (_24005_, _24004_, _23932_);
  and (_24006_, _24005_, _23995_);
  nor (_24007_, _24006_, _24002_);
  not (_24008_, _24007_);
  and (_24009_, _23995_, _23923_);
  and (_24010_, _23971_, _23948_);
  and (_24011_, _24010_, _23923_);
  or (_24012_, _24011_, _24009_);
  or (_24013_, _24012_, _24008_);
  or (_24014_, _24013_, _24001_);
  and (_24015_, _23947_, _23929_);
  nor (_24016_, _24015_, _23998_);
  nor (_24017_, _24016_, _23955_);
  and (_24018_, _23972_, _23943_);
  nor (_24019_, _24018_, _24017_);
  nand (_24020_, _24015_, _23999_);
  nand (_24021_, _24020_, _24019_);
  and (_24022_, _24005_, _23930_);
  and (_24023_, _23956_, _23923_);
  nor (_24024_, _24023_, _24022_);
  not (_24025_, _24024_);
  and (_24026_, _23945_, _22804_);
  and (_24027_, _23926_, _23928_);
  and (_24029_, _24027_, _23923_);
  or (_24030_, _24029_, _24026_);
  or (_24031_, _24030_, _24025_);
  or (_24032_, _24031_, _24021_);
  and (_24033_, _23961_, _23923_);
  nor (_24034_, _23941_, _23934_);
  not (_24035_, _24034_);
  nor (_24036_, _22968_, _22804_);
  and (_24037_, _24036_, _24027_);
  and (_24038_, _24037_, _24035_);
  and (_24039_, _23961_, _22804_);
  or (_24040_, _24039_, _24038_);
  or (_24041_, _24040_, _24033_);
  and (_24042_, _24015_, _23923_);
  and (_24043_, _23971_, _23928_);
  and (_24044_, _24043_, _23936_);
  or (_24046_, _24044_, _24042_);
  or (_24047_, _24046_, _24041_);
  and (_24048_, _24003_, _22777_);
  not (_24049_, _22968_);
  nor (_24050_, _24049_, _22804_);
  and (_24051_, _24050_, _24048_);
  and (_24052_, _24051_, _24027_);
  and (_24053_, _23947_, _23928_);
  and (_24054_, _24051_, _24053_);
  nor (_24055_, _24054_, _24052_);
  or (_24056_, _23998_, _23956_);
  nand (_24057_, _24056_, _23977_);
  nand (_24058_, _24057_, _24055_);
  and (_24059_, _23968_, _22804_);
  and (_24060_, _24043_, _23977_);
  or (_24061_, _24060_, _24059_);
  and (_24062_, _24048_, _24036_);
  and (_24063_, _24062_, _23947_);
  and (_24064_, _22855_, _23932_);
  and (_24065_, _24064_, _23921_);
  or (_24067_, _24065_, _24063_);
  or (_24068_, _24067_, _24061_);
  or (_24069_, _24068_, _24058_);
  or (_24070_, _24069_, _24047_);
  or (_24071_, _24070_, _24032_);
  or (_24072_, _24071_, _24014_);
  nor (_24073_, _24072_, _23994_);
  nor (_24074_, _23862_, _23860_);
  nor (_24075_, _24074_, _23863_);
  not (_24076_, _24075_);
  nor (_24077_, _24076_, _24073_);
  and (_24078_, _24024_, _24019_);
  and (_24079_, _24078_, _24007_);
  nor (_24080_, _24054_, _24039_);
  and (_24081_, _23937_, _23926_);
  and (_24083_, _24081_, _24005_);
  nor (_24084_, _24083_, _24011_);
  and (_24085_, _24084_, _24080_);
  and (_24086_, _24085_, _23986_);
  and (_24087_, _24086_, _24079_);
  not (_24088_, _24087_);
  nor (_24089_, _24088_, _24073_);
  not (_24091_, _24089_);
  nor (_24092_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_24093_, _24092_, _23860_);
  and (_24094_, _24093_, _24091_);
  and (_24095_, _24076_, _24073_);
  nor (_24096_, _24095_, _24077_);
  and (_24097_, _24096_, _24094_);
  nor (_24098_, _24097_, _24077_);
  not (_24099_, _24098_);
  and (_24100_, _23867_, _23864_);
  nor (_24101_, _24100_, _23868_);
  and (_24102_, _24101_, _24099_);
  and (_24103_, _24102_, _23920_);
  not (_24104_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_24105_, _23916_, _24104_);
  or (_24106_, _24105_, _23912_);
  and (_24107_, _24106_, _24103_);
  and (_24108_, _24107_, _23914_);
  and (_24109_, _24108_, _23911_);
  and (_24110_, _24109_, _23908_);
  nor (_24112_, _23902_, _23901_);
  or (_24113_, _24112_, _23903_);
  and (_24114_, _24113_, _24110_);
  and (_24115_, _24114_, _23905_);
  and (_24116_, _24115_, _23899_);
  and (_24117_, _24116_, _23897_);
  nor (_24118_, _23895_, _23870_);
  or (_24119_, _24118_, _23886_);
  and (_24120_, _24119_, _24117_);
  and (_24121_, _24120_, _23891_);
  not (_24122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_24123_, _23889_, _24122_);
  and (_24124_, _23889_, _24122_);
  or (_24125_, _24124_, _24123_);
  and (_24126_, _24125_, _24121_);
  and (_24127_, _24124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_24128_, _24124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_24129_, _24128_, _24127_);
  and (_24130_, _24129_, _24126_);
  nor (_24131_, _24129_, _24126_);
  or (_24132_, _24131_, _24130_);
  or (_24133_, _24132_, _23856_);
  or (_24134_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_24135_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_24136_, _24135_, _24134_);
  and (_24137_, _24136_, _24133_);
  or (_26922_[15], _24137_, _23854_);
  and (_24138_, _22992_, _22862_);
  and (_24139_, _24138_, _23040_);
  not (_24140_, _24139_);
  and (_24141_, _22975_, _22972_);
  nand (_24142_, _24141_, _22989_);
  not (_24143_, _22808_);
  nand (_24144_, _24141_, _24143_);
  and (_24145_, _24144_, _24142_);
  and (_24146_, _22991_, _22981_);
  and (_24148_, _24146_, _22862_);
  or (_24149_, _24138_, _24148_);
  and (_24150_, _22860_, _22835_);
  and (_24151_, _24150_, _23051_);
  and (_24152_, _24151_, _23018_);
  and (_24153_, _24151_, _24141_);
  and (_24154_, _23052_, _24141_);
  or (_24155_, _24154_, _24153_);
  or (_24156_, _24155_, _24152_);
  nor (_24157_, _24156_, _24149_);
  nand (_24158_, _24157_, _24145_);
  nand (_24159_, _24158_, _22944_);
  and (_24160_, _24159_, _24140_);
  not (_24161_, _22944_);
  and (_24162_, _23030_, _22862_);
  nor (_24163_, _24162_, _23056_);
  nor (_24164_, _22973_, _22808_);
  and (_24165_, _24164_, _23017_);
  nor (_24166_, _24165_, _22985_);
  and (_24167_, _24166_, _24163_);
  nor (_24168_, _24167_, _24161_);
  not (_24169_, _24168_);
  and (_24170_, _24169_, _24160_);
  and (_24171_, _23027_, _22997_);
  and (_24172_, _24171_, _23040_);
  nor (_24173_, _24172_, _23043_);
  and (_24174_, _24173_, _24159_);
  nand (_24175_, _24174_, _24140_);
  and (_24176_, _24150_, _22809_);
  nor (_24177_, _24176_, _24171_);
  nor (_24178_, _24177_, _23061_);
  and (_24179_, _22985_, _22944_);
  nor (_24180_, _24179_, _24178_);
  nor (_24182_, _24180_, _24175_);
  nor (_24183_, _24182_, _24170_);
  not (_24184_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_24185_, _22739_, _23253_);
  and (_24186_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24188_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_24189_, _22746_, _24188_);
  nor (_24191_, _22751_, _22895_);
  or (_24192_, _24191_, _24189_);
  and (_24193_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_24194_, _22767_, _22901_);
  or (_24195_, _24194_, _24193_);
  or (_24196_, _24195_, _24192_);
  and (_24198_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_24199_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_24200_, _24199_, _24198_);
  or (_24201_, _24200_, _24196_);
  and (_24202_, _24201_, _22743_);
  or (_24203_, _24202_, _24186_);
  and (_24204_, _24203_, _22739_);
  nor (_24205_, _24204_, _24185_);
  and (_24206_, _24205_, _24175_);
  and (_24207_, _24174_, _24140_);
  nor (_24208_, _22739_, _23250_);
  nor (_24209_, _22746_, _22901_);
  nor (_24210_, _22767_, _22895_);
  nor (_24211_, _24210_, _24209_);
  and (_24212_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_24213_, _22751_, _22897_);
  nor (_24214_, _24213_, _24212_);
  and (_24216_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_24217_, _22759_, _24188_);
  nor (_24218_, _24217_, _24216_);
  and (_24219_, _24218_, _24214_);
  and (_24220_, _24219_, _24211_);
  nor (_24221_, _24220_, _23856_);
  nor (_24222_, _24221_, _24208_);
  and (_24223_, _24222_, _24207_);
  nor (_24224_, _24223_, _24206_);
  and (_24225_, _24224_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_24226_, _24224_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_24227_, _24226_);
  nor (_24228_, _22739_, _23555_);
  or (_24230_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22743_);
  and (_24231_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_24232_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_24233_, _24232_, _24231_);
  nor (_24234_, _22751_, _22919_);
  not (_24235_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_24236_, _22746_, _24235_);
  nor (_24237_, _22767_, _22914_);
  or (_24238_, _24237_, _24236_);
  or (_24239_, _24238_, _24234_);
  or (_24240_, _24239_, _24233_);
  and (_24241_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_24242_, _24241_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_24243_, _24242_, _24240_);
  and (_24244_, _24243_, _22739_);
  and (_24245_, _24244_, _24230_);
  nor (_24247_, _24245_, _24228_);
  and (_24248_, _24247_, _24175_);
  nor (_24249_, _22739_, _23553_);
  nor (_24250_, _22746_, _22914_);
  nor (_24251_, _22767_, _22919_);
  nor (_24252_, _24251_, _24250_);
  and (_24253_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_24254_, _22751_, _22921_);
  nor (_24255_, _24254_, _24253_);
  and (_24256_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_24257_, _22759_, _24235_);
  nor (_24258_, _24257_, _24256_);
  and (_24259_, _24258_, _24255_);
  and (_24260_, _24259_, _24252_);
  nor (_24261_, _24260_, _23856_);
  nor (_24262_, _24261_, _24249_);
  and (_24263_, _24262_, _24207_);
  nor (_24264_, _24263_, _24248_);
  and (_24265_, _24264_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_24266_, _24265_);
  nor (_24267_, _24264_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_24268_, _24267_, _24265_);
  nor (_24269_, _22739_, _23294_);
  and (_24270_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24271_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_24272_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_24273_, _24272_, _24271_);
  and (_24274_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_24275_, _22767_, _22875_);
  or (_24276_, _24275_, _24274_);
  nor (_24277_, _22751_, _22868_);
  not (_24278_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_24279_, _22746_, _24278_);
  or (_24280_, _24279_, _24277_);
  or (_24281_, _24280_, _24276_);
  or (_24282_, _24281_, _24273_);
  and (_24283_, _24282_, _22743_);
  or (_24284_, _24283_, _24270_);
  and (_24285_, _24284_, _22739_);
  nor (_24286_, _24285_, _24269_);
  and (_24287_, _24286_, _24175_);
  nor (_24288_, _22739_, _23292_);
  nor (_24289_, _22746_, _22875_);
  nor (_24290_, _22767_, _22868_);
  nor (_24291_, _24290_, _24289_);
  and (_24292_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_24293_, _22751_, _22871_);
  nor (_24294_, _24293_, _24292_);
  and (_24295_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_24296_, _22759_, _24278_);
  nor (_24297_, _24296_, _24295_);
  and (_24298_, _24297_, _24294_);
  and (_24299_, _24298_, _24291_);
  nor (_24300_, _24299_, _23856_);
  nor (_24301_, _24300_, _24288_);
  and (_24302_, _24301_, _24207_);
  nor (_24303_, _24302_, _24287_);
  nor (_24304_, _24303_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_24305_, _24303_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_24306_, _22739_, _23331_);
  not (_24307_, _22739_);
  and (_24308_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_24310_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_24311_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_24313_, _24311_, _24310_);
  and (_24314_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_24315_, _22842_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_24316_, _24315_, _24314_);
  and (_24317_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_24318_, _22951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_24319_, _24318_, _24317_);
  and (_24320_, _24319_, _24316_);
  and (_24321_, _24320_, _24313_);
  nor (_24322_, _24321_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_24323_, _24322_, _24308_);
  nor (_24324_, _24323_, _24307_);
  nor (_24325_, _24324_, _24306_);
  and (_24326_, _24325_, _24175_);
  nor (_24327_, _22739_, _23333_);
  and (_24328_, _22951_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_24329_, _22842_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_24330_, _24329_, _24328_);
  and (_24331_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_24332_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_24333_, _24332_, _24331_);
  and (_24334_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_24335_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_24336_, _24335_, _24334_);
  and (_24337_, _24336_, _24333_);
  and (_24338_, _24337_, _24330_);
  nor (_24339_, _24338_, _23856_);
  nor (_24340_, _24339_, _24327_);
  and (_24341_, _24340_, _24207_);
  nor (_24342_, _24341_, _24326_);
  nand (_24343_, _24342_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_24344_, _22739_, _23363_);
  and (_24345_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24346_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_24347_, _22746_, _24346_);
  nor (_24348_, _22751_, _22785_);
  or (_24349_, _24348_, _24347_);
  and (_24350_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_24351_, _22767_, _22794_);
  or (_24352_, _24351_, _24350_);
  or (_24353_, _24352_, _24349_);
  and (_24354_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_24355_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_24356_, _24355_, _24354_);
  or (_24357_, _24356_, _24353_);
  and (_24358_, _24357_, _22743_);
  or (_24359_, _24358_, _24345_);
  and (_24360_, _24359_, _22739_);
  nor (_24361_, _24360_, _24344_);
  and (_24362_, _24361_, _24175_);
  nor (_24363_, _22739_, _23361_);
  nor (_24364_, _22746_, _22794_);
  nor (_24365_, _22767_, _22785_);
  nor (_24366_, _24365_, _24364_);
  and (_24367_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_24369_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_24370_, _24369_, _24367_);
  nor (_24372_, _22759_, _24346_);
  nor (_24373_, _22751_, _22788_);
  nor (_24374_, _24373_, _24372_);
  and (_24375_, _24374_, _24370_);
  and (_24376_, _24375_, _24366_);
  nor (_24377_, _24376_, _23856_);
  nor (_24378_, _24377_, _24363_);
  and (_24379_, _24378_, _24207_);
  nor (_24380_, _24379_, _24362_);
  and (_24381_, _24380_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_24382_, _24380_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_24383_, _24382_, _24381_);
  nor (_24384_, _22739_, _23407_);
  or (_24385_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _22743_);
  and (_24386_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_24387_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_24388_, _24387_, _24386_);
  nor (_24389_, _22751_, _22744_);
  not (_24390_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_24391_, _22746_, _24390_);
  nor (_24392_, _22767_, _22758_);
  or (_24393_, _24392_, _24391_);
  or (_24394_, _24393_, _24389_);
  or (_24395_, _24394_, _24388_);
  and (_24396_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_24397_, _24396_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_24398_, _24397_, _24395_);
  and (_24399_, _24398_, _22739_);
  and (_24400_, _24399_, _24385_);
  nor (_24401_, _24400_, _24384_);
  not (_24402_, _24401_);
  or (_24403_, _24402_, _24207_);
  nor (_24404_, _22739_, _23405_);
  nor (_24405_, _22746_, _22758_);
  nor (_24406_, _22767_, _22744_);
  nor (_24407_, _24406_, _24405_);
  and (_24408_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_24409_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_24410_, _24409_, _24408_);
  nor (_24411_, _22759_, _24390_);
  nor (_24412_, _22751_, _22765_);
  nor (_24413_, _24412_, _24411_);
  and (_24414_, _24413_, _24410_);
  and (_24415_, _24414_, _24407_);
  nor (_24416_, _24415_, _23856_);
  nor (_24417_, _24416_, _24404_);
  not (_24418_, _24417_);
  or (_24419_, _24418_, _24175_);
  nand (_24420_, _24419_, _24403_);
  or (_24421_, _24420_, _23391_);
  not (_24422_, _24421_);
  nor (_24423_, _22739_, _23428_);
  and (_24424_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24425_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_24426_, _22746_, _24425_);
  nor (_24427_, _22751_, _22839_);
  or (_24428_, _24427_, _24426_);
  and (_24429_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_24430_, _22767_, _22837_);
  or (_24431_, _24430_, _24429_);
  or (_24432_, _24431_, _24428_);
  and (_24433_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_24434_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_24435_, _24434_, _24433_);
  or (_24436_, _24435_, _24432_);
  and (_24437_, _24436_, _22743_);
  or (_24438_, _24437_, _24424_);
  and (_24439_, _24438_, _22739_);
  nor (_24440_, _24439_, _24423_);
  not (_24441_, _24440_);
  or (_24442_, _24441_, _24207_);
  nor (_24443_, _22739_, _23430_);
  nor (_24444_, _22746_, _22837_);
  nor (_24445_, _22767_, _22839_);
  nor (_24446_, _24445_, _24444_);
  and (_24447_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_24448_, _22752_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_24449_, _24448_, _24447_);
  and (_24450_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_24451_, _22759_, _24425_);
  nor (_24452_, _24451_, _24450_);
  and (_24453_, _24452_, _24449_);
  and (_24454_, _24453_, _24446_);
  nor (_24455_, _24454_, _23856_);
  nor (_24456_, _24455_, _24443_);
  not (_24457_, _24456_);
  or (_24458_, _24457_, _24175_);
  and (_24460_, _24458_, _24442_);
  nand (_24461_, _24460_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_24462_, _22739_, _23459_);
  and (_24464_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24465_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_24466_, _22746_, _24465_);
  nor (_24467_, _22751_, _22819_);
  or (_24468_, _24467_, _24466_);
  and (_24469_, _22960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_24470_, _22767_, _22815_);
  or (_24471_, _24470_, _24469_);
  or (_24473_, _24471_, _24468_);
  and (_24474_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_24475_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_24476_, _24475_, _24474_);
  or (_24477_, _24476_, _24473_);
  and (_24478_, _24477_, _22743_);
  or (_24479_, _24478_, _24464_);
  and (_24480_, _24479_, _22739_);
  nor (_24481_, _24480_, _24462_);
  not (_24482_, _24481_);
  or (_24483_, _24482_, _24207_);
  nor (_24484_, _22739_, _23461_);
  nor (_24485_, _22746_, _22815_);
  nor (_24486_, _22767_, _22819_);
  nor (_24487_, _24486_, _24485_);
  and (_24489_, _22756_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_24490_, _22763_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_24491_, _24490_, _24489_);
  nor (_24492_, _22759_, _24465_);
  nor (_24493_, _22751_, _22811_);
  nor (_24494_, _24493_, _24492_);
  and (_24495_, _24494_, _24491_);
  and (_24496_, _24495_, _24487_);
  nor (_24497_, _24496_, _23856_);
  nor (_24498_, _24497_, _24484_);
  not (_24499_, _24498_);
  or (_24500_, _24499_, _24175_);
  and (_24502_, _24500_, _24483_);
  and (_24503_, _24502_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_24504_, _24460_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_24505_, _24504_, _24461_);
  and (_24506_, _24505_, _24503_);
  not (_24507_, _24506_);
  nand (_24508_, _24507_, _24461_);
  nand (_24509_, _24420_, _23391_);
  and (_24510_, _24509_, _24421_);
  and (_24512_, _24510_, _24508_);
  or (_24513_, _24512_, _24422_);
  and (_24514_, _24513_, _24383_);
  or (_24515_, _24514_, _24381_);
  or (_24516_, _24342_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_24517_, _24516_, _24343_);
  nand (_24518_, _24517_, _24515_);
  nand (_24519_, _24518_, _24343_);
  nor (_24520_, _24519_, _24305_);
  nor (_24521_, _24520_, _24304_);
  nand (_24522_, _24521_, _24268_);
  nand (_24523_, _24522_, _24266_);
  and (_24524_, _24523_, _24227_);
  or (_24525_, _24524_, _24225_);
  or (_24526_, _24525_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_24527_, _24526_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_24528_, _24527_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_24529_, _24528_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_24530_, _24529_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_24531_, _24530_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_24532_, _24531_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_24533_, _24532_, _24224_);
  not (_24534_, _24224_);
  not (_24535_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_24536_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_24537_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_24538_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_24539_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_24540_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_24541_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_24542_, _24524_, _24225_);
  or (_24543_, _24542_, _24541_);
  or (_24544_, _24543_, _24540_);
  or (_24545_, _24544_, _24539_);
  or (_24546_, _24545_, _24538_);
  or (_24547_, _24546_, _24537_);
  or (_24548_, _24547_, _24536_);
  or (_24549_, _24548_, _24535_);
  and (_24550_, _24549_, _24534_);
  or (_24551_, _24550_, _24533_);
  nand (_24552_, _24551_, _24184_);
  or (_24553_, _24551_, _24184_);
  and (_24554_, _24553_, _24552_);
  and (_24555_, _24554_, _24183_);
  nor (_24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24557_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_24558_, _24557_);
  nand (_24559_, _24556_, _23279_);
  and (_24560_, _24559_, _24558_);
  not (_24561_, _24560_);
  or (_24562_, _23483_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_24564_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24565_, _23419_, _24564_);
  and (_24566_, _24565_, _24562_);
  or (_24567_, _24566_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24568_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24569_, _23609_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24570_, _23576_, _24564_);
  and (_24571_, _24570_, _24569_);
  or (_24572_, _24571_, _24568_);
  and (_24573_, _24572_, _24567_);
  or (_24574_, _24573_, _24561_);
  nand (_24575_, _24556_, _23570_);
  nor (_24576_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_24577_, _24576_);
  and (_24578_, _24577_, _24575_);
  not (_24579_, _24578_);
  and (_24580_, _23454_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24581_, _24580_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24582_, _23647_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24583_, _23322_, _24564_);
  and (_24584_, _24583_, _24582_);
  or (_24585_, _24584_, _24568_);
  and (_24586_, _24585_, _24581_);
  or (_24587_, _24586_, _24579_);
  nand (_24588_, _24572_, _24567_);
  or (_24589_, _24588_, _24560_);
  and (_24590_, _24589_, _24574_);
  not (_24591_, _24590_);
  or (_24592_, _24591_, _24587_);
  and (_24593_, _24592_, _24574_);
  nand (_24594_, _24585_, _24581_);
  or (_24595_, _24594_, _24578_);
  and (_24596_, _24595_, _24587_);
  and (_24597_, _24596_, _24590_);
  not (_24598_, _24556_);
  or (_24599_, _24598_, _23316_);
  nor (_24600_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_24601_, _24600_);
  nand (_24603_, _24601_, _24599_);
  and (_24604_, _23483_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24605_, _24604_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24606_, _23419_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24607_, _23609_, _24564_);
  and (_24608_, _24607_, _24606_);
  or (_24609_, _24608_, _24568_);
  and (_24610_, _24609_, _24605_);
  or (_24611_, _24610_, _24603_);
  or (_24612_, _23454_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_24613_, _23647_, _24564_);
  and (_24614_, _24613_, _24612_);
  and (_24615_, _24614_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24616_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_24617_, _24616_);
  nand (_24618_, _24556_, _23348_);
  and (_24619_, _24618_, _24617_);
  not (_24620_, _24619_);
  or (_24621_, _24620_, _24615_);
  and (_24622_, _24601_, _24599_);
  nand (_24623_, _24609_, _24605_);
  or (_24624_, _24623_, _24622_);
  nand (_24625_, _24624_, _24611_);
  or (_24626_, _24625_, _24621_);
  nand (_24627_, _24626_, _24611_);
  nand (_24628_, _24627_, _24597_);
  and (_24629_, _24628_, _24593_);
  and (_24630_, _24566_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_24631_, _24630_);
  nand (_24632_, _24556_, _23378_);
  nor (_24633_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_24634_, _24633_);
  and (_24635_, _24634_, _24632_);
  nand (_24636_, _24635_, _24631_);
  or (_24637_, _24635_, _24631_);
  nand (_24638_, _24637_, _24636_);
  nand (_24639_, _24580_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24640_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_24641_, _24640_);
  or (_24642_, _24598_, _23412_);
  and (_24643_, _24642_, _24641_);
  nand (_24644_, _24643_, _24639_);
  and (_24645_, _24604_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_24646_, _24598_, _23448_);
  nor (_24647_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_24649_, _24647_);
  nand (_24650_, _24649_, _24646_);
  and (_24651_, _24650_, _24645_);
  or (_24652_, _24643_, _24639_);
  nand (_24653_, _24652_, _24644_);
  or (_24654_, _24653_, _24651_);
  and (_24655_, _24654_, _24644_);
  or (_24656_, _24655_, _24638_);
  nand (_24657_, _24656_, _24636_);
  not (_24658_, _24615_);
  or (_24659_, _24619_, _24658_);
  and (_24660_, _24659_, _24621_);
  and (_24661_, _24624_, _24611_);
  and (_24662_, _24661_, _24660_);
  and (_24663_, _24662_, _24597_);
  nand (_24664_, _24663_, _24657_);
  nand (_24665_, _24664_, _24629_);
  and (_24666_, _23577_, _23289_);
  nor (_24667_, _24666_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_24668_, _24584_, _24571_);
  or (_24669_, _23322_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_24670_, _23289_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_24671_, _24670_, _24669_);
  nor (_24672_, _24671_, _24608_);
  nand (_24673_, _24672_, _24668_);
  and (_24674_, _24673_, _24568_);
  nor (_24675_, _24674_, _24667_);
  nor (_24676_, _24614_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_24677_, _24671_, _24568_);
  nor (_24678_, _24677_, _24676_);
  not (_24679_, _24678_);
  and (_24681_, _24679_, _24675_);
  nand (_24682_, _24681_, _24665_);
  and (_24683_, _24682_, _24560_);
  not (_24684_, _24683_);
  and (_24685_, _24681_, _24665_);
  and (_24686_, _24610_, _24603_);
  not (_24687_, _24621_);
  and (_24688_, _24660_, _24657_);
  nor (_24689_, _24688_, _24687_);
  or (_24690_, _24689_, _24686_);
  and (_24691_, _24690_, _24611_);
  not (_24692_, _24691_);
  nand (_24693_, _24692_, _24596_);
  and (_24694_, _24693_, _24587_);
  nand (_24695_, _24694_, _24590_);
  or (_24696_, _24694_, _24590_);
  nand (_24697_, _24696_, _24695_);
  nand (_24698_, _24697_, _24685_);
  and (_24700_, _24698_, _24684_);
  nand (_24701_, _24698_, _24684_);
  or (_24703_, _24701_, _24679_);
  or (_24704_, _24700_, _24678_);
  or (_24705_, _24692_, _24596_);
  nand (_24706_, _24705_, _24693_);
  nand (_24707_, _24706_, _24685_);
  and (_24708_, _24682_, _24579_);
  not (_24709_, _24708_);
  and (_24710_, _24709_, _24707_);
  and (_24711_, _24710_, _24588_);
  not (_24712_, _24711_);
  nand (_24713_, _24712_, _24704_);
  nand (_24714_, _24713_, _24703_);
  and (_24715_, _24704_, _24703_);
  or (_24716_, _24710_, _24588_);
  and (_24717_, _24716_, _24712_);
  and (_24718_, _24717_, _24715_);
  nand (_24719_, _24625_, _24689_);
  or (_24720_, _24625_, _24689_);
  nand (_24721_, _24720_, _24719_);
  nand (_24722_, _24721_, _24685_);
  and (_24723_, _24682_, _24603_);
  not (_24724_, _24723_);
  and (_24725_, _24724_, _24722_);
  and (_24726_, _24725_, _24594_);
  nor (_24727_, _24660_, _24657_);
  or (_24728_, _24727_, _24688_);
  and (_24729_, _24728_, _24685_);
  and (_24730_, _24682_, _24620_);
  nor (_24731_, _24730_, _24729_);
  and (_24732_, _24731_, _24623_);
  nor (_24733_, _24725_, _24594_);
  or (_24734_, _24733_, _24726_);
  not (_24735_, _24734_);
  and (_24736_, _24735_, _24732_);
  nor (_24737_, _24736_, _24726_);
  and (_24738_, _24655_, _24638_);
  not (_24739_, _24738_);
  and (_24740_, _24739_, _24656_);
  or (_24741_, _24740_, _24682_);
  or (_24742_, _24685_, _24635_);
  and (_24743_, _24742_, _24741_);
  nor (_24744_, _24743_, _24658_);
  not (_24745_, _24744_);
  not (_24746_, _24645_);
  or (_24747_, _24682_, _24746_);
  nand (_24748_, _24747_, _24650_);
  or (_24749_, _24747_, _24650_);
  and (_24750_, _24749_, _24748_);
  nand (_24751_, _24750_, _24639_);
  or (_24752_, _24750_, _24639_);
  and (_24753_, _24752_, _24751_);
  and (_24754_, _24556_, _23476_);
  nor (_24755_, _24556_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_24756_, _24755_, _24754_);
  nor (_24757_, _24756_, _24746_);
  not (_24758_, _24757_);
  nand (_24759_, _24758_, _24753_);
  and (_24760_, _24759_, _24751_);
  and (_24761_, _24653_, _24651_);
  not (_24762_, _24761_);
  and (_24763_, _24762_, _24654_);
  or (_24764_, _24763_, _24682_);
  or (_24765_, _24685_, _24643_);
  and (_24766_, _24765_, _24764_);
  nand (_24767_, _24766_, _24631_);
  or (_24768_, _24766_, _24631_);
  and (_24769_, _24768_, _24767_);
  not (_24770_, _24769_);
  or (_24771_, _24770_, _24760_);
  and (_24772_, _24743_, _24658_);
  not (_24773_, _24772_);
  and (_24774_, _24773_, _24767_);
  nand (_24775_, _24774_, _24771_);
  and (_24776_, _24775_, _24745_);
  nor (_24777_, _24731_, _24623_);
  nor (_24778_, _24777_, _24732_);
  and (_24779_, _24735_, _24778_);
  nand (_24780_, _24779_, _24776_);
  nand (_24781_, _24780_, _24737_);
  nand (_24782_, _24781_, _24718_);
  nand (_24783_, _24782_, _24714_);
  and (_24784_, _24783_, _24675_);
  or (_24785_, _24784_, _24700_);
  nand (_24786_, _24781_, _24717_);
  and (_24787_, _24786_, _24712_);
  nand (_24788_, _24787_, _24715_);
  or (_24789_, _24787_, _24715_);
  nand (_24790_, _24789_, _24788_);
  nand (_24791_, _24790_, _24784_);
  nand (_24792_, _24791_, _24785_);
  nand (_24793_, _24792_, _23752_);
  and (_24794_, _23690_, _23234_);
  nor (_24795_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_24796_, _24795_);
  and (_24797_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_24798_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  or (_24799_, _24796_, _23576_);
  not (_24800_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_24801_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _24800_);
  not (_24802_, _24801_);
  or (_24803_, _24802_, _23354_);
  not (_24804_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_24805_, _24804_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_24806_, _24805_);
  or (_24807_, _24806_, _23628_);
  and (_24808_, _24807_, _24803_);
  nor (_24809_, _24805_, _24801_);
  or (_24810_, _23483_, _24800_);
  nand (_24811_, _24810_, _24809_);
  nand (_24812_, _24811_, _24808_);
  nand (_24813_, _24812_, _24799_);
  or (_24814_, _24813_, _23378_);
  nand (_24815_, _24795_, _23289_);
  or (_24816_, _24802_, _23607_);
  or (_24817_, _24806_, _23384_);
  and (_24818_, _24817_, _24816_);
  or (_24819_, _23454_, _24800_);
  nand (_24820_, _24819_, _24809_);
  nand (_24821_, _24820_, _24818_);
  nand (_24822_, _24821_, _24815_);
  or (_24823_, _24822_, _23348_);
  or (_24824_, _24823_, _24814_);
  not (_24825_, _24824_);
  or (_24826_, _24813_, _23669_);
  or (_24827_, _24826_, _24823_);
  nand (_24828_, _24826_, _24823_);
  and (_24829_, _24828_, _24827_);
  nand (_24830_, _24829_, _24825_);
  not (_24831_, _24830_);
  or (_24832_, _24827_, _23570_);
  and (_24833_, _24821_, _24815_);
  and (_24834_, _24833_, _23316_);
  not (_24835_, _23570_);
  and (_24836_, _24812_, _24799_);
  and (_24837_, _24836_, _24835_);
  not (_24838_, _24837_);
  nand (_24839_, _24838_, _24827_);
  and (_24840_, _24839_, _24834_);
  nand (_24841_, _24840_, _24832_);
  or (_24842_, _24837_, _24834_);
  and (_24843_, _24842_, _24841_);
  and (_24844_, _24843_, _24831_);
  not (_24845_, _24840_);
  or (_24846_, _24813_, _23279_);
  or (_24847_, _24822_, _23570_);
  or (_24848_, _24847_, _24846_);
  nand (_24849_, _24847_, _24846_);
  and (_24850_, _24849_, _24848_);
  nand (_24851_, _24850_, _24845_);
  or (_24852_, _24850_, _24845_);
  nand (_24853_, _24852_, _24851_);
  nand (_24854_, _24853_, _24844_);
  and (_24855_, _24833_, _23448_);
  and (_24856_, _24836_, _23412_);
  nand (_24857_, _24856_, _24855_);
  and (_24858_, _24836_, _23795_);
  not (_24859_, _23448_);
  or (_24860_, _24813_, _24859_);
  and (_24861_, _24833_, _23412_);
  and (_24862_, _24861_, _24860_);
  nand (_24863_, _24862_, _24858_);
  nand (_24864_, _24863_, _24857_);
  or (_24865_, _24813_, _23348_);
  or (_24866_, _24822_, _23378_);
  nand (_24867_, _24866_, _24865_);
  and (_24868_, _24867_, _24824_);
  and (_24869_, _24868_, _24864_);
  or (_24870_, _24829_, _24825_);
  and (_24871_, _24870_, _24830_);
  nand (_24872_, _24871_, _24869_);
  not (_24873_, _24872_);
  nand (_24874_, _24843_, _24831_);
  or (_24875_, _24843_, _24831_);
  and (_24876_, _24875_, _24874_);
  nand (_24877_, _24876_, _24873_);
  not (_24878_, _24877_);
  or (_24879_, _24853_, _24844_);
  and (_24880_, _24879_, _24854_);
  nand (_24881_, _24880_, _24878_);
  and (_24882_, _24881_, _24854_);
  and (_24883_, _24836_, _23448_);
  and (_24884_, _24833_, _23717_);
  and (_24885_, _24884_, _24883_);
  or (_24886_, _24856_, _24855_);
  and (_24887_, _24886_, _24857_);
  and (_24888_, _24887_, _24885_);
  or (_24889_, _24862_, _24858_);
  and (_24890_, _24889_, _24863_);
  and (_24891_, _24890_, _24888_);
  nand (_24892_, _24868_, _24864_);
  or (_24893_, _24868_, _24864_);
  and (_24894_, _24893_, _24892_);
  and (_24895_, _24894_, _24891_);
  or (_24896_, _24871_, _24869_);
  and (_24897_, _24896_, _24872_);
  nand (_24898_, _24897_, _24895_);
  not (_24899_, _24898_);
  or (_24900_, _24876_, _24873_);
  and (_24901_, _24900_, _24877_);
  and (_24902_, _24880_, _24901_);
  nand (_24903_, _24902_, _24899_);
  nand (_24904_, _24903_, _24882_);
  and (_24905_, _24833_, _23714_);
  and (_24906_, _24905_, _24838_);
  and (_24907_, _24850_, _24840_);
  and (_24908_, _24907_, _24906_);
  nor (_24909_, _24907_, _24906_);
  nor (_24910_, _24909_, _24908_);
  nand (_24911_, _24910_, _24904_);
  not (_24912_, _24908_);
  and (_24913_, _24912_, _24848_);
  nand (_24914_, _24913_, _24911_);
  nand (_24915_, _24914_, _24798_);
  or (_24916_, _24914_, _24798_);
  nand (_24917_, _24916_, _24915_);
  and (_24918_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_24919_, _24910_, _24904_);
  and (_24920_, _24919_, _24911_);
  nand (_24921_, _24920_, _24918_);
  or (_24922_, _24921_, _24917_);
  nand (_24923_, _24922_, _24915_);
  and (_24924_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_24925_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_24926_, _24925_, _24924_);
  and (_24927_, _24926_, _24923_);
  and (_24928_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_24929_, _24901_, _24899_);
  nand (_24930_, _24929_, _24877_);
  nand (_24931_, _24880_, _24930_);
  or (_24932_, _24880_, _24930_);
  and (_24933_, _24932_, _24931_);
  nand (_24934_, _24933_, _24928_);
  or (_24935_, _24933_, _24928_);
  and (_24936_, _24935_, _24934_);
  and (_24937_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_24938_, _24901_, _24899_);
  and (_24939_, _24938_, _24929_);
  nand (_24940_, _24939_, _24937_);
  or (_24941_, _24939_, _24937_);
  and (_24942_, _24941_, _24940_);
  and (_24943_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_24944_, _24897_, _24895_);
  and (_24945_, _24944_, _24898_);
  nand (_24946_, _24945_, _24943_);
  or (_24947_, _24945_, _24943_);
  and (_24948_, _24947_, _24946_);
  and (_24949_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nand (_24950_, _24894_, _24891_);
  or (_24951_, _24894_, _24891_);
  and (_24952_, _24951_, _24950_);
  nand (_24953_, _24952_, _24949_);
  and (_24954_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand (_24955_, _24890_, _24888_);
  or (_24956_, _24890_, _24888_);
  and (_24957_, _24956_, _24955_);
  nand (_24958_, _24957_, _24954_);
  and (_24959_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_24960_, _24887_, _24885_);
  nor (_24961_, _24960_, _24888_);
  and (_24962_, _24961_, _24959_);
  or (_24963_, _24957_, _24954_);
  and (_24964_, _24963_, _24958_);
  nand (_24965_, _24964_, _24962_);
  nand (_24966_, _24965_, _24958_);
  or (_24967_, _24952_, _24949_);
  and (_24968_, _24967_, _24953_);
  nand (_24969_, _24968_, _24966_);
  nand (_24970_, _24969_, _24953_);
  nand (_24971_, _24970_, _24948_);
  nand (_24972_, _24971_, _24946_);
  nand (_24973_, _24972_, _24942_);
  nand (_24974_, _24973_, _24940_);
  nand (_24975_, _24974_, _24936_);
  nand (_24976_, _24975_, _24934_);
  and (_24977_, _24916_, _24915_);
  or (_24978_, _24920_, _24918_);
  and (_24979_, _24978_, _24921_);
  and (_24980_, _24979_, _24977_);
  and (_24981_, _24926_, _24980_);
  and (_24982_, _24981_, _24976_);
  or (_24983_, _24982_, _24927_);
  and (_24984_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_24985_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_24986_, _24985_, _24984_);
  and (_24987_, _24986_, _24983_);
  nand (_24988_, _24987_, _24797_);
  and (_24989_, _24796_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_24990_, _24989_, _24988_);
  or (_24991_, _24988_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_24992_, _24991_, _24990_);
  nand (_24993_, _24992_, _24794_);
  not (_24994_, _23605_);
  and (_24995_, _23656_, _24994_);
  nor (_24996_, _23656_, _24994_);
  nor (_24997_, _24996_, _24995_);
  and (_24998_, _24997_, _23601_);
  not (_24999_, _24998_);
  nor (_25000_, _23605_, _23590_);
  and (_25001_, _23605_, _23590_);
  or (_25002_, _25001_, _25000_);
  and (_25003_, _25002_, _23238_);
  nor (_25004_, _23736_, _23591_);
  and (_25005_, _23705_, _23605_);
  nor (_25006_, _25005_, _25004_);
  and (_25007_, _23697_, _23717_);
  nor (_25008_, _23748_, _23570_);
  nor (_25009_, _25008_, _25007_);
  and (_25010_, _23718_, _23710_);
  and (_25011_, _23691_, _23290_);
  and (_25012_, _23700_, _23279_);
  nor (_25013_, _25012_, _25011_);
  and (_25014_, _23711_, _23714_);
  not (_25015_, _25014_);
  nand (_25017_, _25015_, _25013_);
  nor (_25018_, _25017_, _25010_);
  and (_25019_, _25018_, _25009_);
  not (_25020_, _23742_);
  nor (_25021_, _23536_, _23603_);
  or (_25022_, _25021_, _25020_);
  nor (_25023_, _25022_, _23680_);
  and (_25024_, _23798_, _23661_);
  and (_25025_, _25024_, _23316_);
  nor (_25026_, _25025_, _23710_);
  and (_25027_, _23793_, _23348_);
  and (_25028_, _25027_, _23670_);
  nor (_25029_, _25028_, _23536_);
  or (_25030_, _25029_, _23677_);
  nor (_25031_, _25030_, _25026_);
  nor (_25032_, _25031_, _23714_);
  and (_25033_, _25031_, _23714_);
  nor (_25034_, _25033_, _25032_);
  and (_25035_, _25034_, _23744_);
  nor (_25036_, _25035_, _25023_);
  nor (_25037_, _23670_, _23279_);
  nor (_25038_, _25037_, _23667_);
  and (_25039_, _25038_, _23536_);
  nor (_25040_, _25039_, _23672_);
  and (_25041_, _25040_, _23279_);
  nor (_25042_, _25040_, _23279_);
  nor (_25043_, _25042_, _25041_);
  nor (_25044_, _25043_, _23679_);
  not (_25045_, _25044_);
  and (_25046_, _25045_, _25036_);
  and (_25047_, _25046_, _25019_);
  and (_25048_, _25047_, _25006_);
  not (_25049_, _25048_);
  nor (_25050_, _25049_, _25003_);
  and (_25051_, _25050_, _24999_);
  and (_25052_, _25051_, _24993_);
  nand (_25053_, _25052_, _24793_);
  and (_25055_, _25053_, _23043_);
  not (_25056_, _23041_);
  and (_25057_, _24149_, _25056_);
  not (_25058_, _23048_);
  nand (_25059_, _23010_, _22948_);
  not (_25060_, _25059_);
  and (_25061_, _24151_, _23010_);
  nor (_25062_, _25061_, _25060_);
  and (_25063_, _22976_, _22862_);
  and (_25064_, _23027_, _22984_);
  nor (_25065_, _25064_, _25063_);
  and (_25066_, _25065_, _25062_);
  and (_25068_, _24141_, _22862_);
  not (_25069_, _25068_);
  and (_25070_, _23027_, _24141_);
  and (_25071_, _23017_, _22973_);
  and (_25072_, _23027_, _25071_);
  nor (_25073_, _25072_, _25070_);
  and (_25074_, _24146_, _24151_);
  nor (_25075_, _25074_, _24152_);
  and (_25076_, _25075_, _25073_);
  and (_25077_, _25076_, _25069_);
  and (_25078_, _25077_, _25066_);
  and (_25079_, _23030_, _23027_);
  and (_25080_, _22994_, _22948_);
  nor (_25081_, _25080_, _25079_);
  and (_25082_, _24151_, _23009_);
  and (_25083_, _22976_, _24143_);
  or (_25084_, _25083_, _25082_);
  nor (_25085_, _25084_, _24153_);
  and (_25086_, _25085_, _25081_);
  and (_25087_, _23027_, _23018_);
  and (_25088_, _23027_, _22976_);
  nor (_25089_, _25088_, _25087_);
  and (_25090_, _23027_, _22982_);
  and (_25091_, _24151_, _23030_);
  nor (_25092_, _25091_, _25090_);
  and (_25093_, _25092_, _25089_);
  and (_25094_, _25093_, _25086_);
  nand (_25095_, _23032_, _22948_);
  and (_25096_, _23017_, _22862_);
  not (_25097_, _25096_);
  and (_25098_, _25097_, _25095_);
  and (_25099_, _24151_, _23032_);
  and (_25100_, _24151_, _25071_);
  or (_25101_, _25100_, _25099_);
  and (_25102_, _24151_, _22995_);
  nor (_25103_, _25102_, _25101_);
  and (_25104_, _25103_, _25098_);
  and (_25105_, _24151_, _22982_);
  and (_25106_, _22997_, _22973_);
  and (_25107_, _25106_, _24151_);
  or (_25108_, _25107_, _25105_);
  nor (_25109_, _25108_, _23028_);
  and (_25110_, _22989_, _22973_);
  and (_25111_, _25110_, _22975_);
  nor (_25112_, _24149_, _25111_);
  and (_25113_, _25112_, _25109_);
  and (_25114_, _25113_, _25104_);
  and (_25115_, _25114_, _25094_);
  nand (_25116_, _25115_, _25078_);
  nand (_25117_, _25116_, _23040_);
  nor (_25118_, _23057_, _23043_);
  nand (_25119_, _25118_, _25117_);
  nand (_25120_, _25119_, _22734_);
  and (_25121_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_25122_, _25121_);
  and (_25123_, _25122_, _25120_);
  and (_25124_, _25123_, _25058_);
  and (_25125_, _25124_, _23065_);
  nor (_25126_, _23183_, _23098_);
  nor (_25127_, _23071_, _23068_);
  and (_25128_, _25127_, _23763_);
  and (_25129_, _25128_, _23153_);
  and (_25130_, _23167_, _23137_);
  and (_25131_, _25130_, _23215_);
  and (_25132_, _25131_, _25129_);
  and (_25133_, _25132_, _25126_);
  nor (_25134_, _23202_, _23122_);
  and (_25135_, _25134_, _25133_);
  not (_25136_, _25135_);
  and (_25137_, _25136_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_25138_, _25136_, _23824_);
  nor (_25139_, _25138_, _25137_);
  not (_25140_, _25139_);
  and (_25141_, _25136_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_25142_, _23811_, _23378_);
  nor (_25143_, _23797_, _23795_);
  nor (_25144_, _25143_, _23799_);
  nor (_25145_, _23792_, _23378_);
  nor (_25146_, _25145_, _23793_);
  nor (_25147_, _25146_, _23536_);
  or (_25148_, _25147_, _25144_);
  and (_25149_, _25148_, _23744_);
  and (_25150_, _23705_, _23387_);
  nor (_25151_, _23736_, _23386_);
  and (_25152_, _23691_, _23385_);
  and (_25153_, _23742_, _23647_);
  and (_25154_, _23700_, _23378_);
  or (_25155_, _25154_, _25153_);
  or (_25156_, _25155_, _25152_);
  or (_25157_, _25156_, _25151_);
  or (_25158_, _25157_, _25150_);
  or (_25159_, _25158_, _25149_);
  nor (_25160_, _25159_, _25142_);
  nor (_25161_, _25136_, _25160_);
  nor (_25162_, _25161_, _25141_);
  and (_25163_, _25162_, _22835_);
  and (_25164_, _25163_, _25140_);
  and (_25165_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_25166_, _25162_, _22835_);
  and (_25167_, _25166_, _25139_);
  and (_25168_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_25169_, _25168_, _25165_);
  nor (_25170_, _25162_, _22836_);
  and (_25171_, _25170_, _25139_);
  and (_25172_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_25173_, _25162_, _22836_);
  and (_25174_, _25173_, _25139_);
  and (_25175_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_25176_, _25175_, _25172_);
  and (_25177_, _25176_, _25169_);
  and (_25178_, _23122_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_25179_, _25139_, _23123_);
  nor (_25180_, _25179_, _25178_);
  not (_25181_, _23167_);
  and (_25182_, _25181_, _23137_);
  nor (_25183_, _25182_, _22836_);
  nor (_25184_, _25130_, _22835_);
  nor (_25185_, _25184_, _25183_);
  and (_25186_, _23183_, _23098_);
  and (_25187_, _23067_, _23763_);
  and (_25188_, _25187_, _23215_);
  and (_25189_, _25188_, _23201_);
  and (_25190_, _25189_, _25186_);
  and (_25191_, _25190_, _25185_);
  and (_25192_, _25162_, _23154_);
  nor (_25193_, _25162_, _23154_);
  nor (_25194_, _25193_, _25192_);
  and (_25195_, _25194_, _25191_);
  and (_25196_, _25195_, _25180_);
  not (_25197_, _25196_);
  and (_25198_, _25170_, _25140_);
  and (_25199_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_25200_, _25173_, _25140_);
  and (_25201_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_25202_, _25201_, _25199_);
  and (_25203_, _25166_, _25140_);
  and (_25204_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_25205_, _25163_, _25139_);
  and (_25206_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_25207_, _25206_, _25204_);
  and (_25208_, _25207_, _25202_);
  and (_25209_, _25208_, _25197_);
  and (_25210_, _25209_, _25177_);
  and (_25211_, _25196_, _25160_);
  nor (_25212_, _25211_, _25210_);
  and (_25213_, _25212_, _25125_);
  not (_25214_, _24378_);
  not (_25215_, _25123_);
  and (_25216_, _23065_, _23048_);
  and (_25217_, _25216_, _25215_);
  and (_25218_, _25217_, _25214_);
  nor (_25219_, _25218_, _25213_);
  nor (_25220_, _25123_, _23048_);
  and (_25221_, _25220_, _23065_);
  not (_25222_, _25221_);
  and (_25223_, _23215_, _23137_);
  and (_25224_, _25223_, _25181_);
  and (_25225_, _23201_, _23122_);
  and (_25226_, _25225_, _23777_);
  and (_25227_, _25226_, _25129_);
  and (_25228_, _25227_, _25224_);
  not (_25230_, _25228_);
  nor (_25231_, _25160_, _25230_);
  and (_25232_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_25233_, _25231_, _25232_);
  and (_25234_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_25235_, _23742_, _23419_);
  and (_25236_, _23476_, _24859_);
  or (_25237_, _25236_, _23536_);
  or (_25238_, _23796_, _23710_);
  and (_25239_, _25238_, _25237_);
  nand (_25240_, _25239_, _23412_);
  or (_25241_, _25239_, _23412_);
  and (_25242_, _25241_, _25240_);
  and (_25243_, _25242_, _23744_);
  nor (_25244_, _25243_, _25235_);
  not (_25245_, _23811_);
  and (_25246_, _25245_, _23412_);
  not (_25247_, _25246_);
  and (_25248_, _23705_, _23422_);
  nor (_25249_, _23736_, _23421_);
  not (_25250_, _25249_);
  and (_25251_, _23691_, _23420_);
  not (_25252_, _23412_);
  and (_25253_, _23700_, _25252_);
  nor (_25254_, _25253_, _25251_);
  nand (_25255_, _25254_, _25250_);
  nor (_25256_, _25255_, _25248_);
  and (_25257_, _25256_, _25247_);
  nand (_25258_, _25257_, _25244_);
  and (_25259_, _25258_, _25228_);
  nor (_25260_, _25259_, _25234_);
  and (_25261_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_25262_, _23742_, _23454_);
  nor (_25263_, _23796_, _25236_);
  nand (_25264_, _25263_, _23710_);
  or (_25265_, _25263_, _23710_);
  and (_25266_, _25265_, _23744_);
  and (_25267_, _25266_, _25264_);
  nor (_25268_, _25267_, _25262_);
  and (_25269_, _25245_, _23448_);
  and (_25270_, _23705_, _23487_);
  nor (_25271_, _23736_, _23486_);
  not (_25272_, _25271_);
  and (_25273_, _23691_, _23455_);
  and (_25274_, _23700_, _24859_);
  nor (_25275_, _25274_, _25273_);
  nand (_25276_, _25275_, _25272_);
  or (_25277_, _25276_, _25270_);
  nor (_25278_, _25277_, _25269_);
  and (_25279_, _25278_, _25268_);
  nor (_25280_, _25279_, _25230_);
  nor (_25281_, _25280_, _25261_);
  or (_25282_, _25228_, _23159_);
  not (_25283_, _23761_);
  nand (_25284_, _25228_, _25283_);
  and (_25285_, _25284_, _25282_);
  and (_25286_, _25285_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_25287_, _25286_, _25281_);
  and (_25288_, _25287_, _25260_);
  and (_25289_, _25288_, _25233_);
  nor (_25290_, _25288_, _25233_);
  nor (_25291_, _25290_, _25289_);
  nor (_25292_, _25291_, _23072_);
  nor (_25293_, _25292_, _23144_);
  nor (_25294_, _25293_, _25228_);
  nor (_25295_, _25294_, _25231_);
  nor (_25296_, _25295_, _25222_);
  not (_25297_, _25162_);
  and (_25298_, _25216_, _25123_);
  and (_25299_, _25298_, _25297_);
  nor (_25300_, _25299_, _25296_);
  and (_25301_, _25300_, _25219_);
  nor (_25302_, _25301_, _23153_);
  and (_25303_, _25301_, _23153_);
  nor (_25304_, _25303_, _25302_);
  not (_25305_, _25304_);
  and (_25306_, _25027_, _23669_);
  nor (_25307_, _25306_, _23536_);
  or (_25308_, _25307_, _25026_);
  and (_25309_, _25308_, _23570_);
  not (_25310_, _25309_);
  not (_25311_, _23744_);
  nor (_25312_, _25308_, _23570_);
  nor (_25313_, _25312_, _25311_);
  and (_25314_, _25313_, _25310_);
  nor (_25316_, _23576_, _23536_);
  not (_25317_, _25316_);
  nor (_25318_, _25020_, _23677_);
  and (_25319_, _25318_, _25317_);
  nor (_25320_, _25319_, _25314_);
  and (_25322_, _23691_, _23578_);
  and (_25323_, _23700_, _23570_);
  nor (_25324_, _25323_, _25322_);
  nor (_25325_, _23811_, _23570_);
  and (_25326_, _23705_, _23580_);
  nor (_25328_, _23736_, _23579_);
  or (_25329_, _25328_, _25326_);
  nor (_25330_, _25329_, _25325_);
  and (_25331_, _25330_, _25324_);
  and (_25332_, _25331_, _25320_);
  nor (_25333_, _25332_, _25230_);
  and (_25334_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_25335_, _25230_, _23824_);
  nor (_25336_, _25335_, _25334_);
  and (_25337_, _25336_, _25289_);
  and (_25338_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_25339_, _23536_, _23316_);
  nor (_25340_, _23536_, _23607_);
  nor (_25341_, _25340_, _25339_);
  nor (_25342_, _25341_, _25020_);
  nor (_25343_, _25027_, _23536_);
  not (_25344_, _25343_);
  or (_25345_, _25024_, _23710_);
  and (_25346_, _25345_, _25344_);
  and (_25347_, _25346_, _23316_);
  or (_25348_, _25346_, _23316_);
  nand (_25349_, _25348_, _23744_);
  nor (_25350_, _25349_, _25347_);
  nor (_25351_, _25350_, _25342_);
  nor (_25352_, _23736_, _23324_);
  and (_25353_, _23705_, _23325_);
  nor (_25354_, _25353_, _25352_);
  and (_25355_, _23691_, _23323_);
  and (_25356_, _23700_, _23669_);
  nor (_25357_, _25356_, _25355_);
  and (_25358_, _25245_, _23316_);
  not (_25359_, _25358_);
  and (_25360_, _25359_, _25357_);
  and (_25361_, _25360_, _25354_);
  and (_25362_, _25361_, _25351_);
  nor (_25363_, _25362_, _25230_);
  nor (_25364_, _25363_, _25338_);
  and (_25365_, _25364_, _25337_);
  and (_25366_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_25367_, _25366_, _25333_);
  and (_25368_, _25367_, _25365_);
  nor (_25369_, _25367_, _25365_);
  nor (_25370_, _25369_, _25368_);
  nor (_25371_, _25370_, _23072_);
  nor (_25372_, _25371_, _23175_);
  nor (_25373_, _25372_, _25228_);
  nor (_25374_, _25373_, _25333_);
  nor (_25375_, _25374_, _25222_);
  not (_25376_, _25375_);
  and (_25377_, _25196_, _25332_);
  and (_25378_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_25379_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_25380_, _25379_, _25378_);
  and (_25381_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_25382_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_25383_, _25382_, _25381_);
  and (_25384_, _25383_, _25380_);
  and (_25385_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_25386_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_25387_, _25386_, _25385_);
  and (_25388_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_25389_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_25390_, _25389_, _25388_);
  and (_25391_, _25390_, _25387_);
  and (_25392_, _25391_, _25197_);
  and (_25393_, _25392_, _25384_);
  nor (_25394_, _25393_, _25377_);
  and (_25395_, _25394_, _25125_);
  not (_25396_, _24262_);
  and (_25397_, _25217_, _25396_);
  nor (_25398_, _25124_, _23065_);
  nor (_25399_, _25398_, _25397_);
  not (_25400_, _25399_);
  nor (_25401_, _25400_, _25395_);
  and (_25402_, _25401_, _25376_);
  nor (_25403_, _25402_, _23183_);
  and (_25404_, _25402_, _23183_);
  nor (_25405_, _25404_, _25403_);
  and (_25406_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_25407_, _25406_, _25368_);
  or (_25408_, _25406_, _25368_);
  and (_25409_, _25408_, _23111_);
  nand (_25410_, _25409_, _25407_);
  nor (_25411_, _25228_, _23082_);
  and (_25412_, _25411_, _25410_);
  nor (_25413_, _23811_, _23279_);
  not (_25414_, _25413_);
  and (_25415_, _25414_, _25013_);
  and (_25416_, _25415_, _25006_);
  and (_25417_, _25416_, _25036_);
  and (_25418_, _25417_, _25228_);
  nor (_25419_, _25418_, _25412_);
  nand (_25420_, _25419_, _25220_);
  and (_25421_, _25417_, _25196_);
  and (_25422_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_25423_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_25424_, _25423_, _25422_);
  and (_25425_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_25426_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_25427_, _25426_, _25425_);
  and (_25428_, _25427_, _25424_);
  nand (_25429_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_25430_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_25431_, _25430_, _25429_);
  nand (_25432_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_25433_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_25434_, _25433_, _25432_);
  and (_25435_, _25434_, _25431_);
  and (_25436_, _25435_, _25197_);
  and (_25437_, _25436_, _25428_);
  nor (_25438_, _25437_, _25421_);
  nand (_25439_, _25438_, _25124_);
  not (_25440_, _24222_);
  and (_25441_, _25215_, _23048_);
  nand (_25442_, _25441_, _25440_);
  and (_25443_, _25442_, _23065_);
  and (_25444_, _25443_, _25439_);
  nand (_25445_, _25444_, _25420_);
  and (_25446_, _25445_, _23226_);
  nor (_25447_, _25445_, _23226_);
  nor (_25448_, _25447_, _25446_);
  nor (_25449_, _25448_, _25405_);
  nor (_25450_, _25336_, _25289_);
  nor (_25451_, _25450_, _25337_);
  nor (_25452_, _25451_, _23072_);
  nor (_25453_, _25452_, _23113_);
  nor (_25454_, _25453_, _25228_);
  nor (_25455_, _25454_, _25335_);
  nor (_25456_, _25455_, _25222_);
  not (_25457_, _25456_);
  and (_25458_, _25196_, _23824_);
  and (_25459_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_25460_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_25461_, _25460_, _25459_);
  and (_25462_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_25463_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_25464_, _25463_, _25462_);
  and (_25465_, _25464_, _25461_);
  and (_25466_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_25467_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_25468_, _25467_, _25466_);
  and (_25469_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_25470_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_25471_, _25470_, _25469_);
  and (_25472_, _25471_, _25468_);
  and (_25473_, _25472_, _25197_);
  and (_25474_, _25473_, _25465_);
  nor (_25475_, _25474_, _25458_);
  and (_25476_, _25475_, _25125_);
  and (_25477_, _25298_, _25140_);
  not (_25478_, _25477_);
  or (_25479_, _24340_, _25123_);
  and (_25481_, _25479_, _23065_);
  or (_25482_, _25481_, _25058_);
  nand (_25483_, _25482_, _25478_);
  nor (_25484_, _25483_, _25476_);
  and (_25485_, _25484_, _25457_);
  nor (_25486_, _25485_, _23122_);
  and (_25487_, _25485_, _23122_);
  nor (_25488_, _25487_, _25486_);
  not (_25489_, _25441_);
  and (_25490_, _25398_, _25489_);
  not (_25491_, _25490_);
  nor (_25492_, _25364_, _25337_);
  nor (_25493_, _25492_, _25365_);
  nor (_25494_, _25493_, _23072_);
  nor (_25495_, _25494_, _23193_);
  nor (_25496_, _25495_, _25228_);
  nor (_25497_, _25496_, _25363_);
  nor (_25498_, _25497_, _25222_);
  not (_25499_, _25498_);
  and (_25500_, _25196_, _25362_);
  and (_25502_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_25503_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_25504_, _25503_, _25502_);
  and (_25505_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_25506_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_25507_, _25506_, _25505_);
  and (_25508_, _25507_, _25504_);
  and (_25509_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_25510_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_25511_, _25510_, _25509_);
  and (_25512_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_25513_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_25514_, _25513_, _25512_);
  and (_25515_, _25514_, _25511_);
  and (_25516_, _25515_, _25197_);
  and (_25517_, _25516_, _25508_);
  nor (_25518_, _25517_, _25500_);
  and (_25519_, _25518_, _25125_);
  not (_25520_, _24301_);
  and (_25521_, _25217_, _25520_);
  nor (_25523_, _25521_, _25519_);
  and (_25524_, _25523_, _25499_);
  and (_25525_, _25524_, _25491_);
  nor (_25526_, _25525_, _23201_);
  and (_25528_, _25525_, _23201_);
  nor (_25529_, _25528_, _25526_);
  nor (_25530_, _25529_, _25488_);
  and (_25531_, _25530_, _25449_);
  and (_25532_, _25531_, _25305_);
  not (_25533_, _25128_);
  not (_25534_, _23215_);
  nor (_25535_, _23167_, _23137_);
  and (_25536_, _25535_, _25534_);
  nor (_25537_, _25536_, _25533_);
  and (_25538_, _25537_, _25532_);
  and (_25539_, _25538_, _25057_);
  not (_25540_, _25539_);
  or (_25541_, _24162_, _22985_);
  nor (_25542_, _23652_, _23357_);
  and (_25543_, _23652_, _23357_);
  nor (_25544_, _25543_, _25542_);
  not (_25545_, _25544_);
  nor (_25547_, _23654_, _23617_);
  nor (_25548_, _25547_, _23655_);
  and (_25549_, _25548_, _25545_);
  nor (_25550_, _25057_, _23057_);
  nor (_25551_, _23653_, _23620_);
  nor (_25552_, _25551_, _23654_);
  and (_25553_, _23645_, _23633_);
  nor (_25554_, _25553_, _23646_);
  and (_25555_, _23540_, _23536_);
  nor (_25556_, _25555_, _23541_);
  not (_25557_, _25556_);
  nor (_25558_, _23643_, _23636_);
  nor (_25559_, _25558_, _23644_);
  and (_25560_, _25559_, _25557_);
  and (_25561_, _25560_, _25554_);
  and (_25562_, _25561_, _23640_);
  and (_25563_, _25562_, _25552_);
  nand (_25564_, _25563_, _25550_);
  nor (_25565_, _25564_, _24997_);
  and (_25566_, _25565_, _25549_);
  not (_25567_, _25566_);
  and (_25568_, _25057_, _23685_);
  not (_25569_, _25568_);
  nor (_25570_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_25571_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_25572_, _25571_, _25570_);
  nor (_25573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_25574_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_25575_, _25574_, _25573_);
  and (_25576_, _25575_, _25572_);
  and (_25577_, _25576_, _22946_);
  nor (_25578_, _24149_, _22980_);
  nor (_25579_, _25578_, _23058_);
  and (_25580_, _25579_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25581_, _25580_, _25577_);
  and (_25582_, _25581_, _25569_);
  and (_25583_, _25582_, _25567_);
  and (_25584_, _22992_, _22972_);
  or (_25585_, _25584_, _22994_);
  or (_25586_, _25585_, _22984_);
  and (_25587_, _25586_, _22862_);
  not (_25588_, _25587_);
  nor (_25589_, _24165_, _24156_);
  and (_25590_, _25589_, _24145_);
  and (_25591_, _25590_, _25588_);
  and (_25592_, _25591_, _25583_);
  and (_25593_, _24138_, _22973_);
  and (_25594_, _23056_, _22973_);
  or (_25595_, _25594_, _24148_);
  or (_25596_, _25595_, _25593_);
  nor (_25597_, _25596_, _25583_);
  nor (_25598_, _25597_, _25592_);
  nor (_25599_, _25598_, _25541_);
  and (_25600_, _25599_, _23029_);
  nor (_25601_, _23043_, _22944_);
  nor (_25602_, _25601_, _25600_);
  nor (_25603_, _25602_, _24178_);
  not (_25604_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_25605_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _22734_);
  and (_25606_, _25605_, _25604_);
  not (_25607_, _25606_);
  not (_25608_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_25609_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22734_);
  and (_25610_, _25609_, _25608_);
  and (_25611_, _23202_, _23122_);
  and (_25612_, _25611_, _25133_);
  nor (_25613_, _25612_, _25610_);
  and (_25614_, _25613_, _25607_);
  nor (_25615_, _23154_, _23098_);
  and (_25616_, _25615_, _23122_);
  nor (_25617_, _23201_, _23183_);
  and (_25618_, _25127_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_25619_, _25618_, _25617_);
  and (_25620_, _25619_, _25616_);
  not (_25621_, _25620_);
  and (_25622_, _25621_, _25614_);
  not (_25623_, _25622_);
  and (_25624_, _25623_, _22946_);
  nor (_25625_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_25626_, _25625_);
  and (_25627_, _25615_, _23123_);
  nand (_25628_, _25618_, _23201_);
  nor (_25629_, _25628_, _23183_);
  and (_25630_, _25629_, _25627_);
  nor (_25631_, _25630_, _25626_);
  and (_25632_, _25631_, _25136_);
  not (_25633_, _25632_);
  and (_25634_, _25633_, _25579_);
  or (_25635_, _25634_, _25624_);
  nor (_25636_, _25635_, _25603_);
  not (_25637_, _25532_);
  and (_25638_, _25196_, _23761_);
  and (_25639_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_25640_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_25641_, _25640_, _25639_);
  and (_25642_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_25643_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_25644_, _25643_, _25642_);
  and (_25645_, _25644_, _25641_);
  and (_25646_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_25647_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_25648_, _25647_, _25646_);
  and (_25649_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_25650_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_25651_, _25650_, _25649_);
  and (_25652_, _25651_, _25648_);
  and (_25653_, _25652_, _25197_);
  and (_25654_, _25653_, _25645_);
  nor (_25655_, _25654_, _25638_);
  and (_25656_, _25655_, _25125_);
  not (_25657_, _25656_);
  and (_25658_, _25298_, _22835_);
  nor (_25659_, _25285_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_25660_, _25659_, _25286_);
  nor (_25661_, _25660_, _23072_);
  nor (_25662_, _25661_, _23160_);
  nor (_25663_, _25662_, _25228_);
  not (_25664_, _25663_);
  and (_25665_, _25664_, _25284_);
  not (_25666_, _25665_);
  nand (_25667_, _25666_, _25221_);
  nand (_25668_, _25217_, _24499_);
  nand (_25669_, _25668_, _25667_);
  nor (_25670_, _25669_, _25658_);
  and (_25671_, _25670_, _25657_);
  and (_25672_, _25671_, _25181_);
  not (_25673_, _25672_);
  nor (_25674_, _25197_, _25258_);
  and (_25675_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_25677_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_25678_, _25677_, _25675_);
  and (_25679_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_25680_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_25681_, _25680_, _25679_);
  and (_25682_, _25681_, _25678_);
  and (_25683_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_25684_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_25685_, _25684_, _25683_);
  and (_25686_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_25687_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_25688_, _25687_, _25686_);
  and (_25689_, _25688_, _25685_);
  and (_25691_, _25689_, _25197_);
  and (_25692_, _25691_, _25682_);
  nor (_25693_, _25692_, _25674_);
  and (_25694_, _25693_, _25125_);
  and (_25695_, _25217_, _24418_);
  nor (_25696_, _25695_, _25694_);
  nor (_25697_, _25287_, _25260_);
  nor (_25698_, _25697_, _25288_);
  nor (_25699_, _25698_, _23072_);
  nor (_25700_, _25699_, _23207_);
  nor (_25701_, _25700_, _25228_);
  nor (_25702_, _25701_, _25259_);
  not (_25703_, _25702_);
  and (_25704_, _25703_, _25221_);
  and (_25705_, _25298_, _22782_);
  nor (_25706_, _25705_, _25704_);
  and (_25707_, _25706_, _25696_);
  and (_25708_, _25707_, _25534_);
  nor (_25709_, _25707_, _25534_);
  nor (_25710_, _25709_, _25708_);
  nand (_25711_, _25710_, _25673_);
  not (_25712_, _23137_);
  and (_25713_, _25217_, _24457_);
  nor (_25714_, _25286_, _25281_);
  nor (_25715_, _25714_, _25287_);
  nor (_25716_, _25715_, _23072_);
  nor (_25717_, _25716_, _23127_);
  nor (_25718_, _25717_, _25228_);
  nor (_25719_, _25718_, _25280_);
  not (_25720_, _25719_);
  nand (_25721_, _25720_, _25220_);
  and (_25722_, _25721_, _23065_);
  nor (_25723_, _25722_, _25398_);
  and (_25724_, _25196_, _25279_);
  and (_25725_, _25198_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_25727_, _25203_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_25728_, _25727_, _25725_);
  and (_25729_, _25164_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_25730_, _25205_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_25731_, _25730_, _25729_);
  and (_25732_, _25731_, _25728_);
  and (_25733_, _25171_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_25734_, _25167_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_25735_, _25734_, _25733_);
  and (_25736_, _25200_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_25737_, _25174_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_25738_, _25737_, _25736_);
  and (_25739_, _25738_, _25735_);
  and (_25740_, _25739_, _25197_);
  and (_25741_, _25740_, _25732_);
  nor (_25742_, _25741_, _25724_);
  and (_25743_, _25742_, _25125_);
  and (_25744_, _25298_, _22947_);
  or (_25745_, _25744_, _25743_);
  or (_25746_, _25745_, _25723_);
  nor (_25748_, _25746_, _25713_);
  and (_25749_, _25748_, _25712_);
  nor (_25750_, _25748_, _25712_);
  not (_25751_, _25127_);
  nor (_25752_, _25671_, _25181_);
  or (_25753_, _25752_, _25751_);
  or (_25754_, _25753_, _25750_);
  or (_25755_, _25754_, _25749_);
  or (_25756_, _25755_, _25711_);
  nor (_25757_, _25756_, _25637_);
  nor (_25758_, _23098_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_25759_, _25758_, _25757_);
  not (_25760_, _25759_);
  and (_25761_, _25760_, _25636_);
  and (_25762_, _25761_, _25540_);
  and (_25763_, _23711_, _23603_);
  and (_25764_, _23715_, _23795_);
  nor (_25766_, _23570_, _23279_);
  and (_25767_, _25766_, _23316_);
  and (_25768_, _25767_, _25024_);
  and (_25769_, _25768_, _23483_);
  and (_25770_, _25769_, _23454_);
  and (_25771_, _25770_, _23419_);
  and (_25772_, _23536_, _23647_);
  and (_25773_, _25772_, _25771_);
  nor (_25774_, _23536_, _23322_);
  and (_25775_, _25028_, _23279_);
  and (_25776_, _23628_, _23384_);
  nor (_25777_, _23483_, _23454_);
  and (_25778_, _25777_, _25776_);
  and (_25779_, _25778_, _25775_);
  and (_25780_, _25779_, _23354_);
  and (_25781_, _25780_, _25774_);
  or (_25782_, _25781_, _25773_);
  and (_25783_, _23536_, _23607_);
  and (_25784_, _23536_, _23354_);
  nor (_25785_, _25784_, _25783_);
  and (_25786_, _25785_, _25782_);
  nor (_25787_, _23577_, _23536_);
  and (_25788_, _23577_, _23536_);
  nor (_25789_, _25788_, _25787_);
  and (_25790_, _25789_, _25786_);
  nor (_25791_, _25790_, _23603_);
  and (_25792_, _25790_, _23603_);
  nor (_25793_, _25792_, _25791_);
  and (_25794_, _25793_, _23744_);
  and (_25795_, _23536_, _23603_);
  nor (_25796_, _25795_, _23674_);
  nor (_25797_, _25796_, _25020_);
  or (_25798_, _25797_, _25794_);
  or (_25799_, _25798_, _25764_);
  and (_25800_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_25801_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25802_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24536_);
  nor (_25803_, _25802_, _25801_);
  not (_25804_, _25803_);
  nor (_25805_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25806_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24538_);
  nor (_25807_, _25806_, _25805_);
  nor (_25808_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25809_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24541_);
  nor (_25810_, _25809_, _25808_);
  and (_25811_, _25810_, _23594_);
  nor (_25812_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25813_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24540_);
  nor (_25814_, _25813_, _25812_);
  and (_25815_, _25814_, _25811_);
  nor (_25816_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25817_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24539_);
  nor (_25818_, _25817_, _25816_);
  and (_25819_, _25818_, _25815_);
  and (_25820_, _25819_, _25807_);
  nor (_25821_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25822_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24537_);
  nor (_25824_, _25822_, _25821_);
  nand (_25825_, _25824_, _25820_);
  or (_25826_, _25825_, _25804_);
  nor (_25827_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_25828_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _24535_);
  nor (_25829_, _25828_, _25827_);
  not (_25830_, _25829_);
  or (_25831_, _25830_, _25826_);
  nor (_25832_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_25833_, _24184_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_25834_, _25833_, _25832_);
  nor (_25835_, _25834_, _25831_);
  and (_25836_, _25834_, _25831_);
  or (_25837_, _25836_, _25835_);
  nand (_25838_, _25837_, _23238_);
  or (_25839_, _24974_, _24936_);
  and (_25840_, _25839_, _24975_);
  and (_25841_, _25840_, _24794_);
  not (_25842_, _25841_);
  nand (_25843_, _25842_, _25838_);
  or (_25844_, _25843_, _25800_);
  or (_25845_, _25844_, _25799_);
  or (_25846_, _25845_, _25763_);
  and (_25847_, _25846_, _24179_);
  and (_25848_, _25440_, _24172_);
  and (_25849_, _24170_, _24174_);
  and (_25850_, _25849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_25851_, _25850_, _25848_);
  nor (_25852_, _25851_, _25847_);
  nand (_25853_, _25852_, _25762_);
  or (_25854_, _25853_, _25055_);
  or (_25855_, _25854_, _24555_);
  and (_25856_, _22745_, _22748_);
  nor (_25857_, _25856_, _24307_);
  nor (_25858_, _25857_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_25859_, _25858_);
  and (_25860_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_25861_, _25860_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_25862_, _25861_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_25863_, _25862_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_25864_, _25863_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_25865_, _25864_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_25866_, _25865_, _25859_);
  and (_25867_, _25866_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_25868_, _25867_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_25869_, _25868_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_25870_, _25869_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_25871_, _25870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_25872_, _25871_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_25873_, _25872_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_25874_, _25872_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_25875_, _25874_, _25873_);
  or (_25876_, _25875_, _25762_);
  and (_25877_, _25876_, _23049_);
  and (_26921_[15], _25877_, _25855_);
  and (_26920_, _23049_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r );
  nor (_25878_, _23043_, rst);
  and (_26919_, _25878_, _25762_);
  and (_26918_[7], _25438_, _23049_);
  nor (_26917_[4], _25139_, rst);
  and (_26916_, _25445_, _23049_);
  and (_25879_, _23731_, _23512_);
  and (_25880_, _25879_, _23730_);
  nor (_25881_, _25160_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_25882_, _23519_, _23763_);
  and (_25883_, _25882_, _23369_);
  or (_25884_, _25883_, _25881_);
  or (_25885_, _25884_, _25880_);
  and (_25886_, _25885_, _23100_);
  and (_25887_, _25886_, _23849_);
  and (_25888_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_19750_, _25888_, _25887_);
  and (_25889_, _23154_, _23122_);
  and (_25890_, _25889_, _23226_);
  and (_25891_, _25890_, _25629_);
  and (_25892_, _23167_, _25712_);
  and (_25894_, _25892_, _23215_);
  not (_25895_, _25894_);
  nor (_25896_, _25895_, _23729_);
  and (_25897_, _25223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_25898_, _25897_, _25896_);
  and (_25899_, _25898_, _25891_);
  and (_25900_, _25126_, _25225_);
  nor (_25901_, _25533_, _23153_);
  and (_25902_, _25901_, _25131_);
  and (_25903_, _25902_, _25900_);
  or (_25904_, _25535_, _25534_);
  not (_25905_, _25904_);
  nand (_25906_, _25905_, _25891_);
  and (_25907_, _25906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_25908_, _25907_, _25903_);
  or (_25909_, _25908_, _25899_);
  not (_25910_, _25903_);
  or (_25911_, _25910_, _25258_);
  and (_25912_, _25911_, _23049_);
  and (_22232_, _25912_, _25909_);
  nor (_25913_, _23772_, _23140_);
  and (_25914_, _25913_, _23774_);
  and (_25915_, _25914_, _23779_);
  not (_25916_, _25915_);
  and (_25917_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nand (_25918_, _23731_, _23498_);
  nor (_25919_, _25918_, _23729_);
  nor (_25920_, _25279_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_25921_, _25879_, _23784_);
  and (_25922_, _23731_, _23502_);
  or (_25923_, _25922_, _25921_);
  and (_25924_, _25923_, _23438_);
  or (_25925_, _25924_, _25920_);
  or (_25926_, _25925_, _25919_);
  and (_25927_, _25926_, _23100_);
  and (_25928_, _25927_, _25915_);
  or (_22597_, _25928_, _25917_);
  and (_25930_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_25931_, _25915_, _23768_);
  or (_22601_, _25931_, _25930_);
  and (_25932_, _25913_, _23219_);
  not (_25933_, _23221_);
  nor (_25934_, _23202_, _23102_);
  not (_25935_, _25934_);
  and (_25936_, _25935_, _23100_);
  and (_25937_, _25936_, _25933_);
  and (_25938_, _25937_, _23229_);
  and (_25939_, _25938_, _25932_);
  and (_25940_, _25939_, _23768_);
  not (_25941_, _25939_);
  and (_25942_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_22671_, _25942_, _25940_);
  and (_25943_, _22740_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_25944_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_25945_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_25946_, _25943_, _25945_);
  or (_25947_, _25946_, _25944_);
  and (_26914_[0], _25947_, _23049_);
  and (_25948_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_25949_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_25950_, _25943_, _25949_);
  or (_25951_, _25950_, _25948_);
  and (_26914_[1], _25951_, _23049_);
  and (_25952_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_25953_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_25955_, _25943_, _25953_);
  or (_25956_, _25955_, _25952_);
  and (_26914_[2], _25956_, _23049_);
  and (_25957_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_25958_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_25959_, _25943_, _25958_);
  or (_25960_, _25959_, _25957_);
  and (_26914_[3], _25960_, _23049_);
  and (_25961_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_25962_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_25963_, _25943_, _25962_);
  or (_25964_, _25963_, _25961_);
  and (_26914_[4], _25964_, _23049_);
  and (_25965_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_25966_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_25967_, _25943_, _25966_);
  or (_25969_, _25967_, _25965_);
  and (_26914_[5], _25969_, _23049_);
  and (_25970_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_25971_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_25972_, _25943_, _25971_);
  or (_25973_, _25972_, _25970_);
  and (_26914_[6], _25973_, _23049_);
  and (_25974_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_25976_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_25977_, _25943_, _25976_);
  or (_25978_, _25977_, _25974_);
  and (_26914_[7], _25978_, _23049_);
  and (_25979_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_25981_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_25982_, _25943_, _25981_);
  or (_25983_, _25982_, _25979_);
  and (_26914_[8], _25983_, _23049_);
  and (_25984_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_25985_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_25987_, _25943_, _25985_);
  or (_25988_, _25987_, _25984_);
  and (_26914_[9], _25988_, _23049_);
  and (_25989_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_25990_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_25991_, _25943_, _25990_);
  or (_25992_, _25991_, _25989_);
  and (_26914_[10], _25992_, _23049_);
  and (_25994_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_25996_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_25997_, _25943_, _25996_);
  or (_25998_, _25997_, _25994_);
  and (_26914_[11], _25998_, _23049_);
  and (_25999_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_26001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_26002_, _25943_, _26001_);
  or (_26003_, _26002_, _25999_);
  and (_26914_[12], _26003_, _23049_);
  and (_26004_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_26005_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_26006_, _25943_, _26005_);
  or (_26007_, _26006_, _26004_);
  and (_26914_[13], _26007_, _23049_);
  and (_26008_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_26009_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_26010_, _25943_, _26009_);
  or (_26011_, _26010_, _26008_);
  and (_26914_[14], _26011_, _23049_);
  and (_26012_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_26013_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_26014_, _25943_, _26013_);
  or (_26015_, _26014_, _26012_);
  and (_26915_[0], _26015_, _23049_);
  and (_26016_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_26017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_26018_, _25943_, _26017_);
  or (_26019_, _26018_, _26016_);
  and (_26915_[1], _26019_, _23049_);
  and (_26020_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_26021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_26022_, _25943_, _26021_);
  or (_26023_, _26022_, _26020_);
  and (_26915_[2], _26023_, _23049_);
  and (_26024_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_26025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_26026_, _25943_, _26025_);
  or (_26027_, _26026_, _26024_);
  and (_26915_[3], _26027_, _23049_);
  or (_26028_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_26029_, _25943_, _25962_);
  and (_26030_, _26029_, _23049_);
  and (_26915_[4], _26030_, _26028_);
  and (_26031_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_26032_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_26033_, _25943_, _26032_);
  or (_26034_, _26033_, _26031_);
  and (_26915_[5], _26034_, _23049_);
  and (_26035_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_26036_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_26037_, _25943_, _26036_);
  or (_26038_, _26037_, _26035_);
  and (_26915_[6], _26038_, _23049_);
  and (_26039_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_26040_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_26041_, _25943_, _26040_);
  or (_26042_, _26041_, _26039_);
  and (_26915_[7], _26042_, _23049_);
  or (_26044_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand (_26045_, _25943_, _25981_);
  and (_26046_, _26045_, _23049_);
  and (_26915_[8], _26046_, _26044_);
  and (_26047_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_26048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_26049_, _25943_, _26048_);
  or (_26050_, _26049_, _26047_);
  and (_26915_[9], _26050_, _23049_);
  and (_26051_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not (_26052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_26053_, _25943_, _26052_);
  or (_26054_, _26053_, _26051_);
  and (_26915_[10], _26054_, _23049_);
  and (_26055_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_26056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_26057_, _25943_, _26056_);
  or (_26058_, _26057_, _26055_);
  and (_26915_[11], _26058_, _23049_);
  or (_26059_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand (_26060_, _25943_, _26001_);
  and (_26061_, _26060_, _23049_);
  and (_26915_[12], _26061_, _26059_);
  and (_26062_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_26063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_26065_, _25943_, _26063_);
  or (_26066_, _26065_, _26062_);
  and (_26915_[13], _26066_, _23049_);
  and (_26067_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not (_26068_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_26069_, _25943_, _26068_);
  or (_26070_, _26069_, _26067_);
  and (_26915_[14], _26070_, _23049_);
  and (_26071_, _23772_, _23139_);
  and (_26072_, _26071_, _23219_);
  and (_26073_, _26072_, _23230_);
  and (_26074_, _26073_, _25886_);
  not (_26075_, _26073_);
  and (_26076_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_23781_, _26076_, _26074_);
  nand (_26077_, _23784_, _23498_);
  nor (_26078_, _26077_, _23729_);
  nor (_26079_, _25362_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_26080_, _23498_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26081_, _23305_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_26082_, _26081_, _26080_);
  or (_26083_, _26082_, _26079_);
  or (_26084_, _26083_, _26078_);
  and (_26085_, _26084_, _23100_);
  and (_26086_, _26085_, _26073_);
  and (_26087_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_24045_, _26087_, _26086_);
  not (_26088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor (_26089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_26090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_26092_, _26090_, _26089_);
  and (_26093_, _26092_, _26088_);
  and (_26094_, _26093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  not (_26095_, _26093_);
  and (_26096_, _26089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_26097_, _26096_);
  and (_26098_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_26099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_26100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_26102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _26100_);
  and (_26103_, _26102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_26104_, _26103_, _26099_);
  and (_26105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_26106_, _26105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_26107_, _26106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_26108_, _26107_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_26109_, _26108_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_26110_, _26109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_26111_, _26110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_26112_, _26111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_26113_, _26112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_26114_, _26113_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_26115_, _26114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_26116_, _26115_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_26117_, _26116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_26118_, _26117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_26119_, _26118_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_26120_, _26119_, _26104_);
  and (_26121_, _26120_, _26098_);
  and (_26122_, _26105_, _26104_);
  or (_26123_, _26122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_26124_, _26106_, _26104_);
  and (_26125_, _26124_, _26123_);
  or (_26126_, _26125_, _26121_);
  and (_26127_, _26126_, _26095_);
  or (_26128_, _26127_, _26094_);
  and (_26130_, _25130_, _25534_);
  and (_26131_, _25901_, _26130_);
  and (_26132_, _26131_, _25900_);
  not (_26133_, _26132_);
  and (_26134_, _26133_, _26128_);
  and (_26136_, _25182_, _25534_);
  and (_26137_, _25901_, _26136_);
  and (_26138_, _26137_, _25900_);
  and (_26139_, _26132_, _25258_);
  or (_26140_, _26139_, _26138_);
  or (_26141_, _26140_, _26134_);
  not (_26142_, _26138_);
  or (_26143_, _26142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_26144_, _26143_, _23049_);
  and (_24066_, _26144_, _26141_);
  and (_26145_, _26073_, _23830_);
  and (_26146_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_24246_, _26146_, _26145_);
  and (_26147_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_26148_, _25915_, _23830_);
  or (_27060_, _26148_, _26147_);
  and (_26149_, _23217_, _23189_);
  and (_26150_, _26149_, _26071_);
  and (_26151_, _26150_, _25938_);
  and (_26152_, _26151_, _23830_);
  not (_26153_, _26151_);
  and (_26154_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_25054_, _26154_, _26152_);
  and (_26156_, _26151_, _25886_);
  and (_26157_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_27246_, _26157_, _26156_);
  and (_26158_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_26159_, _25915_, _25886_);
  or (_25480_, _26159_, _26158_);
  and (_26160_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nand (_26161_, _23731_, _23503_);
  nor (_26162_, _26161_, _23729_);
  and (_26163_, _25258_, _23763_);
  and (_26164_, _23731_, _23497_);
  or (_26165_, _26164_, _25921_);
  and (_26166_, _26165_, _23400_);
  or (_26167_, _26166_, _26163_);
  or (_26168_, _26167_, _26162_);
  and (_26170_, _26168_, _23100_);
  and (_26171_, _26170_, _25915_);
  or (_25501_, _26171_, _26160_);
  and (_26172_, _26151_, _26085_);
  and (_26173_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_25522_, _26173_, _26172_);
  and (_26174_, _23225_, _23098_);
  and (_26175_, _26174_, _25937_);
  and (_26176_, _26175_, _23220_);
  nand (_26177_, _23784_, _23503_);
  nor (_26178_, _26177_, _23729_);
  nor (_26179_, _25332_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_26180_, _23503_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26181_, _23506_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_26182_, _26181_, _26180_);
  or (_26183_, _26182_, _26179_);
  or (_26184_, _26183_, _26178_);
  and (_26185_, _26184_, _23100_);
  and (_26186_, _26185_, _26176_);
  not (_26188_, _26176_);
  and (_26189_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_26330_, _26189_, _26186_);
  and (_26190_, _26071_, _23774_);
  nor (_26191_, _25936_, _23222_);
  and (_26192_, _25126_, _23100_);
  and (_26193_, _26192_, _26191_);
  and (_26194_, _26193_, _26190_);
  and (_26195_, _26194_, _23830_);
  not (_26196_, _26194_);
  and (_26197_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_26358_, _26197_, _26195_);
  and (_26198_, _26176_, _26085_);
  and (_26199_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_26396_, _26199_, _26198_);
  and (_26200_, _26194_, _25886_);
  and (_26201_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or (_27104_, _26201_, _26200_);
  and (_26202_, _23773_, _23219_);
  and (_26204_, _25937_, _23777_);
  and (_26205_, _26204_, _26202_);
  not (_26206_, _26205_);
  and (_26207_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_26208_, _26205_, _26085_);
  or (_26490_, _26208_, _26207_);
  and (_26209_, _26151_, _25927_);
  and (_26210_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_26509_, _26210_, _26209_);
  and (_26211_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_26212_, _26205_, _23830_);
  or (_00887_, _26212_, _26211_);
  and (_26213_, _23774_, _23170_);
  and (_26214_, _26213_, _23779_);
  not (_26215_, _26214_);
  and (_26216_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  and (_26217_, _26214_, _25927_);
  or (_00920_, _26217_, _26216_);
  and (_26219_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_26220_, _26205_, _25886_);
  or (_00972_, _26220_, _26219_);
  and (_26221_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_26222_, _26205_, _26170_);
  or (_00992_, _26222_, _26221_);
  and (_26224_, _26149_, _25913_);
  and (_26225_, _26224_, _25938_);
  and (_26227_, _26225_, _26085_);
  not (_26228_, _26225_);
  and (_26230_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_02445_, _26230_, _26227_);
  and (_26231_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_26233_, _23784_, _23512_);
  not (_26234_, _26233_);
  nor (_26235_, _26234_, _23729_);
  nand (_26236_, _25417_, _23763_);
  or (_26237_, _23264_, _23763_);
  and (_26239_, _26237_, _26234_);
  and (_26240_, _26239_, _26236_);
  or (_26241_, _26240_, _26235_);
  and (_26242_, _26241_, _23100_);
  and (_26243_, _26242_, _26205_);
  or (_27059_, _26243_, _26231_);
  and (_26244_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_26245_, _26205_, _26185_);
  or (_02673_, _26245_, _26244_);
  and (_26246_, _26242_, _26225_);
  and (_26247_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_02758_, _26247_, _26246_);
  and (_26248_, _26225_, _26185_);
  and (_26249_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_02810_, _26249_, _26248_);
  and (_26250_, _26225_, _26170_);
  and (_26252_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_03119_, _26252_, _26250_);
  and (_26254_, _26204_, _23220_);
  not (_26255_, _26254_);
  and (_26256_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_26257_, _26254_, _26185_);
  or (_03364_, _26257_, _26256_);
  and (_26258_, _26071_, _23846_);
  and (_26260_, _25937_, _25126_);
  and (_26261_, _26260_, _26258_);
  not (_26262_, _26261_);
  and (_26263_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_26264_, _26261_, _26185_);
  or (_03398_, _26264_, _26263_);
  and (_26265_, _26225_, _23830_);
  and (_26267_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_03458_, _26267_, _26265_);
  and (_26268_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_26269_, _26254_, _26085_);
  or (_03533_, _26269_, _26268_);
  and (_26270_, _26225_, _25886_);
  and (_26271_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_03555_, _26271_, _26270_);
  and (_26273_, _26174_, _23776_);
  and (_26275_, _26273_, _26258_);
  and (_26276_, _26275_, _23768_);
  not (_26277_, _26275_);
  and (_26278_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_03594_, _26278_, _26276_);
  and (_26279_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_26281_, _26254_, _23830_);
  or (_27057_, _26281_, _26279_);
  and (_26283_, _23846_, _23773_);
  and (_26284_, _26283_, _25938_);
  and (_26285_, _26284_, _25886_);
  not (_26286_, _26284_);
  and (_26287_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_04138_, _26287_, _26285_);
  and (_26290_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_26291_, _26205_, _23768_);
  or (_27058_, _26291_, _26290_);
  and (_26292_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_26293_, _26254_, _26242_);
  or (_04739_, _26293_, _26292_);
  and (_26294_, _26273_, _26190_);
  and (_26295_, _26294_, _25927_);
  not (_26296_, _26294_);
  and (_26297_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_04772_, _26297_, _26295_);
  and (_26298_, _26294_, _26170_);
  and (_26299_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_04799_, _26299_, _26298_);
  and (_26301_, _25938_, _23847_);
  and (_26302_, _26301_, _26185_);
  not (_26303_, _26301_);
  and (_26305_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_04935_, _26305_, _26302_);
  and (_26308_, _26072_, _23848_);
  and (_26310_, _26308_, _26185_);
  not (_26311_, _26308_);
  and (_26312_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_05061_, _26312_, _26310_);
  and (_26313_, _26284_, _23768_);
  and (_26314_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_05104_, _26314_, _26313_);
  and (_26315_, _26308_, _26085_);
  and (_26316_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_05137_, _26316_, _26315_);
  and (_26318_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_26320_, _26254_, _23768_);
  or (_05243_, _26320_, _26318_);
  and (_26321_, _26204_, _26072_);
  not (_26322_, _26321_);
  and (_26323_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and (_26324_, _26321_, _26242_);
  or (_05570_, _26324_, _26323_);
  and (_26326_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_26327_, _26321_, _26185_);
  or (_27056_, _26327_, _26326_);
  and (_26329_, _26258_, _23848_);
  and (_26331_, _26329_, _26170_);
  not (_26332_, _26329_);
  and (_26333_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_05627_, _26333_, _26331_);
  and (_26334_, _26284_, _26185_);
  and (_26335_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_05683_, _26335_, _26334_);
  and (_26336_, _26284_, _26085_);
  and (_26337_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_05785_, _26337_, _26336_);
  and (_26338_, _26225_, _23768_);
  and (_26339_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_06031_, _26339_, _26338_);
  and (_26340_, _26149_, _23773_);
  and (_26341_, _26340_, _25938_);
  and (_26343_, _26341_, _26242_);
  not (_26345_, _26341_);
  and (_26346_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_06192_, _26346_, _26343_);
  and (_26348_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_26349_, _26254_, _26170_);
  or (_06294_, _26349_, _26348_);
  and (_26351_, _26202_, _23848_);
  and (_26352_, _26351_, _23830_);
  not (_26353_, _26351_);
  and (_26354_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_06366_, _26354_, _26352_);
  and (_26355_, _26191_, _26174_);
  and (_26356_, _26355_, _23847_);
  and (_26357_, _26356_, _23768_);
  not (_26359_, _26356_);
  and (_26360_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_06398_, _26360_, _26357_);
  and (_26361_, _26329_, _25927_);
  and (_26362_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_06491_, _26362_, _26361_);
  and (_26363_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_26364_, _26254_, _25927_);
  or (_06565_, _26364_, _26363_);
  and (_26366_, _26355_, _26258_);
  and (_26367_, _26366_, _26242_);
  not (_26368_, _26366_);
  and (_26369_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_27288_, _26369_, _26367_);
  and (_26370_, _26190_, _26175_);
  and (_26371_, _26370_, _26242_);
  not (_26372_, _26370_);
  and (_26373_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_07040_, _26373_, _26371_);
  and (_26374_, _25913_, _23846_);
  and (_26375_, _26174_, _23223_);
  and (_26376_, _26375_, _26374_);
  and (_26377_, _26376_, _23830_);
  not (_26378_, _26376_);
  and (_26379_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_07169_, _26379_, _26377_);
  and (_26380_, _26370_, _23830_);
  and (_26381_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_07257_, _26381_, _26380_);
  and (_26382_, _26301_, _25927_);
  and (_26383_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_07318_, _26383_, _26382_);
  and (_26384_, _26370_, _26185_);
  and (_26385_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_07374_, _26385_, _26384_);
  and (_26386_, _26356_, _23830_);
  and (_26387_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_07487_, _26387_, _26386_);
  and (_26388_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_26389_, _26321_, _26170_);
  or (_07513_, _26389_, _26388_);
  and (_26390_, _26356_, _25886_);
  and (_26391_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_07632_, _26391_, _26390_);
  and (_26392_, _26356_, _26170_);
  and (_26393_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_07688_, _26393_, _26392_);
  and (_26394_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_26395_, _26321_, _25927_);
  or (_07707_, _26395_, _26394_);
  and (_26397_, _26366_, _26170_);
  and (_26398_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_08000_, _26398_, _26397_);
  and (_26399_, _26366_, _25927_);
  and (_26400_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_08099_, _26400_, _26399_);
  and (_26401_, _26366_, _23768_);
  and (_26402_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_08200_, _26402_, _26401_);
  and (_26403_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_26404_, _26321_, _23830_);
  or (_08293_, _26404_, _26403_);
  and (_26405_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_26406_, _26321_, _25886_);
  or (_08527_, _26406_, _26405_);
  and (_26407_, _26366_, _26085_);
  and (_26408_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_08569_, _26408_, _26407_);
  and (_26409_, _26366_, _23830_);
  and (_26410_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_08626_, _26410_, _26409_);
  and (_26411_, _26366_, _25886_);
  and (_26412_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_08715_, _26412_, _26411_);
  and (_26413_, _26374_, _23779_);
  not (_26414_, _26413_);
  and (_26415_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_26416_, _26413_, _26085_);
  or (_27070_, _26416_, _26415_);
  and (_26417_, _26204_, _25932_);
  not (_26418_, _26417_);
  and (_26419_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_26420_, _26417_, _23830_);
  or (_09243_, _26420_, _26419_);
  and (_26421_, _26149_, _23170_);
  and (_26422_, _26421_, _23779_);
  not (_26423_, _26422_);
  and (_26424_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_26425_, _26422_, _25886_);
  or (_27082_, _26425_, _26424_);
  and (_26426_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_26427_, _26261_, _26085_);
  or (_09436_, _26427_, _26426_);
  and (_26428_, _26213_, _26175_);
  and (_26429_, _26428_, _23830_);
  not (_26430_, _26428_);
  and (_26431_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_09482_, _26431_, _26429_);
  and (_26432_, _26375_, _26258_);
  and (_26433_, _26432_, _23768_);
  not (_26434_, _26432_);
  and (_26435_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_09520_, _26435_, _26433_);
  and (_26436_, _26428_, _23768_);
  and (_26437_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_09695_, _26437_, _26436_);
  and (_26438_, _26428_, _26170_);
  and (_26439_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_09768_, _26439_, _26438_);
  and (_26440_, _26242_, _26194_);
  and (_26441_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_09875_, _26441_, _26440_);
  and (_26442_, _26175_, _25914_);
  and (_26443_, _26442_, _23830_);
  not (_26444_, _26442_);
  and (_26445_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_09944_, _26445_, _26443_);
  and (_26446_, _26175_, _23775_);
  and (_26447_, _26446_, _25927_);
  not (_26448_, _26446_);
  and (_26449_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_09976_, _26449_, _26447_);
  and (_26450_, _26294_, _26085_);
  and (_26451_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_10181_, _26451_, _26450_);
  and (_26452_, _26428_, _26185_);
  and (_26453_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_10241_, _26453_, _26452_);
  and (_26454_, _26428_, _26085_);
  and (_26455_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_10505_, _26455_, _26454_);
  and (_26456_, _26194_, _26185_);
  and (_26457_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_10743_, _26457_, _26456_);
  and (_26458_, _26355_, _26224_);
  and (_26459_, _26458_, _25927_);
  not (_26460_, _26458_);
  and (_26461_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_10787_, _26461_, _26459_);
  and (_26462_, _26458_, _23768_);
  and (_26463_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_10919_, _26463_, _26462_);
  and (_26464_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_26465_, _26417_, _26242_);
  or (_11342_, _26465_, _26464_);
  and (_26466_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_26467_, _26417_, _26185_);
  or (_11359_, _26467_, _26466_);
  nor (_26468_, _23153_, _23122_);
  and (_26469_, _23202_, _23183_);
  and (_26470_, _25618_, _23226_);
  and (_26471_, _26470_, _26469_);
  and (_26472_, _26471_, _26468_);
  and (_26473_, _25535_, _23215_);
  not (_26474_, _26473_);
  nor (_26475_, _26474_, _23729_);
  not (_26476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_26477_, _25904_, _26476_);
  or (_26478_, _26477_, _26475_);
  and (_26479_, _26478_, _26472_);
  nand (_26480_, _26472_, _23215_);
  and (_26481_, _26480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_26482_, _25536_, _25129_);
  nor (_26483_, _23201_, _23122_);
  and (_26484_, _26483_, _23777_);
  and (_26485_, _26484_, _26482_);
  or (_26486_, _26485_, _26481_);
  or (_26487_, _26486_, _26479_);
  nand (_26488_, _26485_, _25160_);
  and (_26489_, _26488_, _23049_);
  and (_11487_, _26489_, _26487_);
  and (_26491_, _25223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_26492_, _26491_, _25896_);
  and (_26493_, _26492_, _26472_);
  not (_26494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_26495_, _26472_, _25905_);
  nor (_26496_, _26495_, _26494_);
  or (_26497_, _26496_, _26485_);
  or (_26498_, _26497_, _26493_);
  not (_26499_, _26485_);
  or (_26500_, _26499_, _25258_);
  and (_26501_, _26500_, _23049_);
  and (_11532_, _26501_, _26498_);
  and (_26502_, _26472_, _25224_);
  or (_26503_, _26502_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_26504_, _26503_, _26499_);
  nand (_26505_, _26502_, _23729_);
  and (_26506_, _26505_, _26504_);
  nor (_26507_, _26499_, _25279_);
  or (_26508_, _26507_, _26506_);
  and (_11560_, _26508_, _23049_);
  and (_26510_, _26472_, _25131_);
  or (_26511_, _26510_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_26512_, _26511_, _26499_);
  nand (_26513_, _26510_, _23729_);
  and (_26514_, _26513_, _26512_);
  and (_26515_, _26485_, _25283_);
  or (_26516_, _26515_, _26514_);
  and (_11591_, _26516_, _23049_);
  and (_26517_, _26458_, _23830_);
  and (_26518_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_11683_, _26518_, _26517_);
  and (_26519_, _26458_, _25886_);
  and (_26520_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_11754_, _26520_, _26519_);
  and (_26521_, _26458_, _26170_);
  and (_26522_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_11774_, _26522_, _26521_);
  nor (_26523_, _23215_, _23137_);
  and (_26524_, _26523_, _23167_);
  and (_26525_, _26524_, _26472_);
  nand (_26526_, _26525_, _23729_);
  or (_26527_, _26525_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_26528_, _26527_, _26499_);
  and (_26529_, _26528_, _26526_);
  nor (_26530_, _26499_, _25332_);
  or (_26531_, _26530_, _26529_);
  and (_11795_, _26531_, _23049_);
  and (_26532_, _26472_, _26136_);
  nand (_26533_, _26532_, _23729_);
  or (_26534_, _26532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_26535_, _26534_, _26499_);
  and (_26536_, _26535_, _26533_);
  nor (_26537_, _26499_, _25362_);
  or (_26538_, _26537_, _26536_);
  and (_11846_, _26538_, _23049_);
  and (_26539_, _26242_, _26176_);
  and (_26540_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_11927_, _26540_, _26539_);
  and (_26541_, _26260_, _23775_);
  not (_26542_, _26541_);
  and (_26543_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  and (_26544_, _26541_, _25927_);
  or (_11958_, _26544_, _26543_);
  and (_26545_, _25611_, _23777_);
  and (_26546_, _26545_, _25902_);
  not (_26547_, _26546_);
  and (_26548_, _26471_, _25889_);
  and (_26549_, _26548_, _25224_);
  or (_26550_, _26549_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_26551_, _26550_, _26547_);
  nand (_26552_, _26549_, _23729_);
  and (_26553_, _26552_, _26551_);
  nor (_26554_, _26547_, _25279_);
  or (_26555_, _26554_, _26553_);
  and (_11999_, _26555_, _23049_);
  not (_26556_, _26130_);
  nor (_26557_, _26556_, _23729_);
  nor (_26558_, _25130_, _25534_);
  and (_26559_, _26558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_26560_, _26559_, _26557_);
  and (_26561_, _26560_, _26548_);
  not (_26562_, _26548_);
  nor (_26563_, _25130_, _23215_);
  or (_26564_, _26563_, _25131_);
  or (_26565_, _26564_, _26562_);
  and (_26566_, _26565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_26567_, _26566_, _26546_);
  or (_26568_, _26567_, _26561_);
  nand (_26569_, _26546_, _23824_);
  and (_26570_, _26569_, _23049_);
  and (_12030_, _26570_, _26568_);
  and (_26571_, _26548_, _26475_);
  nand (_26572_, _26548_, _23215_);
  and (_26573_, _26548_, _25905_);
  or (_26574_, _26573_, _26572_);
  and (_26575_, _26574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_26576_, _26575_, _26546_);
  or (_26577_, _26576_, _26571_);
  nand (_26578_, _26546_, _25160_);
  and (_26579_, _26578_, _23049_);
  and (_12084_, _26579_, _26577_);
  and (_26580_, _25223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_26581_, _26580_, _25896_);
  and (_26582_, _26581_, _26548_);
  not (_26583_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor (_26584_, _26573_, _26583_);
  or (_26585_, _26584_, _26546_);
  or (_26586_, _26585_, _26582_);
  or (_26587_, _26547_, _25258_);
  and (_26588_, _26587_, _23049_);
  and (_12107_, _26588_, _26586_);
  and (_26589_, _26548_, _25131_);
  or (_26590_, _26589_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_26591_, _26590_, _26547_);
  nand (_26592_, _26589_, _23729_);
  and (_26593_, _26592_, _26591_);
  and (_26594_, _26546_, _25283_);
  or (_26595_, _26594_, _26593_);
  and (_12128_, _26595_, _23049_);
  and (_26596_, _26355_, _26283_);
  and (_26597_, _26596_, _23768_);
  not (_26598_, _26596_);
  and (_26599_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_12189_, _26599_, _26597_);
  and (_26600_, _26596_, _26170_);
  and (_26601_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_12252_, _26601_, _26600_);
  and (_26602_, _26340_, _26204_);
  not (_26603_, _26602_);
  and (_26604_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_26605_, _26602_, _26242_);
  or (_12305_, _26605_, _26604_);
  and (_26606_, _26596_, _25927_);
  and (_26607_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_12346_, _26607_, _26606_);
  and (_26608_, _26548_, _26524_);
  nand (_26609_, _26608_, _23729_);
  or (_26610_, _26608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_26611_, _26610_, _26547_);
  and (_26612_, _26611_, _26609_);
  nor (_26613_, _26547_, _25332_);
  or (_26614_, _26613_, _26612_);
  and (_12397_, _26614_, _23049_);
  and (_26615_, _23848_, _23220_);
  and (_26616_, _26615_, _23768_);
  not (_26617_, _26615_);
  and (_26618_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_12508_, _26618_, _26616_);
  and (_26619_, _23201_, _23183_);
  and (_26620_, _25618_, _26619_);
  and (_26621_, _26620_, _25890_);
  and (_26622_, _26621_, _26130_);
  nand (_26623_, _26622_, _23729_);
  and (_26624_, _25902_, _25226_);
  not (_26625_, _26624_);
  or (_26626_, _26622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_26627_, _26626_, _26625_);
  and (_26628_, _26627_, _26623_);
  nor (_26629_, _26625_, _23824_);
  or (_26630_, _26629_, _26628_);
  and (_12608_, _26630_, _23049_);
  and (_26631_, _26621_, _25894_);
  or (_26632_, _26631_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_26633_, _26632_, _26625_);
  nand (_26634_, _26631_, _23729_);
  and (_26635_, _26634_, _26633_);
  and (_26636_, _26624_, _25258_);
  or (_26637_, _26636_, _26635_);
  and (_12623_, _26637_, _23049_);
  and (_26638_, _26621_, _25131_);
  or (_26639_, _26638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_26640_, _26639_, _26625_);
  nand (_26641_, _26638_, _23729_);
  and (_26642_, _26641_, _26640_);
  and (_26643_, _26624_, _25283_);
  or (_26644_, _26643_, _26642_);
  and (_12637_, _26644_, _23049_);
  and (_26645_, _26596_, _23830_);
  and (_26646_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_12750_, _26646_, _26645_);
  and (_26647_, _26596_, _26185_);
  and (_26648_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_27291_, _26648_, _26647_);
  and (_26649_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_26650_, _26417_, _26170_);
  or (_12791_, _26650_, _26649_);
  and (_26651_, _26596_, _26085_);
  and (_26652_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_12812_, _26652_, _26651_);
  and (_26653_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_26654_, _26417_, _25927_);
  or (_12923_, _26654_, _26653_);
  and (_26655_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  and (_26656_, _26214_, _26185_);
  or (_12944_, _26656_, _26655_);
  and (_26657_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_26658_, _26657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_26659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_26660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_26661_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _26660_);
  and (_26662_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_26663_, _26662_, _26661_);
  and (_26664_, _26663_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_26665_, _26664_, _26659_);
  not (_26666_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_26667_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_26668_, _26667_, _26666_);
  nand (_26669_, _26668_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_26670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_26671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_26672_, _26671_, _26670_);
  and (_26673_, _26672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_26674_, _26673_);
  and (_26675_, _26674_, _26669_);
  and (_26676_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_26677_, _26676_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_26678_, _26677_);
  and (_26679_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_26680_, _26679_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_26681_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_26682_, _26681_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_26683_, _26682_, _26680_);
  and (_26684_, _26683_, _26678_);
  and (_26685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_26686_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_26687_, _26686_);
  and (_26688_, _26687_, _26684_);
  and (_26689_, _26688_, _26675_);
  nor (_26690_, _26689_, _26665_);
  and (_26691_, _26690_, _26658_);
  not (_26692_, _26658_);
  and (_26693_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _26659_);
  not (_26694_, _26693_);
  not (_26695_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_26696_, _26668_, _26695_);
  not (_26697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_26698_, _26672_, _26697_);
  nor (_26699_, _26698_, _26696_);
  and (_26700_, _26685_, _26476_);
  not (_26701_, _26700_);
  and (_26702_, _26701_, _26699_);
  nor (_26703_, _26702_, _26694_);
  not (_26704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_26705_, _26676_, _26704_);
  not (_26706_, _26705_);
  not (_26707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_26708_, _26679_, _26707_);
  and (_26709_, _26681_, _26494_);
  nor (_26710_, _26709_, _26708_);
  and (_26711_, _26710_, _26706_);
  nor (_26712_, _26711_, _26694_);
  nor (_26713_, _26712_, _26703_);
  or (_26714_, _26713_, _26692_);
  and (_26715_, _26714_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_26716_, _26715_, _26691_);
  and (_13095_, _26716_, _23049_);
  and (_26717_, _26356_, _26242_);
  and (_26718_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_27290_, _26718_, _26717_);
  and (_26719_, _26356_, _26185_);
  and (_26720_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_13216_, _26720_, _26719_);
  and (_26721_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_26722_, _26602_, _25886_);
  or (_13327_, _26722_, _26721_);
  nor (_26723_, _26657_, _26660_);
  and (_26724_, _26723_, _26690_);
  not (_26725_, _26723_);
  or (_26726_, _26725_, _26713_);
  and (_26727_, _26726_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_26728_, _26727_, _26724_);
  and (_13348_, _26728_, _23049_);
  and (_26729_, _26170_, _26073_);
  and (_26730_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_13379_, _26730_, _26729_);
  not (_26731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_26732_, _26690_);
  and (_26733_, _26713_, _26732_);
  nor (_26734_, _26733_, _26657_);
  nor (_26735_, _26734_, _26731_);
  not (_26736_, _26657_);
  and (_26737_, _26673_, _26660_);
  or (_26738_, _26737_, _26731_);
  nor (_26739_, _26669_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_26740_, _26739_, _26686_);
  nand (_26741_, _26740_, _26738_);
  and (_26742_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_26743_, _26742_);
  nand (_26744_, _26743_, _26686_);
  and (_26745_, _26744_, _26741_);
  or (_26746_, _26745_, _26682_);
  not (_26747_, _26680_);
  not (_26748_, _26682_);
  or (_26749_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _26660_);
  or (_26750_, _26749_, _26748_);
  and (_26751_, _26750_, _26747_);
  and (_26752_, _26751_, _26746_);
  and (_26753_, _26742_, _26680_);
  or (_26754_, _26753_, _26677_);
  or (_26755_, _26754_, _26752_);
  or (_26756_, _26749_, _26678_);
  and (_26757_, _26756_, _26690_);
  and (_26758_, _26757_, _26755_);
  and (_26759_, _26698_, _26660_);
  or (_26760_, _26759_, _26731_);
  and (_26761_, _26696_, _26660_);
  nor (_26762_, _26761_, _26700_);
  nand (_26763_, _26762_, _26760_);
  nand (_26764_, _26743_, _26700_);
  and (_26765_, _26764_, _26763_);
  or (_26766_, _26765_, _26709_);
  not (_26767_, _26708_);
  not (_26768_, _26709_);
  or (_26769_, _26749_, _26768_);
  and (_26770_, _26769_, _26767_);
  and (_26771_, _26770_, _26766_);
  and (_26772_, _26742_, _26708_);
  or (_26773_, _26772_, _26705_);
  or (_26774_, _26773_, _26771_);
  nor (_26775_, _26713_, _26690_);
  and (_26776_, _26775_, _26706_);
  and (_26777_, _26749_, _26775_);
  or (_26778_, _26777_, _26776_);
  and (_26779_, _26778_, _26774_);
  or (_26780_, _26779_, _26758_);
  and (_26781_, _26780_, _26736_);
  or (_26782_, _26781_, _26735_);
  and (_13488_, _26782_, _23049_);
  and (_26783_, _26355_, _23775_);
  and (_26784_, _26783_, _23830_);
  not (_26785_, _26783_);
  and (_26786_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_27284_, _26786_, _26784_);
  nand (_26787_, _26733_, _26658_);
  nor (_26788_, _26690_, _26657_);
  or (_26789_, _26788_, _26660_);
  and (_26790_, _26789_, _23049_);
  and (_13569_, _26790_, _26787_);
  and (_26791_, _26783_, _25886_);
  and (_26792_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_27283_, _26792_, _26791_);
  and (_26793_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_26794_, _26602_, _26170_);
  or (_13620_, _26794_, _26793_);
  not (_26795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_26796_, _26734_, _26795_);
  and (_26797_, _26673_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_26798_, _26797_, _26795_);
  nor (_26799_, _26669_, _26660_);
  nor (_26800_, _26799_, _26686_);
  nand (_26801_, _26800_, _26798_);
  and (_26802_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _26660_);
  or (_26803_, _26802_, _26687_);
  and (_26804_, _26803_, _26801_);
  or (_26805_, _26804_, _26682_);
  or (_26806_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_26807_, _26806_, _26748_);
  and (_26808_, _26807_, _26747_);
  and (_26809_, _26808_, _26805_);
  and (_26810_, _26802_, _26680_);
  or (_26811_, _26810_, _26677_);
  or (_26812_, _26811_, _26809_);
  or (_26813_, _26806_, _26678_);
  and (_26814_, _26813_, _26690_);
  and (_26815_, _26814_, _26812_);
  and (_26816_, _26698_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_26817_, _26816_, _26795_);
  and (_26818_, _26696_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_26819_, _26818_, _26700_);
  nand (_26820_, _26819_, _26817_);
  or (_26821_, _26802_, _26701_);
  and (_26822_, _26821_, _26820_);
  or (_26823_, _26822_, _26709_);
  or (_26824_, _26806_, _26768_);
  and (_26825_, _26824_, _26767_);
  and (_26826_, _26825_, _26823_);
  and (_26827_, _26802_, _26708_);
  or (_26828_, _26827_, _26705_);
  or (_26829_, _26828_, _26826_);
  and (_26830_, _26806_, _26775_);
  or (_26831_, _26830_, _26776_);
  and (_26832_, _26831_, _26829_);
  or (_26833_, _26832_, _26815_);
  and (_26834_, _26833_, _26736_);
  or (_26835_, _26834_, _26796_);
  and (_13761_, _26835_, _23049_);
  and (_26836_, _26783_, _26242_);
  and (_26837_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_14032_, _26837_, _26836_);
  and (_26838_, _26783_, _26185_);
  and (_26839_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_14073_, _26839_, _26838_);
  and (_26840_, _26657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_26841_, _26840_, _26734_);
  and (_14164_, _26841_, _23049_);
  nor (_26842_, _26708_, _26705_);
  nor (_26843_, _26709_, _26700_);
  and (_26844_, _26843_, _26842_);
  nand (_26845_, _26844_, _26693_);
  or (_26846_, _26845_, _26699_);
  nor (_26847_, _26846_, _26690_);
  and (_26848_, _26657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_26849_, _26665_, _26657_);
  not (_26850_, _26675_);
  and (_26851_, _26688_, _26850_);
  and (_26852_, _26851_, _26849_);
  or (_26853_, _26852_, _26848_);
  or (_26854_, _26853_, _26847_);
  and (_14185_, _26854_, _23049_);
  nand (_26855_, _26699_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand (_26856_, _26855_, _26843_);
  and (_26857_, _26856_, _26842_);
  and (_26858_, _26857_, _26775_);
  nor (_26859_, _26680_, _26677_);
  or (_26860_, _26686_, _26682_);
  and (_26861_, _26675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_26862_, _26861_, _26860_);
  and (_26863_, _26862_, _26859_);
  and (_26864_, _26863_, _26690_);
  or (_26865_, _26864_, _26858_);
  or (_26866_, _26865_, _26657_);
  or (_26867_, _26736_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26868_, _26867_, _23049_);
  and (_14206_, _26868_, _26866_);
  nor (_26869_, _26698_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_26870_, _26869_, _26696_);
  or (_26871_, _26870_, _26700_);
  and (_26872_, _26871_, _26768_);
  or (_26873_, _26872_, _26708_);
  and (_00001_, _26873_, _26776_);
  or (_00002_, _26673_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_00003_, _00002_, _26669_);
  or (_00004_, _00003_, _26686_);
  and (_00005_, _00004_, _26748_);
  or (_00006_, _00005_, _26680_);
  and (_00007_, _26690_, _26678_);
  and (_00008_, _00007_, _00006_);
  or (_00009_, _00008_, _26657_);
  or (_00010_, _00009_, _00001_);
  nand (_00011_, _26657_, _23832_);
  and (_00012_, _00011_, _23049_);
  and (_14243_, _00012_, _00010_);
  and (_00013_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_00014_, _26602_, _26085_);
  or (_27055_, _00014_, _00013_);
  and (_00015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _23049_);
  and (_14273_, _00015_, _26657_);
  and (_00016_, _26355_, _26213_);
  and (_00017_, _00016_, _26185_);
  not (_00018_, _00016_);
  and (_00019_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_27280_, _00019_, _00017_);
  and (_00020_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_00021_, _26413_, _25927_);
  or (_27068_, _00021_, _00020_);
  and (_00022_, _26283_, _26204_);
  not (_00023_, _00022_);
  and (_00024_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and (_00025_, _00022_, _25886_);
  or (_14576_, _00025_, _00024_);
  and (_00026_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_00027_, _00022_, _26170_);
  or (_14602_, _00027_, _00026_);
  and (_00028_, _26783_, _25927_);
  and (_00029_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_14716_, _00029_, _00028_);
  and (_00030_, _26783_, _23768_);
  and (_00031_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_14751_, _00031_, _00030_);
  and (_00032_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and (_00033_, _00022_, _26242_);
  or (_15030_, _00033_, _00032_);
  and (_00034_, _26615_, _26170_);
  and (_00035_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_15068_, _00035_, _00034_);
  and (_00036_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_00037_, _00022_, _26185_);
  or (_15082_, _00037_, _00036_);
  and (_00038_, _26374_, _26355_);
  and (_00039_, _00038_, _25886_);
  not (_00041_, _00038_);
  and (_00042_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_27286_, _00042_, _00039_);
  and (_00043_, _26329_, _23830_);
  and (_00044_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_15151_, _00044_, _00043_);
  and (_00045_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_00046_, _00022_, _26085_);
  or (_15165_, _00046_, _00045_);
  and (_00047_, _00038_, _26170_);
  and (_00048_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_15180_, _00048_, _00047_);
  and (_00049_, _25938_, _25914_);
  and (_00050_, _00049_, _25927_);
  not (_00051_, _00049_);
  and (_00052_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_15240_, _00052_, _00050_);
  and (_00053_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_00055_, _25927_, _23780_);
  or (_15256_, _00055_, _00053_);
  and (_00056_, _00038_, _26185_);
  and (_00057_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_15616_, _00057_, _00056_);
  and (_00059_, _26204_, _23847_);
  not (_00060_, _00059_);
  and (_00061_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_00063_, _00059_, _26185_);
  or (_15637_, _00063_, _00061_);
  and (_00064_, _00038_, _26085_);
  and (_00065_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_15758_, _00065_, _00064_);
  and (_00066_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_00067_, _00059_, _26085_);
  or (_15839_, _00067_, _00066_);
  and (_00068_, _25901_, _25894_);
  and (_00069_, _00068_, _25226_);
  not (_00070_, _00069_);
  and (_00071_, _26131_, _25226_);
  and (_00072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_00073_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_00074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00076_, _00074_, _23049_);
  and (_00077_, _00076_, _00073_);
  not (_00078_, _00072_);
  and (_00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00080_, _00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00081_, _00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00082_, _00081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00083_, _00082_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00084_, _00083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00085_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_00086_, _00085_, _00078_);
  nand (_00087_, _00086_, _00077_);
  nor (_00088_, _00087_, _00071_);
  and (_15990_, _00088_, _00070_);
  and (_00089_, _26283_, _26260_);
  not (_00090_, _00089_);
  and (_00091_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  and (_00092_, _00089_, _23768_);
  or (_27166_, _00092_, _00091_);
  and (_00093_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_00094_, _00059_, _26242_);
  or (_16454_, _00094_, _00093_);
  and (_00095_, _26191_, _23229_);
  and (_00096_, _00095_, _26150_);
  and (_00097_, _00096_, _26242_);
  not (_00099_, _00096_);
  and (_00100_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_27325_, _00100_, _00097_);
  and (_00101_, _00096_, _26185_);
  and (_00102_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_16605_, _00102_, _00101_);
  and (_00103_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_00104_, _00022_, _23768_);
  or (_16646_, _00104_, _00103_);
  and (_00105_, _26258_, _23230_);
  and (_00106_, _00105_, _25927_);
  not (_00107_, _00105_);
  and (_00108_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_16927_, _00108_, _00106_);
  and (_00109_, _00105_, _25886_);
  and (_00110_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_16948_, _00110_, _00109_);
  and (_00111_, _00105_, _23830_);
  and (_00112_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_17068_, _00112_, _00111_);
  and (_00113_, _00105_, _26185_);
  and (_00114_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_17089_, _00114_, _00113_);
  and (_00115_, _26190_, _23230_);
  and (_00116_, _00115_, _26242_);
  not (_00117_, _00115_);
  and (_00118_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_17400_, _00118_, _00116_);
  and (_00119_, _26213_, _23230_);
  and (_00120_, _00119_, _23768_);
  not (_00121_, _00119_);
  and (_00122_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_17431_, _00122_, _00120_);
  and (_00123_, _00119_, _26170_);
  and (_00124_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_17452_, _00124_, _00123_);
  and (_00125_, _00119_, _23830_);
  and (_00126_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_27090_, _00126_, _00125_);
  and (_00127_, _26308_, _26242_);
  and (_00128_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_27271_, _00128_, _00127_);
  and (_00129_, _26301_, _23768_);
  and (_00130_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_27242_, _00130_, _00129_);
  and (_00131_, _00119_, _26185_);
  and (_00132_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_27091_, _00132_, _00131_);
  and (_00133_, _23775_, _23230_);
  and (_00134_, _00133_, _25927_);
  not (_00135_, _00133_);
  and (_00136_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_18851_, _00136_, _00134_);
  not (_00137_, _22738_);
  or (_00138_, _22909_, _00137_);
  or (_00139_, _22738_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_00140_, _00139_, _23049_);
  and (_26896_[7], _00140_, _00138_);
  and (_00141_, _26258_, _26204_);
  not (_00142_, _00141_);
  and (_00143_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_00144_, _00141_, _26242_);
  or (_27052_, _00144_, _00143_);
  and (_00145_, _00133_, _26170_);
  and (_00146_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_19316_, _00146_, _00145_);
  and (_00147_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_00148_, _26422_, _26085_);
  or (_27083_, _00148_, _00147_);
  and (_00149_, _00133_, _26085_);
  and (_00150_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_19380_, _00150_, _00149_);
  and (_00151_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_00152_, _00059_, _23768_);
  or (_19450_, _00152_, _00151_);
  and (_00153_, _00133_, _26185_);
  and (_00154_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_19708_, _00154_, _00153_);
  and (_00155_, _26374_, _23230_);
  and (_00156_, _00155_, _23768_);
  not (_00157_, _00155_);
  and (_00158_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_19729_, _00158_, _00156_);
  and (_00159_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_00160_, _26413_, _23768_);
  or (_19784_, _00160_, _00159_);
  and (_00161_, _00155_, _25927_);
  and (_00162_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_19825_, _00162_, _00161_);
  and (_00163_, _00155_, _23830_);
  and (_00164_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_21660_, _00164_, _00163_);
  and (_00165_, _00155_, _26085_);
  and (_00166_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_21981_, _00166_, _00165_);
  and (_00167_, _00155_, _26242_);
  and (_00168_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_27132_, _00168_, _00167_);
  and (_00169_, _00105_, _23768_);
  and (_00170_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_27151_, _00170_, _00169_);
  and (_00171_, _23847_, _23230_);
  and (_00172_, _00171_, _23768_);
  not (_00173_, _00171_);
  and (_00174_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_22253_, _00174_, _00172_);
  and (_00175_, _00171_, _25927_);
  and (_00176_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_22592_, _00176_, _00175_);
  and (_00177_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  and (_00178_, _26541_, _23768_);
  or (_22593_, _00178_, _00177_);
  and (_00179_, _00171_, _25886_);
  and (_00180_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_22594_, _00180_, _00179_);
  and (_00181_, _00171_, _26085_);
  and (_00182_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_22595_, _00182_, _00181_);
  and (_00183_, _00171_, _26242_);
  and (_00184_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_22596_, _00184_, _00183_);
  and (_00185_, _26283_, _23230_);
  and (_00186_, _00185_, _23768_);
  not (_00187_, _00185_);
  and (_00188_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_27182_, _00188_, _00186_);
  and (_00189_, _26473_, _25901_);
  and (_00190_, _00189_, _25226_);
  nand (_00191_, _00190_, _25332_);
  not (_00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00193_, _00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00194_);
  nor (_00196_, _00195_, _00193_);
  not (_00197_, _00196_);
  not (_00199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_00200_, t1_i);
  and (_00201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00200_);
  nor (_00202_, _00201_, _00199_);
  not (_00203_, _00202_);
  not (_00204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00205_, _00204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_00206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_00207_, _00206_);
  and (_00208_, _00207_, _00205_);
  and (_00209_, _00208_, _00203_);
  and (_00210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00212_, _00211_, _00210_);
  and (_00213_, _00212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00214_, _00213_, _00209_);
  and (_00215_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00216_, _00215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00217_, _00215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00218_, _00217_, _00216_);
  and (_00219_, _00218_, _00197_);
  and (_00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00221_, _00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00222_, _00221_, _00214_);
  and (_00223_, _00222_, _00193_);
  and (_00224_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00225_, _00224_, _00219_);
  and (_00226_, _26137_, _25226_);
  nor (_00227_, _00226_, _00225_);
  or (_00228_, _00226_, _00196_);
  and (_00229_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_00230_, _00229_, _00227_);
  or (_00231_, _00230_, _00190_);
  and (_00232_, _00231_, _23049_);
  and (_22598_, _00232_, _00191_);
  and (_00234_, _00185_, _26170_);
  and (_00235_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_27184_, _00235_, _00234_);
  and (_00236_, _00185_, _23830_);
  and (_00237_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_22599_, _00237_, _00236_);
  and (_00238_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  and (_00239_, _26214_, _26085_);
  or (_22600_, _00239_, _00238_);
  and (_00241_, _00185_, _26242_);
  and (_00242_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_22602_, _00242_, _00241_);
  not (_00243_, _26524_);
  nor (_00244_, _00243_, _23729_);
  and (_00246_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_00247_, _00246_, _00244_);
  and (_00249_, _26469_, _25627_);
  and (_00250_, _00249_, _00247_);
  not (_00251_, _00249_);
  and (_00252_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_00253_, _00252_, _00250_);
  and (_00254_, _00253_, _25618_);
  and (_00255_, _25131_, _23153_);
  and (_00256_, _26483_, _00255_);
  and (_00257_, _00256_, _23777_);
  nand (_00258_, _00257_, _25332_);
  or (_00259_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_00260_, _00259_, _25128_);
  and (_00261_, _00260_, _00258_);
  and (_00263_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_00264_, _00263_, rst);
  or (_00265_, _00264_, _00261_);
  or (_22603_, _00265_, _00254_);
  and (_00266_, _26224_, _23230_);
  and (_00267_, _00266_, _23768_);
  not (_00268_, _00266_);
  and (_00269_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_22604_, _00269_, _00267_);
  and (_00270_, _00249_, _26136_);
  or (_00271_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00272_, _00271_, _25618_);
  nand (_00273_, _00270_, _23729_);
  and (_00274_, _00273_, _00272_);
  nand (_00275_, _00257_, _25362_);
  or (_00276_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00277_, _00276_, _25128_);
  and (_00278_, _00277_, _00275_);
  and (_00279_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_00280_, _00279_, rst);
  or (_00281_, _00280_, _00278_);
  or (_22605_, _00281_, _00274_);
  and (_00282_, _00266_, _26170_);
  and (_00283_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_22606_, _00283_, _00282_);
  and (_00284_, _26615_, _23830_);
  and (_00285_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_22607_, _00285_, _00284_);
  and (_00286_, _00266_, _25886_);
  and (_00287_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_27203_, _00287_, _00286_);
  and (_00288_, _00266_, _26185_);
  and (_00289_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_22608_, _00289_, _00288_);
  and (_00290_, _00266_, _26242_);
  and (_00291_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_27204_, _00291_, _00290_);
  and (_00292_, _26150_, _23230_);
  and (_00293_, _00292_, _25927_);
  not (_00294_, _00292_);
  and (_00295_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_27216_, _00295_, _00293_);
  and (_00296_, _00292_, _26170_);
  and (_00297_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_22609_, _00297_, _00296_);
  and (_00298_, _00292_, _26185_);
  and (_00299_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_22610_, _00299_, _00298_);
  and (_00300_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_00301_, _00059_, _25886_);
  or (_22611_, _00301_, _00300_);
  and (_26917_[0], _22835_, _23049_);
  nor (_26917_[1], _22860_, rst);
  and (_26917_[2], _22782_, _23049_);
  nor (_26917_[3], _25162_, rst);
  or (_00302_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_00303_, _25858_, _22815_);
  and (_00304_, _00303_, _23049_);
  and (_26935_[0], _00304_, _00302_);
  or (_00305_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_00306_, _25858_, _22837_);
  and (_00307_, _00306_, _23049_);
  and (_26935_[1], _00307_, _00305_);
  or (_00308_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_00309_, _25858_, _22758_);
  and (_00310_, _00309_, _23049_);
  and (_26935_[2], _00310_, _00308_);
  or (_00311_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_00312_, _25858_, _22794_);
  and (_00313_, _00312_, _23049_);
  and (_26935_[3], _00313_, _00311_);
  and (_00314_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00315_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_00316_, _00315_, _00314_);
  and (_26935_[4], _00316_, _23049_);
  or (_00317_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_00318_, _25858_, _22875_);
  and (_00319_, _00318_, _23049_);
  and (_26935_[5], _00319_, _00317_);
  or (_00320_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_00321_, _25858_, _22914_);
  and (_00322_, _00321_, _23049_);
  and (_26935_[6], _00322_, _00320_);
  or (_00323_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_00324_, _25858_, _22901_);
  and (_00325_, _00324_, _23049_);
  and (_26935_[7], _00325_, _00323_);
  or (_00326_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_00327_, _25858_, _24465_);
  and (_00328_, _00327_, _23049_);
  and (_26935_[8], _00328_, _00326_);
  or (_00329_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_00330_, _25858_, _24425_);
  and (_00331_, _00330_, _23049_);
  and (_26935_[9], _00331_, _00329_);
  or (_00332_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_00333_, _25858_, _24390_);
  and (_00334_, _00333_, _23049_);
  and (_26935_[10], _00334_, _00332_);
  or (_00335_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_00336_, _25858_, _24346_);
  and (_00337_, _00336_, _23049_);
  and (_26935_[11], _00337_, _00335_);
  and (_00338_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00339_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or (_00340_, _00339_, _00338_);
  and (_26935_[12], _00340_, _23049_);
  or (_00341_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_00342_, _25858_, _24278_);
  and (_00344_, _00342_, _23049_);
  and (_26935_[13], _00344_, _00341_);
  or (_00345_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_00347_, _25858_, _24235_);
  and (_00348_, _00347_, _23049_);
  and (_26935_[14], _00348_, _00345_);
  or (_00349_, _25858_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_00350_, _25858_, _24188_);
  and (_00351_, _00350_, _23049_);
  and (_26935_[15], _00351_, _00349_);
  and (_00352_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00353_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_00354_, _00353_, _00352_);
  and (_26935_[16], _00354_, _23049_);
  and (_00355_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00356_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_00357_, _00356_, _00355_);
  and (_26935_[17], _00357_, _23049_);
  and (_00358_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00359_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or (_00360_, _00359_, _00358_);
  and (_26935_[18], _00360_, _23049_);
  and (_00361_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00362_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or (_00363_, _00362_, _00361_);
  and (_26935_[19], _00363_, _23049_);
  and (_00364_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00365_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_00366_, _00365_, _00364_);
  and (_26935_[20], _00366_, _23049_);
  and (_00367_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00368_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_00369_, _00368_, _00367_);
  and (_26935_[21], _00369_, _23049_);
  and (_00370_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00371_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_00372_, _00371_, _00370_);
  and (_26935_[22], _00372_, _23049_);
  and (_00373_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00374_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_00375_, _00374_, _00373_);
  and (_26935_[23], _00375_, _23049_);
  and (_00376_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00377_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_00378_, _00377_, _00376_);
  and (_26935_[24], _00378_, _23049_);
  and (_00379_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00380_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_00381_, _00380_, _00379_);
  and (_26935_[25], _00381_, _23049_);
  and (_00382_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00383_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_00384_, _00383_, _00382_);
  and (_26935_[26], _00384_, _23049_);
  and (_00385_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00387_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_00388_, _00387_, _00385_);
  and (_26935_[27], _00388_, _23049_);
  and (_00389_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00390_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or (_00391_, _00390_, _00389_);
  and (_26935_[28], _00391_, _23049_);
  and (_00392_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00393_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_00394_, _00393_, _00392_);
  and (_26935_[29], _00394_, _23049_);
  and (_00395_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00396_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or (_00397_, _00396_, _00395_);
  and (_26935_[30], _00397_, _23049_);
  and (_00398_, _00292_, _26242_);
  and (_00399_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_27217_, _00399_, _00398_);
  and (_00400_, _26421_, _23230_);
  and (_00401_, _00400_, _25927_);
  not (_00402_, _00400_);
  and (_00403_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_27218_, _00403_, _00401_);
  and (_26918_[0], _25655_, _23049_);
  and (_26918_[1], _25742_, _23049_);
  and (_26918_[2], _25693_, _23049_);
  and (_26918_[3], _25212_, _23049_);
  and (_26918_[4], _25475_, _23049_);
  and (_26918_[5], _25518_, _23049_);
  and (_26918_[6], _25394_, _23049_);
  nand (_00404_, _26469_, _25616_);
  nor (_00405_, _00404_, _00243_);
  nand (_00406_, _00405_, _23729_);
  or (_00407_, _00405_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_00408_, _00407_, _25618_);
  and (_00409_, _00408_, _00406_);
  and (_00410_, _26545_, _00255_);
  nand (_00411_, _00410_, _25332_);
  or (_00412_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_00413_, _00412_, _25128_);
  and (_00414_, _00413_, _00411_);
  and (_00415_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_00416_, _00415_, rst);
  or (_00417_, _00416_, _00414_);
  or (_22612_, _00417_, _00409_);
  and (_00418_, _26190_, _23779_);
  not (_00419_, _00418_);
  and (_00420_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  and (_00421_, _00418_, _23768_);
  or (_27063_, _00421_, _00420_);
  and (_00422_, _00400_, _26170_);
  and (_00423_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_27219_, _00423_, _00422_);
  and (_00424_, _00400_, _26085_);
  and (_00425_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_22613_, _00425_, _00424_);
  and (_00426_, _00400_, _26185_);
  and (_00427_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_22614_, _00427_, _00426_);
  and (_00428_, _26340_, _23230_);
  and (_00429_, _00428_, _23768_);
  not (_00430_, _00428_);
  and (_00431_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_22615_, _00431_, _00429_);
  and (_26892_[7], _22909_, _23049_);
  or (_00432_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_00433_, _00432_, _25618_);
  and (_00434_, _00249_, _25131_);
  nand (_00435_, _00434_, _23729_);
  and (_00436_, _00435_, _00433_);
  nand (_00437_, _00257_, _23761_);
  and (_00438_, _00432_, _25128_);
  and (_00439_, _00438_, _00437_);
  not (_00440_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_00441_, _25127_, _00440_);
  or (_00442_, _00441_, rst);
  or (_00443_, _00442_, _00439_);
  or (_22616_, _00443_, _00436_);
  and (_00444_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_00445_, _00059_, _26170_);
  or (_22617_, _00445_, _00444_);
  and (_00446_, _00428_, _25927_);
  and (_00447_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_22618_, _00447_, _00446_);
  nor (_00448_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_00449_, _00448_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_26939_, _00449_, _23049_);
  and (_26932_, _23049_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00450_, _26932_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_26938_, _00450_, _26939_);
  nand (_00451_, _22735_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_26937_, _00451_, _23049_);
  or (_00452_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_00453_, _25858_, _22895_);
  and (_00454_, _00453_, _23049_);
  and (_26936_[31], _00454_, _00452_);
  and (_00455_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_00456_, _25859_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_00457_, _00456_, _00455_);
  and (_26935_[31], _00457_, _23049_);
  and (_00458_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_00459_, _00458_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  or (_00460_, _00459_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_26934_[3], _00460_, _23049_);
  not (_00461_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_00462_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00463_, _00462_, _00461_);
  and (_00464_, _00462_, _00461_);
  nor (_00465_, _00464_, _00463_);
  not (_00466_, _00465_);
  and (_00467_, _00466_, _26934_[3]);
  nor (_00468_, _00463_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00469_, _00463_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_00470_, _00469_, _00468_);
  nor (_00471_, _00458_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00472_, _00471_, _00459_);
  or (_00473_, _00472_, _00462_);
  and (_00474_, _00473_, _00470_);
  and (_26933_, _00474_, _00467_);
  not (_00475_, _24756_);
  and (_00476_, _24784_, _24645_);
  nor (_00477_, _00476_, _00475_);
  and (_00478_, _00476_, _00475_);
  or (_00479_, _00478_, _00477_);
  and (_00480_, _00479_, _23752_);
  nand (_00481_, _24979_, _24976_);
  or (_00482_, _24979_, _24976_);
  and (_00483_, _00482_, _00481_);
  and (_00484_, _00483_, _24794_);
  or (_00485_, _23601_, _23238_);
  and (_00486_, _00485_, _25556_);
  and (_00487_, _23715_, _23710_);
  and (_00488_, _23807_, _23448_);
  or (_00489_, _00488_, _23757_);
  nor (_00490_, _23679_, _23476_);
  and (_00492_, _23689_, _23714_);
  or (_00493_, _00492_, _00490_);
  nor (_00494_, _00493_, _00489_);
  and (_00495_, _00494_, _23746_);
  nand (_00496_, _00495_, _23741_);
  or (_00497_, _00496_, _00487_);
  or (_00498_, _00497_, _00486_);
  or (_00499_, _00498_, _00484_);
  or (_00500_, _00499_, _00480_);
  and (_00501_, _24180_, _24174_);
  and (_00502_, _00501_, _24170_);
  or (_00503_, _00502_, _24179_);
  and (_00504_, _00503_, _00500_);
  and (_00505_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00506_, _24482_, _24172_);
  and (_00507_, _24178_, _24174_);
  and (_00508_, _00507_, _24499_);
  or (_00509_, _00508_, _00506_);
  or (_00510_, _00509_, _00505_);
  nor (_00511_, _24502_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_00512_, _00511_, _24503_);
  and (_00513_, _00512_, _24183_);
  or (_00514_, _00513_, _00510_);
  or (_00515_, _00514_, _00504_);
  and (_00516_, _00515_, _25762_);
  not (_00517_, _25762_);
  and (_00518_, _00517_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_00519_, _00518_, _00516_);
  and (_26921_[0], _00519_, _23049_);
  nand (_00520_, _24783_, _24675_);
  or (_00521_, _24758_, _24753_);
  and (_00522_, _00521_, _24759_);
  or (_00523_, _00522_, _00520_);
  or (_00524_, _24784_, _24750_);
  and (_00525_, _00524_, _00523_);
  and (_00526_, _00525_, _23752_);
  nand (_00527_, _00481_, _24921_);
  nand (_00528_, _00527_, _24977_);
  or (_00529_, _00527_, _24977_);
  and (_00530_, _00529_, _00528_);
  and (_00531_, _00530_, _24794_);
  nor (_00532_, _23487_, _23485_);
  nor (_00533_, _00532_, _23488_);
  or (_00534_, _00533_, _23541_);
  not (_00535_, _23238_);
  nor (_00536_, _23542_, _00535_);
  and (_00537_, _00536_, _00534_);
  nor (_00538_, _23642_, _23640_);
  or (_00539_, _00538_, _23643_);
  and (_00540_, _00539_, _23601_);
  or (_00541_, _00540_, _00537_);
  nor (_00542_, _23666_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_00543_, _00542_, _23448_);
  nor (_00544_, _00542_, _23448_);
  or (_00545_, _00544_, _00543_);
  and (_00546_, _00545_, _23664_);
  nor (_00547_, _23748_, _23476_);
  and (_00548_, _23807_, _23412_);
  and (_00549_, _23711_, _23448_);
  or (_00550_, _00549_, _00548_);
  or (_00551_, _00550_, _00547_);
  or (_00552_, _00551_, _25277_);
  nor (_00553_, _00552_, _00546_);
  nand (_00554_, _00553_, _25268_);
  or (_00555_, _00554_, _00541_);
  or (_00556_, _00555_, _00531_);
  or (_00557_, _00556_, _00526_);
  and (_00558_, _00557_, _00503_);
  and (_00559_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00560_, _24441_, _24172_);
  and (_00561_, _00507_, _24457_);
  or (_00562_, _00561_, _00560_);
  or (_00563_, _00562_, _00559_);
  nor (_00564_, _24505_, _24503_);
  nor (_00565_, _00564_, _24506_);
  and (_00566_, _00565_, _24183_);
  or (_00567_, _00566_, _00563_);
  or (_00568_, _00567_, _00558_);
  and (_00569_, _00568_, _25762_);
  and (_00570_, _00517_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00571_, _00570_, _00569_);
  and (_26921_[1], _00571_, _23049_);
  nand (_00572_, _00528_, _24915_);
  and (_00573_, _00572_, _24924_);
  nor (_00574_, _00572_, _24924_);
  nor (_00575_, _00574_, _00573_);
  nand (_00576_, _00575_, _24794_);
  not (_00577_, _23752_);
  not (_00578_, _24771_);
  and (_00579_, _24770_, _24760_);
  nor (_00580_, _00579_, _00578_);
  nor (_00581_, _00580_, _00520_);
  nor (_00582_, _24784_, _24766_);
  or (_00583_, _00582_, _00581_);
  or (_00584_, _00583_, _00577_);
  nor (_00585_, _25559_, _23602_);
  and (_00586_, _23747_, _23448_);
  not (_00587_, _00586_);
  not (_00588_, _23807_);
  or (_00589_, _00588_, _23378_);
  and (_00590_, _23711_, _23412_);
  not (_00591_, _00590_);
  and (_00592_, _00591_, _00589_);
  and (_00593_, _00592_, _00587_);
  and (_00594_, _00593_, _25256_);
  not (_00595_, _00594_);
  nor (_00596_, _00595_, _00585_);
  nor (_00597_, _23544_, _23542_);
  nor (_00598_, _00597_, _00535_);
  and (_00599_, _00598_, _23546_);
  and (_00600_, _23665_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00601_, _00544_, _25252_);
  nor (_00602_, _00601_, _00600_);
  nor (_00603_, _00602_, _23679_);
  nor (_00604_, _00603_, _00599_);
  and (_00605_, _00604_, _00596_);
  and (_00606_, _00605_, _25244_);
  and (_00607_, _00606_, _00584_);
  and (_00608_, _00607_, _00576_);
  not (_00609_, _00608_);
  and (_00610_, _00609_, _00503_);
  nor (_00611_, _24510_, _24508_);
  nor (_00612_, _00611_, _24512_);
  and (_00613_, _00612_, _24183_);
  and (_00614_, _24402_, _24172_);
  and (_00615_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_00616_, _00507_, _24418_);
  or (_00617_, _00616_, _00615_);
  or (_00618_, _00617_, _00614_);
  or (_00619_, _00618_, _00613_);
  or (_00620_, _00619_, _00610_);
  and (_00621_, _00620_, _25762_);
  not (_00622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00623_, _25858_, _00622_);
  and (_00624_, _25858_, _00622_);
  nor (_00625_, _00624_, _00623_);
  and (_00626_, _00625_, _00517_);
  or (_00627_, _00626_, _00621_);
  and (_26921_[2], _00627_, _23049_);
  or (_00628_, _24772_, _24744_);
  and (_00629_, _24771_, _24767_);
  or (_00630_, _00629_, _00628_);
  nand (_00631_, _00629_, _00628_);
  and (_00632_, _00631_, _00630_);
  or (_00633_, _00632_, _00520_);
  or (_00634_, _24784_, _24743_);
  and (_00635_, _00634_, _00633_);
  and (_00636_, _00635_, _23752_);
  nor (_00637_, _24925_, _00573_);
  nor (_00638_, _00637_, _24983_);
  and (_00639_, _00638_, _24794_);
  nor (_00640_, _25554_, _23602_);
  nand (_00641_, _23546_, _23494_);
  nor (_00642_, _23547_, _00535_);
  and (_00643_, _00642_, _00641_);
  not (_00644_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00645_, _23665_, _00644_);
  or (_00646_, _00645_, _23795_);
  nor (_00647_, _23666_, _23679_);
  and (_00648_, _00647_, _00646_);
  and (_00649_, _23711_, _23795_);
  nor (_00650_, _00588_, _23348_);
  and (_00651_, _23747_, _23412_);
  or (_00652_, _00651_, _00650_);
  or (_00653_, _00652_, _00649_);
  or (_00654_, _00653_, _00648_);
  or (_00655_, _00654_, _25159_);
  or (_00656_, _00655_, _00643_);
  or (_00657_, _00656_, _00640_);
  or (_00658_, _00657_, _00639_);
  or (_00659_, _00658_, _00636_);
  and (_00660_, _00659_, _00503_);
  and (_00661_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not (_00662_, _24361_);
  and (_00663_, _00662_, _24172_);
  and (_00664_, _00507_, _25214_);
  or (_00665_, _00664_, _00663_);
  or (_00666_, _00665_, _00661_);
  or (_00667_, _00666_, _00660_);
  nor (_00668_, _24513_, _24383_);
  nor (_00669_, _00668_, _24514_);
  nand (_00670_, _00669_, _24183_);
  nand (_00671_, _00670_, _25762_);
  or (_00673_, _00671_, _00667_);
  and (_00674_, _00623_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00675_, _00623_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00676_, _00675_, _00674_);
  or (_00677_, _00676_, _25762_);
  and (_00678_, _00677_, _23049_);
  and (_26921_[3], _00678_, _00673_);
  and (_00679_, _24778_, _24776_);
  nor (_00680_, _24778_, _24776_);
  or (_00681_, _00680_, _00679_);
  nand (_00682_, _00681_, _24784_);
  or (_00683_, _24784_, _24731_);
  and (_00684_, _00683_, _00682_);
  nand (_00685_, _00684_, _23752_);
  nand (_00686_, _24984_, _24983_);
  or (_00687_, _24984_, _24983_);
  and (_00688_, _00687_, _00686_);
  nand (_00689_, _00688_, _24794_);
  nor (_00690_, _23550_, _23357_);
  not (_00691_, _00690_);
  nor (_00692_, _23551_, _00535_);
  and (_00693_, _00692_, _00691_);
  not (_00694_, _00693_);
  and (_00695_, _25544_, _23601_);
  nor (_00696_, _23667_, _23661_);
  and (_00697_, _23711_, _23661_);
  nor (_00698_, _23668_, _23679_);
  nor (_00699_, _00698_, _00697_);
  nor (_00700_, _00699_, _00696_);
  nor (_00701_, _23748_, _23378_);
  not (_00702_, _00701_);
  nand (_00703_, _23807_, _23316_);
  and (_00704_, _00703_, _00702_);
  and (_00705_, _00704_, _23822_);
  not (_00706_, _00705_);
  nor (_00707_, _00706_, _00700_);
  and (_00708_, _00707_, _23805_);
  not (_00709_, _00708_);
  nor (_00710_, _00709_, _00695_);
  and (_00711_, _00710_, _00694_);
  and (_00712_, _00711_, _00689_);
  nand (_00713_, _00712_, _00685_);
  and (_00714_, _00713_, _00503_);
  and (_00715_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not (_00716_, _24325_);
  and (_00717_, _00716_, _24172_);
  not (_00718_, _24340_);
  and (_00719_, _00507_, _00718_);
  or (_00720_, _00719_, _00717_);
  or (_00721_, _00720_, _00715_);
  or (_00722_, _24517_, _24515_);
  and (_00723_, _24183_, _24518_);
  and (_00724_, _00723_, _00722_);
  or (_00725_, _00724_, _00721_);
  nor (_00726_, _00725_, _00714_);
  nand (_00727_, _00726_, _25762_);
  and (_00728_, _25861_, _25859_);
  nor (_00729_, _00674_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00730_, _00729_, _00728_);
  or (_00731_, _00730_, _25762_);
  and (_00732_, _00731_, _23049_);
  and (_26921_[4], _00732_, _00727_);
  nor (_00733_, _00679_, _24732_);
  nand (_00734_, _24734_, _00733_);
  or (_00735_, _24734_, _00733_);
  nand (_00736_, _00735_, _00734_);
  nand (_00737_, _00736_, _24784_);
  or (_00738_, _24784_, _24725_);
  and (_00739_, _00738_, _00737_);
  nand (_00740_, _00739_, _23752_);
  not (_00741_, _24985_);
  and (_00742_, _00741_, _00686_);
  nor (_00743_, _00742_, _24987_);
  nand (_00744_, _00743_, _24794_);
  nor (_00745_, _25552_, _23602_);
  not (_00746_, _00745_);
  nor (_00747_, _23355_, _23325_);
  nor (_00748_, _00747_, _23582_);
  nor (_00749_, _00748_, _23551_);
  nor (_00750_, _00749_, _23552_);
  and (_00751_, _00750_, _23238_);
  and (_00752_, _23668_, _23316_);
  nor (_00753_, _00752_, _23676_);
  nor (_00754_, _00753_, _25039_);
  and (_00756_, _25039_, _23316_);
  nor (_00757_, _00756_, _00754_);
  nor (_00758_, _00757_, _23679_);
  or (_00759_, _00588_, _23570_);
  nor (_00760_, _23748_, _23348_);
  and (_00761_, _23711_, _23316_);
  nor (_00762_, _00761_, _00760_);
  and (_00763_, _00762_, _00759_);
  and (_00764_, _00763_, _25357_);
  and (_00765_, _00764_, _25354_);
  not (_00766_, _00765_);
  nor (_00767_, _00766_, _00758_);
  and (_00768_, _00767_, _25351_);
  not (_00769_, _00768_);
  nor (_00770_, _00769_, _00751_);
  and (_00771_, _00770_, _00746_);
  and (_00772_, _00771_, _00744_);
  nand (_00773_, _00772_, _00740_);
  and (_00774_, _00773_, _00503_);
  or (_00775_, _24304_, _24305_);
  not (_00776_, _00775_);
  nand (_00777_, _00776_, _24519_);
  or (_00778_, _00776_, _24519_);
  and (_00779_, _00778_, _24183_);
  and (_00780_, _00779_, _00777_);
  and (_00781_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_00782_, _24286_);
  and (_00783_, _00782_, _24172_);
  and (_00784_, _00507_, _25520_);
  or (_00785_, _00784_, _00783_);
  or (_00786_, _00785_, _00781_);
  nor (_00787_, _00786_, _00780_);
  nand (_00788_, _00787_, _25762_);
  or (_00789_, _00788_, _00774_);
  and (_00790_, _00728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00791_, _00728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00793_, _00791_, _00790_);
  or (_00794_, _00793_, _25762_);
  and (_00795_, _00794_, _23049_);
  and (_26921_[5], _00795_, _00789_);
  or (_00796_, _24781_, _24717_);
  nand (_00797_, _00796_, _24786_);
  nand (_00798_, _00797_, _24784_);
  or (_00799_, _24784_, _24710_);
  and (_00800_, _00799_, _00798_);
  nand (_00801_, _00800_, _23752_);
  or (_00802_, _24987_, _24797_);
  and (_00803_, _00802_, _24988_);
  nand (_00804_, _00803_, _24794_);
  nor (_00805_, _25548_, _23602_);
  not (_00806_, _00805_);
  nor (_00807_, _23676_, _23570_);
  not (_00808_, _00807_);
  and (_00809_, _00808_, _25040_);
  not (_00810_, _25039_);
  and (_00811_, _00752_, _24835_);
  nor (_00812_, _00752_, _24835_);
  nor (_00813_, _00812_, _00811_);
  nor (_00814_, _00813_, _00810_);
  or (_00815_, _00814_, _23679_);
  nor (_00816_, _00815_, _00809_);
  not (_00817_, _00816_);
  or (_00818_, _00588_, _23279_);
  and (_00820_, _23711_, _24835_);
  and (_00821_, _23747_, _23316_);
  nor (_00822_, _00821_, _00820_);
  and (_00823_, _00822_, _00818_);
  not (_00824_, _00823_);
  nor (_00825_, _00824_, _25329_);
  and (_00826_, _00825_, _25324_);
  and (_00827_, _00826_, _25320_);
  and (_00828_, _00827_, _00817_);
  nor (_00830_, _23586_, _23552_);
  or (_00831_, _00830_, _00535_);
  or (_00832_, _00831_, _23587_);
  and (_00833_, _00832_, _00828_);
  and (_00834_, _00833_, _00806_);
  and (_00835_, _00834_, _00804_);
  nand (_00836_, _00835_, _00801_);
  and (_00837_, _00836_, _00503_);
  or (_00838_, _24521_, _24268_);
  and (_00839_, _00838_, _24522_);
  and (_00840_, _00839_, _24183_);
  not (_00841_, _24247_);
  and (_00842_, _00841_, _24172_);
  and (_00843_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_00844_, _00507_, _25396_);
  or (_00846_, _00844_, _00843_);
  or (_00847_, _00846_, _00842_);
  or (_00848_, _00847_, _00840_);
  or (_00849_, _00848_, _00837_);
  and (_00850_, _00849_, _25762_);
  and (_00851_, _00790_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00852_, _00790_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00853_, _00852_, _00851_);
  nor (_00854_, _00853_, _25762_);
  or (_00855_, _00854_, _00850_);
  and (_26921_[6], _00855_, _23049_);
  and (_00856_, _00503_, _25053_);
  and (_00857_, _23043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_00858_, _24205_);
  and (_00859_, _00858_, _24172_);
  and (_00860_, _00507_, _25440_);
  or (_00861_, _00860_, _00859_);
  or (_00862_, _00861_, _00857_);
  or (_00863_, _00862_, _00856_);
  or (_00864_, _24225_, _24226_);
  and (_00866_, _00864_, _24523_);
  nor (_00867_, _00864_, _24523_);
  or (_00868_, _00867_, _00866_);
  nand (_00869_, _00868_, _24183_);
  nand (_00870_, _00869_, _25762_);
  or (_00871_, _00870_, _00863_);
  and (_00872_, _25864_, _25859_);
  nor (_00873_, _00851_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00874_, _00873_, _00872_);
  or (_00875_, _00874_, _25762_);
  and (_00876_, _00875_, _23049_);
  and (_26921_[7], _00876_, _00871_);
  and (_00878_, _00500_, _23043_);
  and (_00879_, _24525_, _24541_);
  and (_00880_, _24542_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00881_, _00880_, _00879_);
  nand (_00882_, _00881_, _24534_);
  or (_00883_, _00881_, _24534_);
  and (_00884_, _00883_, _24183_);
  and (_00885_, _00884_, _00882_);
  and (_00886_, _24784_, _23752_);
  or (_00888_, _25810_, _23594_);
  nor (_00890_, _25811_, _00535_);
  and (_00891_, _00890_, _00888_);
  nor (_00893_, _25775_, _23536_);
  nor (_00894_, _25768_, _23710_);
  nor (_00895_, _00894_, _00893_);
  nand (_00896_, _00895_, _23483_);
  or (_00897_, _00895_, _23483_);
  and (_00898_, _00897_, _23744_);
  and (_00899_, _00898_, _00896_);
  and (_00900_, _24836_, _23717_);
  and (_00901_, _00900_, _24794_);
  and (_00902_, _23715_, _23661_);
  and (_00903_, _23711_, _23483_);
  nor (_00904_, _25020_, _23476_);
  or (_00905_, _00904_, _00903_);
  or (_00906_, _00905_, _00902_);
  or (_00907_, _00906_, _00901_);
  or (_00908_, _00907_, _00899_);
  or (_00909_, _00908_, _00891_);
  or (_00910_, _00909_, _00886_);
  and (_00911_, _00910_, _24179_);
  and (_00912_, _00502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00913_, _24499_, _24172_);
  and (_00914_, _00507_, _23928_);
  or (_00915_, _00914_, _00913_);
  nor (_00916_, _00915_, _00912_);
  nand (_00917_, _00916_, _25762_);
  or (_00918_, _00917_, _00911_);
  or (_00919_, _00918_, _00885_);
  or (_00921_, _00919_, _00878_);
  nor (_00922_, _00872_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00924_, _00922_, _25866_);
  or (_00925_, _00924_, _25762_);
  and (_00926_, _00925_, _23049_);
  and (_26921_[8], _00926_, _00921_);
  and (_00927_, _00557_, _23043_);
  or (_00928_, _24526_, _24534_);
  or (_00929_, _24543_, _24224_);
  and (_00930_, _00929_, _00928_);
  nand (_00931_, _00930_, _24540_);
  or (_00932_, _00930_, _24540_);
  and (_00933_, _00932_, _24183_);
  and (_00934_, _00933_, _00931_);
  or (_00935_, _25814_, _25811_);
  nor (_00936_, _25815_, _00535_);
  and (_00937_, _00936_, _00935_);
  and (_00938_, _24685_, _23752_);
  and (_00939_, _25769_, _23536_);
  and (_00940_, _25775_, _23484_);
  and (_00941_, _00940_, _23710_);
  nor (_00942_, _00941_, _00939_);
  nor (_00943_, _00942_, _23454_);
  and (_00944_, _00942_, _23454_);
  or (_00945_, _00944_, _00943_);
  and (_00946_, _00945_, _23744_);
  nor (_00947_, _24884_, _24883_);
  nor (_00948_, _00947_, _24885_);
  and (_00949_, _00948_, _24794_);
  and (_00950_, _23715_, _23316_);
  and (_00951_, _23711_, _23454_);
  and (_00952_, _23742_, _23448_);
  or (_00953_, _00952_, _00951_);
  or (_00955_, _00953_, _00950_);
  or (_00956_, _00955_, _00949_);
  or (_00957_, _00956_, _00946_);
  or (_00958_, _00957_, _00938_);
  or (_00959_, _00958_, _00937_);
  and (_00960_, _00959_, _24179_);
  and (_00961_, _24457_, _24172_);
  and (_00962_, _00502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_00963_, _00507_, _22934_);
  or (_00964_, _00963_, _00962_);
  or (_00965_, _00964_, _00961_);
  nor (_00966_, _00965_, _00960_);
  nand (_00967_, _00966_, _25762_);
  or (_00968_, _00967_, _00934_);
  or (_00969_, _00968_, _00927_);
  nor (_00970_, _25866_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00971_, _00970_, _25867_);
  or (_00973_, _00971_, _25762_);
  and (_00974_, _00973_, _23049_);
  and (_26921_[9], _00974_, _00969_);
  or (_00975_, _24527_, _24534_);
  or (_00976_, _24544_, _24224_);
  and (_00977_, _00976_, _00975_);
  nand (_00978_, _00977_, _24539_);
  or (_00979_, _00977_, _24539_);
  and (_00980_, _00979_, _00978_);
  and (_00981_, _00980_, _24183_);
  and (_00982_, _00609_, _23043_);
  not (_00983_, _24179_);
  nor (_00984_, _25818_, _25815_);
  nor (_00985_, _00984_, _25819_);
  and (_00986_, _00985_, _23238_);
  not (_00987_, _00986_);
  and (_00988_, _00940_, _23624_);
  and (_00989_, _00988_, _23710_);
  and (_00990_, _25770_, _23536_);
  nor (_00991_, _00990_, _00989_);
  and (_00993_, _00991_, _23628_);
  nor (_00994_, _00991_, _23628_);
  or (_00995_, _00994_, _25311_);
  nor (_00996_, _00995_, _00993_);
  nor (_00997_, _24961_, _24959_);
  nor (_00998_, _00997_, _24962_);
  and (_00999_, _00998_, _24794_);
  and (_01000_, _23711_, _23419_);
  and (_01001_, _23715_, _24835_);
  and (_01002_, _23742_, _23412_);
  and (_01004_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_01005_, _01004_, _01002_);
  or (_01006_, _01005_, _01001_);
  nor (_01007_, _01006_, _01000_);
  not (_01008_, _01007_);
  nor (_01009_, _01008_, _00999_);
  not (_01010_, _01009_);
  nor (_01011_, _01010_, _00996_);
  and (_01012_, _01011_, _00987_);
  nor (_01014_, _01012_, _00983_);
  and (_01015_, _24418_, _24172_);
  and (_01016_, _00502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01017_, _00507_, _22909_);
  or (_01018_, _01017_, _01016_);
  or (_01019_, _01018_, _01015_);
  nor (_01020_, _01019_, _01014_);
  nand (_01021_, _01020_, _25762_);
  or (_01022_, _01021_, _00982_);
  or (_01023_, _01022_, _00981_);
  nor (_01024_, _25867_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01025_, _01024_, _25868_);
  or (_01026_, _01025_, _25762_);
  and (_01027_, _01026_, _23049_);
  and (_26921_[10], _01027_, _01023_);
  or (_01028_, _24545_, _24224_);
  or (_01029_, _24528_, _24534_);
  and (_01030_, _01029_, _01028_);
  nand (_01031_, _01030_, _24538_);
  or (_01032_, _01030_, _24538_);
  and (_01033_, _01032_, _01031_);
  and (_01034_, _01033_, _24183_);
  and (_01035_, _25849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01036_, _00659_, _23043_);
  or (_01037_, _25819_, _25807_);
  nor (_01038_, _25820_, _00535_);
  and (_01039_, _01038_, _01037_);
  or (_01040_, _24964_, _24962_);
  and (_01041_, _01040_, _24965_);
  and (_01042_, _01041_, _24794_);
  and (_01043_, _25771_, _23536_);
  and (_01044_, _00988_, _23628_);
  and (_01045_, _01044_, _23710_);
  nor (_01046_, _01045_, _01043_);
  nand (_01047_, _01046_, _23384_);
  or (_01048_, _01046_, _23384_);
  and (_01049_, _01048_, _23744_);
  and (_01050_, _01049_, _01047_);
  nor (_01051_, _25020_, _23378_);
  and (_01052_, _23711_, _23647_);
  and (_01053_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_01054_, _01053_, _01052_);
  or (_01055_, _01054_, _23716_);
  or (_01056_, _01055_, _01051_);
  or (_01057_, _01056_, _01050_);
  or (_01058_, _01057_, _01042_);
  or (_01059_, _01058_, _01039_);
  and (_01060_, _01059_, _24179_);
  and (_01061_, _25214_, _24172_);
  or (_01062_, _01061_, _01060_);
  or (_01063_, _01062_, _01036_);
  nor (_01064_, _01063_, _01035_);
  nand (_01065_, _01064_, _25762_);
  or (_01066_, _01065_, _01034_);
  nor (_01067_, _25868_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01068_, _01067_, _25869_);
  or (_01070_, _01068_, _25762_);
  and (_01071_, _01070_, _23049_);
  and (_26921_[11], _01071_, _01066_);
  or (_01073_, _24529_, _24534_);
  or (_01074_, _24546_, _24224_);
  and (_01075_, _01074_, _01073_);
  nand (_01076_, _01075_, _24537_);
  or (_01077_, _01075_, _24537_);
  and (_01078_, _01077_, _01076_);
  and (_01079_, _01078_, _24183_);
  and (_01080_, _00713_, _23043_);
  or (_01081_, _25824_, _25820_);
  and (_01082_, _25825_, _23238_);
  and (_01083_, _01082_, _01081_);
  or (_01085_, _24968_, _24966_);
  and (_01086_, _01085_, _24969_);
  and (_01087_, _01086_, _24794_);
  and (_01088_, _25779_, _23710_);
  nor (_01089_, _01088_, _25773_);
  nand (_01090_, _01089_, _23354_);
  or (_01091_, _01089_, _23354_);
  and (_01092_, _01091_, _01090_);
  and (_01093_, _01092_, _23744_);
  or (_01095_, _23536_, _23661_);
  nor (_01096_, _25784_, _25020_);
  and (_01097_, _01096_, _01095_);
  and (_01098_, _23715_, _23717_);
  and (_01099_, _23711_, _23609_);
  and (_01101_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_01102_, _01101_, _01099_);
  or (_01103_, _01102_, _01098_);
  or (_01105_, _01103_, _01097_);
  or (_01106_, _01105_, _01093_);
  or (_01108_, _01106_, _01087_);
  or (_01109_, _01108_, _01083_);
  and (_01110_, _01109_, _24179_);
  and (_01111_, _00718_, _24172_);
  and (_01112_, _25849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01113_, _01112_, _01111_);
  nor (_01114_, _01113_, _01110_);
  nand (_01115_, _01114_, _25762_);
  or (_01116_, _01115_, _01080_);
  or (_01117_, _01116_, _01079_);
  nor (_01118_, _25869_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01120_, _01118_, _25870_);
  or (_01121_, _01120_, _25762_);
  and (_01122_, _01121_, _23049_);
  and (_26921_[12], _01122_, _01117_);
  or (_01123_, _24530_, _24534_);
  or (_01124_, _24547_, _24224_);
  and (_01125_, _01124_, _01123_);
  nor (_01126_, _01125_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01127_, _01125_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01128_, _01127_, _01126_);
  and (_01129_, _01128_, _24183_);
  and (_01130_, _00773_, _23043_);
  and (_01131_, _25825_, _25804_);
  not (_01132_, _01131_);
  and (_01133_, _25826_, _23238_);
  and (_01134_, _01133_, _01132_);
  not (_01135_, _01134_);
  or (_01136_, _24970_, _24948_);
  and (_01137_, _01136_, _24971_);
  and (_01138_, _01137_, _24794_);
  nor (_01139_, _25780_, _25773_);
  nor (_01140_, _01139_, _25784_);
  and (_01141_, _01140_, _23607_);
  nor (_01142_, _01140_, _23607_);
  nor (_01143_, _01142_, _01141_);
  nor (_01144_, _01143_, _25311_);
  and (_01145_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  not (_01146_, _25783_);
  nor (_01148_, _23536_, _23316_);
  nor (_01149_, _01148_, _25020_);
  and (_01150_, _01149_, _01146_);
  and (_01151_, _23715_, _23448_);
  and (_01152_, _23711_, _23322_);
  or (_01153_, _01152_, _01151_);
  or (_01154_, _01153_, _01150_);
  nor (_01155_, _01154_, _01145_);
  not (_01156_, _01155_);
  nor (_01157_, _01156_, _01144_);
  not (_01158_, _01157_);
  nor (_01159_, _01158_, _01138_);
  and (_01160_, _01159_, _01135_);
  nor (_01161_, _01160_, _00983_);
  and (_01162_, _25520_, _24172_);
  or (_01163_, _01162_, _01161_);
  or (_01164_, _01163_, _01130_);
  or (_01165_, _01164_, _01129_);
  nand (_01166_, _25849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_01167_, _01166_, _25762_);
  or (_01168_, _01167_, _01165_);
  nor (_01169_, _25870_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01170_, _01169_, _25871_);
  or (_01171_, _01170_, _25762_);
  and (_01172_, _01171_, _23049_);
  and (_26921_[13], _01172_, _01168_);
  nand (_01173_, _24548_, _24534_);
  nand (_01174_, _24531_, _24224_);
  and (_01175_, _01174_, _01173_);
  nor (_01176_, _01175_, _24535_);
  and (_01177_, _01175_, _24535_);
  or (_01178_, _01177_, _01176_);
  and (_01179_, _01178_, _24183_);
  and (_01180_, _00836_, _23043_);
  and (_01181_, _23711_, _23576_);
  and (_01182_, _23715_, _23412_);
  and (_01183_, _25786_, _23577_);
  nor (_01184_, _25786_, _23577_);
  nor (_01185_, _01184_, _01183_);
  nor (_01186_, _01185_, _25311_);
  nor (_01187_, _24835_, _23536_);
  not (_01188_, _01187_);
  nor (_01189_, _25788_, _25020_);
  and (_01190_, _01189_, _01188_);
  or (_01191_, _01190_, _01186_);
  or (_01192_, _01191_, _01182_);
  and (_01193_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  and (_01194_, _25830_, _25826_);
  not (_01195_, _01194_);
  and (_01196_, _25831_, _23238_);
  and (_01197_, _01196_, _01195_);
  or (_01198_, _24972_, _24942_);
  and (_01199_, _01198_, _24973_);
  and (_01200_, _01199_, _24794_);
  or (_01201_, _01200_, _01197_);
  or (_01202_, _01201_, _01193_);
  or (_01203_, _01202_, _01192_);
  or (_01204_, _01203_, _01181_);
  and (_01205_, _01204_, _24179_);
  and (_01206_, _25396_, _24172_);
  and (_01207_, _25849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01208_, _01207_, _01206_);
  or (_01209_, _01208_, _01205_);
  or (_01210_, _01209_, _01180_);
  or (_01211_, _01210_, _01179_);
  or (_01212_, _01211_, _00517_);
  nor (_01213_, _25871_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01214_, _01213_, _25872_);
  or (_01215_, _01214_, _25762_);
  and (_01216_, _01215_, _23049_);
  and (_26921_[14], _01216_, _01212_);
  and (_01217_, _00428_, _23830_);
  and (_01218_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_22619_, _01218_, _01217_);
  or (_01219_, _24093_, _24091_);
  nor (_01220_, _23856_, _24094_);
  and (_01221_, _01220_, _01219_);
  and (_01222_, _23856_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_01223_, _01222_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01224_, _01223_, _01221_);
  or (_01226_, _23841_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_01227_, _01226_, _23049_);
  and (_26922_[0], _01227_, _01224_);
  nor (_01228_, _24096_, _24094_);
  nor (_01229_, _01228_, _24097_);
  or (_01230_, _01229_, _23856_);
  or (_01231_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01232_, _01231_, _23841_);
  and (_01233_, _01232_, _01230_);
  and (_01234_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_01235_, _01234_, _01233_);
  and (_26922_[1], _01235_, _23049_);
  nor (_01236_, _24101_, _24099_);
  nor (_01237_, _01236_, _24102_);
  or (_01238_, _01237_, _23856_);
  or (_01239_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01240_, _01239_, _23841_);
  and (_01241_, _01240_, _01238_);
  and (_01242_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_01243_, _01242_, _01241_);
  and (_26922_[2], _01243_, _23049_);
  nor (_01244_, _24102_, _23920_);
  nor (_01246_, _01244_, _24103_);
  or (_01247_, _01246_, _23856_);
  or (_01248_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01249_, _01248_, _24135_);
  and (_01250_, _01249_, _01247_);
  and (_01251_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _23049_);
  and (_01252_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_26922_[3], _01252_, _01250_);
  nor (_01253_, _24106_, _24103_);
  nor (_01255_, _01253_, _24107_);
  or (_01256_, _01255_, _23856_);
  or (_01257_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01258_, _01257_, _24135_);
  and (_01260_, _01258_, _01256_);
  and (_01261_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_26922_[4], _01261_, _01260_);
  or (_01262_, _24107_, _23914_);
  nor (_01263_, _23856_, _24108_);
  and (_01264_, _01263_, _01262_);
  nor (_01265_, _23855_, _23298_);
  or (_01266_, _01265_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01267_, _01266_, _01264_);
  or (_01268_, _23841_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01269_, _01268_, _23049_);
  and (_26922_[5], _01269_, _01267_);
  and (_01270_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_01272_, _24108_, _23911_);
  nor (_01273_, _01272_, _24109_);
  or (_01274_, _01273_, _23856_);
  or (_01275_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01276_, _01275_, _24135_);
  and (_01277_, _01276_, _01274_);
  or (_26922_[6], _01277_, _01270_);
  or (_01278_, _24109_, _23908_);
  nor (_01279_, _23856_, _24110_);
  and (_01280_, _01279_, _01278_);
  nor (_01281_, _23855_, _23239_);
  or (_01282_, _01281_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01283_, _01282_, _01280_);
  or (_01284_, _23841_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_01285_, _01284_, _23049_);
  and (_26922_[7], _01285_, _01283_);
  and (_01286_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_01287_, _24113_, _24110_);
  nor (_01288_, _01287_, _24114_);
  or (_01289_, _01288_, _23856_);
  or (_01290_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01291_, _01290_, _24135_);
  and (_01292_, _01291_, _01289_);
  or (_26922_[8], _01292_, _01286_);
  nor (_01293_, _24114_, _23905_);
  nor (_01294_, _01293_, _24115_);
  or (_01295_, _01294_, _23856_);
  or (_01296_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_01297_, _01296_, _24135_);
  and (_01298_, _01297_, _01295_);
  and (_01299_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_26922_[9], _01299_, _01298_);
  nor (_01300_, _24115_, _23899_);
  nor (_01301_, _01300_, _24116_);
  or (_01302_, _01301_, _23856_);
  or (_01303_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01304_, _01303_, _24135_);
  and (_01305_, _01304_, _01302_);
  and (_01306_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_26922_[10], _01306_, _01305_);
  nor (_01307_, _24116_, _23897_);
  nor (_01308_, _01307_, _24117_);
  or (_01309_, _01308_, _23856_);
  or (_01310_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01311_, _01310_, _24135_);
  and (_01312_, _01311_, _01309_);
  and (_01313_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_26922_[11], _01313_, _01312_);
  nor (_01314_, _24119_, _24117_);
  nor (_01315_, _01314_, _24120_);
  or (_01316_, _01315_, _23856_);
  or (_01317_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01318_, _01317_, _24135_);
  and (_01319_, _01318_, _01316_);
  and (_01320_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_26922_[12], _01320_, _01319_);
  and (_01321_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01322_, _24120_, _23891_);
  nor (_01323_, _01322_, _24121_);
  or (_01324_, _01323_, _23856_);
  or (_01326_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01327_, _01326_, _24135_);
  and (_01328_, _01327_, _01324_);
  or (_26922_[13], _01328_, _01321_);
  nor (_01329_, _24125_, _24121_);
  nor (_01330_, _01329_, _24126_);
  or (_01331_, _01330_, _23856_);
  or (_01332_, _23855_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01333_, _01332_, _24135_);
  and (_01334_, _01333_, _01331_);
  and (_01335_, _01251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_26922_[14], _01335_, _01334_);
  and (_01336_, _00428_, _26185_);
  and (_01337_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_27225_, _01337_, _01336_);
  and (_01338_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01339_, _01338_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_26926_[0], _01339_, _23049_);
  and (_01340_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01341_, _01340_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_26926_[1], _01341_, _23049_);
  and (_01342_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_01343_, _01342_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_26926_[2], _01343_, _23049_);
  and (_01344_, _23839_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01345_, _01344_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_26926_[3], _01345_, _23049_);
  and (_01346_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01347_, _01346_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26926_[4], _01347_, _23049_);
  and (_01348_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01349_, _01348_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_26926_[5], _01349_, _23049_);
  and (_01350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _23049_);
  and (_01351_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _23049_);
  and (_01352_, _01351_, _23840_);
  or (_26926_[6], _01352_, _01350_);
  nor (_01353_, _24089_, _24307_);
  nand (_01354_, _01353_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_01355_, _01353_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_01356_, _01355_, _24135_);
  and (_26927_[0], _01356_, _01354_);
  and (_01357_, _24091_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_01358_, _24073_, _22749_);
  and (_01359_, _24073_, _22749_);
  nor (_01360_, _01359_, _01358_);
  and (_01361_, _01360_, _01357_);
  nor (_01362_, _01360_, _01357_);
  nor (_01363_, _01362_, _01361_);
  or (_01364_, _01363_, _24307_);
  or (_01365_, _22739_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01366_, _01365_, _24135_);
  and (_26927_[1], _01366_, _01364_);
  and (_01367_, _25932_, _23230_);
  and (_01368_, _01367_, _25927_);
  not (_01369_, _01367_);
  and (_01370_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_27226_, _01370_, _01368_);
  and (_01371_, _26190_, _25938_);
  and (_01372_, _01371_, _25927_);
  not (_01373_, _01371_);
  and (_01374_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_27233_, _01374_, _01372_);
  and (_01375_, _01367_, _25886_);
  and (_01376_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_27227_, _01376_, _01375_);
  and (_01378_, _01367_, _26085_);
  and (_01379_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_27228_, _01379_, _01378_);
  and (_01380_, _01367_, _26242_);
  and (_01381_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_27230_, _01381_, _01380_);
  and (_01383_, _26073_, _23768_);
  and (_01384_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_27231_, _01384_, _01383_);
  nor (_01386_, _00404_, _26474_);
  nand (_01387_, _01386_, _23729_);
  or (_01388_, _01386_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01389_, _01388_, _25618_);
  and (_01390_, _01389_, _01387_);
  nand (_01391_, _00410_, _25160_);
  or (_01392_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01393_, _01392_, _25128_);
  and (_01394_, _01393_, _01391_);
  and (_01395_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_01396_, _01395_, rst);
  or (_01397_, _01396_, _01394_);
  or (_22620_, _01397_, _01390_);
  nor (_01398_, _00404_, _25895_);
  nand (_01399_, _01398_, _23729_);
  or (_01400_, _01398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_01401_, _01400_, _25618_);
  and (_01402_, _01401_, _01399_);
  not (_01403_, _00410_);
  or (_01404_, _01403_, _25258_);
  or (_01405_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_01406_, _01405_, _25128_);
  and (_01407_, _01406_, _01404_);
  and (_01408_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_01409_, _01408_, rst);
  or (_01410_, _01409_, _01407_);
  or (_22621_, _01410_, _01402_);
  not (_01411_, _25224_);
  nor (_01413_, _00404_, _01411_);
  nand (_01414_, _01413_, _23729_);
  or (_01415_, _01413_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01416_, _01415_, _25618_);
  and (_01417_, _01416_, _01414_);
  nand (_01418_, _00410_, _25279_);
  or (_01419_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01420_, _01419_, _25128_);
  and (_01421_, _01420_, _01418_);
  and (_01422_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_01423_, _01422_, rst);
  or (_01424_, _01423_, _01421_);
  or (_22622_, _01424_, _01417_);
  not (_01425_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_01426_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _01425_);
  and (_01427_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01428_, _01427_, _01426_);
  and (_26931_[0], _01428_, _23049_);
  and (_01429_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _01425_);
  and (_01430_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01431_, _01430_, _01429_);
  and (_26931_[1], _01431_, _23049_);
  and (_01432_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _01425_);
  and (_01433_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01435_, _01433_, _01432_);
  and (_26931_[2], _01435_, _23049_);
  and (_01436_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _01425_);
  and (_01437_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01438_, _01437_, _01436_);
  and (_26931_[3], _01438_, _23049_);
  and (_01439_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _01425_);
  and (_01440_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01441_, _01440_, _01439_);
  and (_26931_[4], _01441_, _23049_);
  and (_01442_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _01425_);
  and (_01443_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01444_, _01443_, _01442_);
  and (_26931_[5], _01444_, _23049_);
  and (_01445_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _01425_);
  and (_01446_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01447_, _01446_, _01445_);
  and (_26931_[6], _01447_, _23049_);
  not (_01448_, _25131_);
  nor (_01449_, _00404_, _01448_);
  nand (_01450_, _01449_, _23729_);
  or (_01451_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_01452_, _01451_, _25618_);
  and (_01453_, _01452_, _01450_);
  nand (_01454_, _00410_, _23761_);
  and (_01455_, _01454_, _25128_);
  and (_01456_, _01455_, _01451_);
  not (_01457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_01458_, _25127_, _01457_);
  or (_01459_, _01458_, rst);
  or (_01460_, _01459_, _01456_);
  or (_22623_, _01460_, _01453_);
  and (_26934_[0], _00465_, _23049_);
  nor (_26934_[1], _00470_, rst);
  and (_26934_[2], _00473_, _23049_);
  and (_01461_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_01462_, _25858_, _22815_);
  or (_01463_, _01462_, _01461_);
  and (_26936_[0], _01463_, _23049_);
  and (_01464_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_01465_, _25858_, _22837_);
  or (_01466_, _01465_, _01464_);
  and (_26936_[1], _01466_, _23049_);
  and (_01467_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_01468_, _25858_, _22758_);
  or (_01469_, _01468_, _01467_);
  and (_26936_[2], _01469_, _23049_);
  and (_01470_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_01471_, _25858_, _22794_);
  or (_01472_, _01471_, _01470_);
  and (_26936_[3], _01472_, _23049_);
  and (_01473_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_01474_, _25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_01475_, _01474_, _01473_);
  and (_26936_[4], _01475_, _23049_);
  and (_01476_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_01477_, _25858_, _22875_);
  or (_01478_, _01477_, _01476_);
  and (_26936_[5], _01478_, _23049_);
  and (_01479_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_01480_, _25858_, _22914_);
  or (_01481_, _01480_, _01479_);
  and (_26936_[6], _01481_, _23049_);
  and (_01482_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_01483_, _25858_, _22901_);
  or (_01484_, _01483_, _01482_);
  and (_26936_[7], _01484_, _23049_);
  and (_01485_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_01486_, _25858_, _24465_);
  or (_01487_, _01486_, _01485_);
  and (_26936_[8], _01487_, _23049_);
  and (_01488_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01489_, _25858_, _24425_);
  or (_01490_, _01489_, _01488_);
  and (_26936_[9], _01490_, _23049_);
  and (_01491_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_01492_, _25858_, _24390_);
  or (_01493_, _01492_, _01491_);
  and (_26936_[10], _01493_, _23049_);
  and (_01494_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01495_, _25858_, _24346_);
  or (_01496_, _01495_, _01494_);
  and (_26936_[11], _01496_, _23049_);
  and (_01497_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_01498_, _25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_01499_, _01498_, _01497_);
  and (_26936_[12], _01499_, _23049_);
  and (_01500_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_01501_, _25858_, _24278_);
  or (_01503_, _01501_, _01500_);
  and (_26936_[13], _01503_, _23049_);
  and (_01506_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_01507_, _25858_, _24235_);
  or (_01509_, _01507_, _01506_);
  and (_26936_[14], _01509_, _23049_);
  and (_01511_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_01512_, _25858_, _24188_);
  or (_01513_, _01512_, _01511_);
  and (_26936_[15], _01513_, _23049_);
  or (_01514_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_01515_, _25858_, _22811_);
  and (_01516_, _01515_, _23049_);
  and (_26936_[16], _01516_, _01514_);
  and (_01517_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_01518_, _25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_01519_, _01518_, _01517_);
  and (_26936_[17], _01519_, _23049_);
  or (_01521_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_01522_, _25858_, _22765_);
  and (_01523_, _01522_, _23049_);
  and (_26936_[18], _01523_, _01521_);
  or (_01525_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_01526_, _25858_, _22788_);
  and (_01527_, _01526_, _23049_);
  and (_26936_[19], _01527_, _01525_);
  and (_01528_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_01530_, _25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_01531_, _01530_, _01528_);
  and (_26936_[20], _01531_, _23049_);
  or (_01532_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_01533_, _25858_, _22871_);
  and (_01534_, _01533_, _23049_);
  and (_26936_[21], _01534_, _01532_);
  or (_01535_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_01536_, _25858_, _22921_);
  and (_01537_, _01536_, _23049_);
  and (_26936_[22], _01537_, _01535_);
  or (_01538_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_01539_, _25858_, _22897_);
  and (_01540_, _01539_, _23049_);
  and (_26936_[23], _01540_, _01538_);
  or (_01541_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_01542_, _25858_, _22819_);
  and (_01543_, _01542_, _23049_);
  and (_26936_[24], _01543_, _01541_);
  or (_01544_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_01545_, _25858_, _22839_);
  and (_01546_, _01545_, _23049_);
  and (_26936_[25], _01546_, _01544_);
  or (_01547_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_01548_, _25858_, _22744_);
  and (_01549_, _01548_, _23049_);
  and (_26936_[26], _01549_, _01547_);
  or (_01550_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_01551_, _25858_, _22785_);
  and (_01552_, _01551_, _23049_);
  and (_26936_[27], _01552_, _01550_);
  and (_01553_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_01554_, _25859_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_01555_, _01554_, _01553_);
  and (_26936_[28], _01555_, _23049_);
  or (_01556_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_01557_, _25858_, _22868_);
  and (_01558_, _01557_, _23049_);
  and (_26936_[29], _01558_, _01556_);
  or (_01559_, _25858_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_01560_, _25858_, _22919_);
  and (_01561_, _01560_, _23049_);
  and (_26936_[30], _01561_, _01559_);
  and (_01562_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_01563_, _00141_, _25886_);
  or (_27051_, _01563_, _01562_);
  and (_01564_, _00095_, _26421_);
  and (_01565_, _01564_, _25927_);
  not (_01566_, _01564_);
  and (_01567_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_22624_, _01567_, _01565_);
  and (_01568_, _25938_, _23775_);
  and (_01569_, _01568_, _26085_);
  not (_01570_, _01568_);
  and (_01571_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_22625_, _01571_, _01569_);
  and (_01572_, _01564_, _23768_);
  and (_01573_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_26969_, _01573_, _01572_);
  nand (_01574_, _25627_, _26619_);
  nor (_01575_, _01574_, _01448_);
  nand (_01576_, _01575_, _23729_);
  and (_01577_, _25134_, _23777_);
  and (_01578_, _01577_, _00255_);
  or (_01579_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01580_, _01579_, _25618_);
  and (_01581_, _01580_, _01576_);
  nand (_01582_, _01578_, _23761_);
  and (_01583_, _01582_, _25128_);
  and (_01584_, _01583_, _01579_);
  not (_01585_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_01586_, _25127_, _01585_);
  or (_01587_, _01586_, rst);
  or (_01588_, _01587_, _01584_);
  or (_22626_, _01588_, _01581_);
  not (_01589_, _00449_);
  or (_01590_, _00500_, _01589_);
  or (_01591_, _00449_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_01592_, _01591_, _23049_);
  and (_26940_[0], _01592_, _01590_);
  or (_01593_, _00557_, _01589_);
  or (_01594_, _00449_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_01595_, _01594_, _23049_);
  and (_26940_[1], _01595_, _01593_);
  nand (_01596_, _00608_, _00449_);
  or (_01597_, _00449_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_01598_, _01597_, _23049_);
  and (_26940_[2], _01598_, _01596_);
  or (_01599_, _00659_, _01589_);
  or (_01600_, _00449_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_01601_, _01600_, _23049_);
  and (_26940_[3], _01601_, _01599_);
  and (_01602_, _26351_, _26242_);
  and (_01603_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_22627_, _01603_, _01602_);
  and (_01604_, _26213_, _25938_);
  and (_01605_, _01604_, _26085_);
  not (_01606_, _01604_);
  and (_01607_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_22628_, _01607_, _01605_);
  and (_01608_, _26260_, _23847_);
  not (_01609_, _01608_);
  and (_01610_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_01611_, _01608_, _23830_);
  or (_27165_, _01611_, _01610_);
  not (_01612_, _00190_);
  or (_01613_, _01612_, _25258_);
  and (_01614_, _00209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_01615_, _01614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_01616_, _01615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_01617_, _01615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_01618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_01619_, _01618_, _01617_);
  and (_01620_, _01619_, _01616_);
  and (_01621_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_01622_, _01621_, _01620_);
  nor (_01624_, _01622_, _00226_);
  nor (_01625_, _01618_, _00226_);
  not (_01627_, _01625_);
  and (_01628_, _01627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_01629_, _01628_, _01624_);
  or (_01630_, _01629_, _00190_);
  and (_01631_, _01630_, _23049_);
  and (_22629_, _01631_, _01613_);
  nor (_01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_01633_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _23049_);
  and (_01635_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_22630_, _01635_, _01633_);
  and (_01636_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_01637_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_22631_, _01637_, _01636_);
  and (_01638_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_01639_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_22632_, _01639_, _01638_);
  and (_01640_, _26242_, _23231_);
  and (_01641_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_22633_, _01641_, _01640_);
  and (_01642_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_01643_, _00141_, _26170_);
  or (_22634_, _01643_, _01642_);
  and (_01644_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_01645_, _00141_, _25927_);
  or (_22635_, _01645_, _01644_);
  not (_01646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_01647_, t0_i);
  and (_01648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01647_);
  nor (_01649_, _01648_, _01646_);
  not (_01650_, _01649_);
  not (_01651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_01652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_01653_, _01652_, _01651_);
  and (_01654_, _01653_, _01650_);
  and (_01655_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_01656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_01657_, _01656_, _01655_);
  and (_01658_, _01657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01659_, _01658_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_01660_, _01659_, _01654_);
  nand (_01661_, _01660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_01662_, _01661_, _00071_);
  or (_01663_, _01662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nor (_01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01665_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_01666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_01667_, _01666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_01668_, _01667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01670_, _01669_, _01660_);
  nand (_01671_, _01670_, _01668_);
  and (_01672_, _01666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_01673_, _01672_, _01667_);
  not (_01674_, _00074_);
  nor (_01675_, _01670_, _01674_);
  or (_01676_, _01675_, _01673_);
  and (_01677_, _01676_, _01671_);
  or (_01678_, _01677_, _01665_);
  or (_01679_, _01678_, _00071_);
  and (_01680_, _01679_, _00070_);
  and (_01681_, _01680_, _01663_);
  nor (_01682_, _00070_, _25417_);
  or (_01683_, _01682_, _01681_);
  and (_22636_, _01683_, _23049_);
  and (_01684_, _00096_, _26170_);
  and (_01685_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_22637_, _01685_, _01684_);
  not (_01686_, _26136_);
  nor (_01687_, _01574_, _01686_);
  nand (_01688_, _01687_, _23729_);
  or (_01689_, _01687_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01690_, _01689_, _25618_);
  and (_01691_, _01690_, _01688_);
  nand (_01692_, _01578_, _25362_);
  or (_01693_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01694_, _01693_, _25128_);
  and (_01695_, _01694_, _01692_);
  and (_01696_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_01697_, _01696_, rst);
  or (_01698_, _01697_, _01695_);
  or (_22638_, _01698_, _01691_);
  nor (_01699_, _01574_, _26556_);
  nand (_01700_, _01699_, _23729_);
  or (_01701_, _01699_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01702_, _01701_, _25618_);
  and (_01703_, _01702_, _01700_);
  nand (_01704_, _01578_, _23824_);
  or (_01705_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01706_, _01705_, _25128_);
  and (_01707_, _01706_, _01704_);
  and (_01708_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_01709_, _01708_, rst);
  or (_01710_, _01709_, _01707_);
  or (_22639_, _01710_, _01703_);
  nor (_01711_, _01574_, _26474_);
  nand (_01712_, _01711_, _23729_);
  or (_01713_, _01711_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_01714_, _01713_, _25618_);
  and (_01715_, _01714_, _01712_);
  nand (_01716_, _01578_, _25160_);
  or (_01717_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_01718_, _01717_, _25128_);
  and (_01719_, _01718_, _01716_);
  and (_01720_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_01721_, _01720_, rst);
  or (_01722_, _01721_, _01719_);
  or (_22640_, _01722_, _01715_);
  and (_01723_, _00096_, _25927_);
  and (_01724_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_27324_, _01724_, _01723_);
  nor (_01725_, _01574_, _25895_);
  nand (_01726_, _01725_, _23729_);
  or (_01727_, _01725_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01728_, _01727_, _25618_);
  and (_01729_, _01728_, _01726_);
  not (_01730_, _01578_);
  or (_01731_, _01730_, _25258_);
  or (_01732_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01733_, _01732_, _25128_);
  and (_01734_, _01733_, _01731_);
  and (_01735_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_01736_, _01735_, rst);
  or (_01737_, _01736_, _01734_);
  or (_22641_, _01737_, _01729_);
  and (_01738_, _00096_, _23768_);
  and (_01739_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_22642_, _01739_, _01738_);
  and (_22643_, _01350_, _26657_);
  and (_01740_, _26657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01741_, _01740_, _26734_);
  and (_22644_, _01741_, _23049_);
  and (_01742_, _26690_, _26736_);
  and (_01743_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _26660_);
  and (_01744_, _26686_, _26683_);
  or (_01745_, _01744_, _26677_);
  and (_01746_, _01745_, _01743_);
  or (_01747_, _26797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01748_, _26800_, _26683_);
  and (_01749_, _01748_, _01747_);
  not (_01750_, _26683_);
  or (_01751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01752_, _01751_, _01750_);
  or (_01753_, _01752_, _01749_);
  and (_01754_, _01753_, _26678_);
  or (_01755_, _01754_, _01746_);
  and (_01756_, _01755_, _01742_);
  not (_01757_, _26713_);
  or (_01758_, _01757_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_01759_, _26816_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01760_, _01759_, _26819_);
  nand (_01761_, _01743_, _26700_);
  nand (_01763_, _01761_, _26710_);
  or (_01764_, _01763_, _01760_);
  or (_01765_, _01751_, _26710_);
  and (_01767_, _01765_, _26706_);
  and (_01768_, _01767_, _01764_);
  and (_01769_, _01743_, _26705_);
  or (_01770_, _01769_, _26713_);
  or (_01771_, _01770_, _01768_);
  and (_01772_, _01771_, _26732_);
  or (_01773_, _01772_, _26657_);
  and (_01774_, _01773_, _01758_);
  or (_01775_, _01774_, _01756_);
  and (_22645_, _01775_, _23049_);
  and (_01776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01777_, _01776_, _01745_);
  or (_01778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _26660_);
  or (_01779_, _01778_, _26683_);
  and (_01780_, _01779_, _26678_);
  or (_01781_, _26737_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01782_, _01781_, _26740_);
  or (_01783_, _01782_, _01750_);
  and (_01784_, _01783_, _01780_);
  or (_01785_, _01784_, _01777_);
  and (_01786_, _01785_, _01742_);
  or (_01787_, _01757_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_01788_, _01778_, _26710_);
  and (_01789_, _01788_, _26706_);
  or (_01790_, _26759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01791_, _01790_, _26762_);
  nand (_01792_, _01776_, _26700_);
  nand (_01793_, _01792_, _26710_);
  or (_01794_, _01793_, _01791_);
  and (_01795_, _01794_, _01789_);
  and (_01796_, _01776_, _26705_);
  or (_01797_, _01796_, _26713_);
  or (_01798_, _01797_, _01795_);
  and (_01799_, _01798_, _26732_);
  or (_01800_, _01799_, _26657_);
  and (_01801_, _01800_, _01787_);
  or (_01802_, _01801_, _01786_);
  and (_22646_, _01802_, _23049_);
  and (_01803_, _26548_, _26136_);
  nand (_01804_, _01803_, _23729_);
  or (_01805_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01806_, _01805_, _26547_);
  and (_01807_, _01806_, _01804_);
  nor (_01808_, _26547_, _25362_);
  or (_01809_, _01808_, _01807_);
  and (_22647_, _01809_, _23049_);
  and (_01810_, _26558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01811_, _01810_, _26557_);
  and (_01812_, _01811_, _26472_);
  not (_01813_, _26472_);
  or (_01814_, _26564_, _01813_);
  and (_01815_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01816_, _01815_, _26485_);
  or (_01817_, _01816_, _01812_);
  nand (_01818_, _26485_, _23824_);
  and (_01819_, _01818_, _23049_);
  and (_22648_, _01819_, _01817_);
  and (_01820_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_01821_, _26422_, _23830_);
  or (_22649_, _01821_, _01820_);
  and (_01822_, _26294_, _23830_);
  and (_01823_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_22650_, _01823_, _01822_);
  and (_01824_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_01825_, _26185_, _23780_);
  or (_22651_, _01825_, _01824_);
  and (_01826_, _25616_, _26619_);
  nand (_01827_, _25905_, _01826_);
  and (_01828_, _01827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_01829_, _25223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_01830_, _01829_, _25896_);
  and (_01831_, _01830_, _01826_);
  or (_01832_, _01831_, _01828_);
  and (_01833_, _01832_, _25618_);
  and (_01834_, _00255_, _25226_);
  not (_01835_, _01834_);
  or (_01836_, _01835_, _25258_);
  or (_01837_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_01838_, _01837_, _25128_);
  and (_01839_, _01838_, _01836_);
  and (_01840_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_01841_, _01840_, rst);
  or (_01842_, _01841_, _01839_);
  or (_22652_, _01842_, _01833_);
  and (_01843_, _25224_, _23153_);
  and (_01844_, _01843_, _25226_);
  nand (_01845_, _01844_, _23729_);
  or (_01846_, _01844_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01847_, _01846_, _25618_);
  and (_01848_, _01847_, _01845_);
  nand (_01849_, _01834_, _25279_);
  or (_01850_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01851_, _01850_, _25128_);
  and (_01852_, _01851_, _01849_);
  and (_01853_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_01854_, _01853_, rst);
  or (_01855_, _01854_, _01852_);
  or (_22653_, _01855_, _01848_);
  and (_01856_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_01857_, _00141_, _26085_);
  or (_22654_, _01857_, _01856_);
  or (_01858_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_01859_, _01858_, _25618_);
  and (_01860_, _25131_, _01826_);
  nand (_01861_, _01860_, _23729_);
  and (_01862_, _01861_, _01859_);
  nand (_01863_, _01834_, _23761_);
  and (_01864_, _01858_, _25128_);
  and (_01865_, _01864_, _01863_);
  not (_01866_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_01868_, _25127_, _01866_);
  or (_01869_, _01868_, rst);
  or (_01870_, _01869_, _01865_);
  or (_22655_, _01870_, _01862_);
  and (_01871_, _23049_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01872_, _01871_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_01873_, _23051_, _22860_);
  and (_01874_, _01873_, _23032_);
  and (_01875_, _01873_, _25071_);
  or (_01876_, _01875_, _25068_);
  or (_01877_, _01876_, _01874_);
  nor (_01878_, _25063_, _25061_);
  not (_01879_, _22998_);
  and (_01880_, _25095_, _01879_);
  nand (_01881_, _01880_, _01878_);
  or (_01882_, _01881_, _01877_);
  and (_01883_, _23052_, _23010_);
  or (_01884_, _01883_, _25060_);
  or (_01885_, _01884_, _25064_);
  and (_01886_, _25110_, _23016_);
  and (_01887_, _23018_, _22989_);
  or (_01888_, _01887_, _23034_);
  or (_01889_, _01888_, _01886_);
  or (_01891_, _01889_, _01885_);
  or (_01892_, _01891_, _01882_);
  and (_01893_, _25106_, _23052_);
  or (_01894_, _24152_, _25107_);
  or (_01895_, _01894_, _01893_);
  and (_01896_, _01873_, _24146_);
  or (_01897_, _01896_, _01895_);
  nor (_01898_, _22972_, _22808_);
  and (_01899_, _01898_, _23016_);
  and (_01900_, _01898_, _22940_);
  or (_01901_, _01900_, _01899_);
  and (_01902_, _01898_, _22997_);
  not (_01903_, _01902_);
  and (_01904_, _24164_, _22997_);
  nor (_01905_, _01904_, _24165_);
  nand (_01907_, _01905_, _01903_);
  and (_01908_, _22991_, _22949_);
  or (_01909_, _01908_, _01907_);
  or (_01910_, _01909_, _01901_);
  or (_01911_, _01910_, _01897_);
  or (_01912_, _01911_, _01892_);
  and (_01913_, _22739_, _23049_);
  and (_01914_, _01913_, _01912_);
  or (_26903_[3], _01914_, _01872_);
  and (_01915_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_01916_, _00141_, _23830_);
  or (_22656_, _01916_, _01915_);
  and (_01917_, _00096_, _23830_);
  and (_01918_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_22657_, _01918_, _01917_);
  and (_01919_, _00096_, _25886_);
  and (_01920_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_22658_, _01920_, _01919_);
  and (_01921_, _26524_, _01826_);
  nand (_01922_, _01921_, _23729_);
  or (_01923_, _01921_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01924_, _01923_, _25618_);
  and (_01925_, _01924_, _01922_);
  nand (_01926_, _01834_, _25332_);
  or (_01927_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01928_, _01927_, _25128_);
  and (_01929_, _01928_, _01926_);
  and (_01930_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_01931_, _01930_, rst);
  or (_01932_, _01931_, _01929_);
  or (_22659_, _01932_, _01925_);
  and (_01933_, _26136_, _01826_);
  nand (_01934_, _01933_, _23729_);
  or (_01935_, _01933_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01936_, _01935_, _25618_);
  and (_01937_, _01936_, _01934_);
  nand (_01938_, _01834_, _25362_);
  or (_01939_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01940_, _01939_, _25128_);
  and (_01941_, _01940_, _01938_);
  and (_01942_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_01943_, _01942_, rst);
  or (_01944_, _01943_, _01941_);
  or (_22660_, _01944_, _01937_);
  not (_01946_, _01826_);
  or (_01947_, _26564_, _01946_);
  and (_01948_, _01947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01949_, _26558_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_01950_, _01949_, _26557_);
  and (_01951_, _01950_, _01826_);
  or (_01952_, _01951_, _01948_);
  and (_01953_, _01952_, _25618_);
  nand (_01954_, _01834_, _23824_);
  or (_01956_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01957_, _01956_, _25128_);
  and (_01958_, _01957_, _01954_);
  and (_01959_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_01960_, _01959_, rst);
  or (_01961_, _01960_, _01958_);
  or (_22661_, _01961_, _01953_);
  and (_01962_, _26374_, _26204_);
  not (_01963_, _01962_);
  and (_01964_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_01965_, _01962_, _23830_);
  or (_22662_, _01965_, _01964_);
  and (_01966_, _00095_, _26224_);
  and (_01967_, _01966_, _23830_);
  not (_01968_, _01966_);
  and (_01969_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_27315_, _01969_, _01967_);
  and (_01970_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_01971_, _01962_, _25886_);
  or (_22663_, _01971_, _01970_);
  and (_01972_, _01966_, _25886_);
  and (_01973_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_22664_, _01973_, _01972_);
  and (_01975_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_01976_, _01962_, _26170_);
  or (_22665_, _01976_, _01975_);
  and (_01977_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_01978_, _01962_, _26185_);
  or (_22666_, _01978_, _01977_);
  and (_01979_, _01966_, _26242_);
  and (_01980_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_22667_, _01980_, _01979_);
  and (_01981_, _01966_, _26185_);
  and (_01982_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_22668_, _01982_, _01981_);
  and (_01984_, _01966_, _26085_);
  and (_01985_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_22669_, _01985_, _01984_);
  and (_01987_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_01988_, _01962_, _26242_);
  or (_22670_, _01988_, _01987_);
  and (_01989_, _26374_, _23848_);
  and (_01990_, _01989_, _26185_);
  not (_01991_, _01989_);
  and (_01992_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_27259_, _01992_, _01990_);
  and (_01993_, _26085_, _25939_);
  and (_01994_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_22672_, _01994_, _01993_);
  and (_01996_, _26340_, _23779_);
  not (_01997_, _01996_);
  and (_01998_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  and (_01999_, _01996_, _25886_);
  or (_22673_, _01999_, _01998_);
  and (_02001_, _26185_, _25939_);
  and (_02002_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_22674_, _02002_, _02001_);
  and (_02003_, _01604_, _26242_);
  and (_02004_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_22675_, _02004_, _02003_);
  and (_02006_, _01568_, _23830_);
  and (_02007_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_22676_, _02007_, _02006_);
  and (_02008_, _25939_, _23830_);
  and (_02009_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_22677_, _02009_, _02008_);
  and (_02010_, _23847_, _23779_);
  not (_02011_, _02010_);
  and (_02012_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  and (_02013_, _02010_, _23768_);
  or (_27073_, _02013_, _02012_);
  and (_02014_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  and (_02015_, _02010_, _25927_);
  or (_22678_, _02015_, _02014_);
  and (_02017_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  and (_02018_, _02010_, _26170_);
  or (_22679_, _02018_, _02017_);
  and (_02019_, _26258_, _23779_);
  not (_02020_, _02019_);
  and (_02021_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  and (_02023_, _02019_, _23830_);
  or (_27071_, _02023_, _02021_);
  and (_02024_, _01568_, _23768_);
  and (_02025_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_22680_, _02025_, _02024_);
  and (_02026_, _00095_, _26283_);
  and (_02028_, _02026_, _26242_);
  not (_02029_, _02026_);
  and (_02030_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_22681_, _02030_, _02028_);
  and (_02031_, _26482_, _25226_);
  nand (_02032_, _02031_, _23761_);
  or (_02034_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_02035_, _02034_, _23049_);
  and (_22682_, _02035_, _02032_);
  or (_02036_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_02037_, _02036_, _23049_);
  not (_02038_, _02031_);
  or (_02040_, _02038_, _25258_);
  and (_22683_, _02040_, _02037_);
  not (_02041_, _25279_);
  not (_02042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_02043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02044_, _25901_, _25224_);
  and (_02045_, _02044_, _01577_);
  and (_02046_, _02045_, _02043_);
  and (_02047_, _02046_, _02042_);
  and (_02049_, _02047_, _02041_);
  nor (_02050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_02051_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_02052_, _02051_, _02050_);
  not (_02053_, _02050_);
  and (_02054_, _02053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_02055_, _02054_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02056_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02058_, _02057_, _02056_);
  and (_02059_, _02058_, _02055_);
  nor (_02060_, _02059_, _02052_);
  not (_02061_, _02060_);
  and (_02062_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_02063_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02064_, _02063_, _02062_);
  nor (_02065_, _02064_, _02045_);
  and (_02066_, _02053_, _02045_);
  and (_02067_, _02066_, _25283_);
  or (_02068_, _02067_, _02065_);
  or (_02069_, _02068_, _02049_);
  and (_22684_, _02069_, _23049_);
  and (_02070_, _02066_, _25258_);
  and (_02071_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02072_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02073_, _02072_, _02071_);
  nor (_02074_, _02073_, _02045_);
  not (_02075_, _25160_);
  and (_02076_, _02047_, _02075_);
  or (_02078_, _02076_, _02074_);
  or (_02079_, _02078_, _02070_);
  and (_22685_, _02079_, _23049_);
  nor (_02081_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02082_, _02081_, _02053_);
  and (_02083_, _02082_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_02084_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_02085_, _02082_, _02084_);
  or (_02087_, _02085_, _02083_);
  and (_02088_, _26468_, _26619_);
  and (_02089_, _02088_, _26470_);
  or (_02090_, _02089_, _02087_);
  or (_02091_, _25894_, _02084_);
  nand (_02092_, _02091_, _02089_);
  or (_02093_, _02092_, _25896_);
  and (_02095_, _02093_, _02090_);
  and (_02096_, _01577_, _25902_);
  or (_02097_, _02096_, _02095_);
  not (_02098_, _02096_);
  or (_02100_, _02098_, _25258_);
  and (_02101_, _02100_, _23049_);
  and (_22686_, _02101_, _02097_);
  and (_02102_, _26273_, _23775_);
  and (_02103_, _02102_, _23830_);
  not (_02104_, _02102_);
  and (_02105_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_22687_, _02105_, _02103_);
  and (_02106_, _01568_, _25927_);
  and (_02107_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_22688_, _02107_, _02106_);
  nand (_02108_, _02066_, _25417_);
  or (_02109_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or (_02110_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and (_02111_, _02110_, _02109_);
  or (_02112_, _02111_, _02045_);
  and (_02113_, _02112_, _23049_);
  and (_22689_, _02113_, _02108_);
  and (_02114_, _02052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_02116_, _02059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_02117_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_02118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02119_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02120_, _02119_, _02118_);
  and (_02121_, _02120_, _02117_);
  nor (_02122_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02123_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02124_, _02123_, _02122_);
  and (_02125_, _02124_, _02052_);
  and (_02126_, _02125_, _02121_);
  and (_02127_, _02126_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_02128_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_02129_, _02128_, _02127_);
  and (_02130_, _02129_, _02116_);
  nor (_02131_, _02130_, _02114_);
  nor (_02132_, _02131_, _02045_);
  and (_02134_, _02047_, _25283_);
  or (_02135_, _02134_, _02132_);
  and (_22690_, _02135_, _23049_);
  not (_02136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_02137_, _02136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02138_, _02137_, _02050_);
  and (_02139_, _02138_, _02081_);
  or (_02140_, _02139_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02141_, _02140_, _02089_);
  nor (_02142_, _01448_, _23729_);
  not (_02143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02144_, _25131_, _02143_);
  nand (_02146_, _02144_, _02089_);
  or (_02147_, _02146_, _02142_);
  and (_02148_, _02147_, _02141_);
  or (_02149_, _02148_, _02096_);
  nand (_02151_, _02096_, _23761_);
  and (_02152_, _02151_, _23049_);
  and (_22691_, _02152_, _02149_);
  or (_02153_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_02154_, _02153_, _23049_);
  nand (_02155_, _02031_, _23824_);
  and (_22692_, _02155_, _02154_);
  not (_02156_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02157_, _02060_, _02156_);
  and (_02158_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_02159_, _02158_, _02157_);
  nor (_02160_, _02159_, _02045_);
  or (_02161_, _02043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02162_, _02161_, _02066_);
  or (_02163_, _02162_, _02160_);
  and (_22693_, _02163_, _23049_);
  and (_02164_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02165_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_02166_, _02165_, _02164_);
  nor (_02167_, _02166_, _02045_);
  not (_02168_, _23824_);
  and (_02169_, _02066_, _02168_);
  or (_02170_, _02169_, _02167_);
  not (_02171_, _25362_);
  and (_02172_, _02047_, _02171_);
  or (_02173_, _02172_, _02170_);
  and (_22694_, _02173_, _23049_);
  or (_02175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_02176_, _02175_, _02089_);
  nor (_02177_, _01411_, _23729_);
  nand (_02178_, _01411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_02179_, _02178_, _02089_);
  or (_02180_, _02179_, _02177_);
  and (_02181_, _02180_, _02176_);
  or (_02182_, _02181_, _02096_);
  nand (_02183_, _02096_, _25279_);
  and (_02184_, _02183_, _23049_);
  and (_22695_, _02184_, _02182_);
  or (_02185_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_02186_, _02185_, _23049_);
  nand (_02187_, _02031_, _25279_);
  and (_22696_, _02187_, _02186_);
  and (_02188_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02189_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02190_, _02189_, _02188_);
  nor (_02191_, _02190_, _02045_);
  and (_02192_, _02066_, _02041_);
  or (_02193_, _02192_, _02191_);
  and (_02195_, _02047_, _25258_);
  or (_02196_, _02195_, _02193_);
  and (_22697_, _02196_, _23049_);
  or (_02197_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_02198_, _02197_, _23049_);
  nand (_02199_, _02031_, _25362_);
  and (_22698_, _02199_, _02198_);
  and (_02200_, _02066_, _02171_);
  and (_02201_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_02202_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_02203_, _02202_, _02201_);
  nor (_02204_, _02203_, _02045_);
  not (_02205_, _25332_);
  and (_02206_, _02047_, _02205_);
  or (_02207_, _02206_, _02204_);
  or (_02208_, _02207_, _02200_);
  and (_22699_, _02208_, _23049_);
  and (_02209_, _02102_, _25886_);
  and (_02210_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_26981_, _02210_, _02209_);
  or (_02211_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_02212_, _02211_, _23049_);
  nand (_02213_, _02031_, _25160_);
  and (_22700_, _02213_, _02212_);
  and (_02214_, _02047_, _02168_);
  and (_02215_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02216_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_02217_, _02216_, _02215_);
  nor (_02218_, _02217_, _02045_);
  and (_02219_, _02066_, _02075_);
  or (_02220_, _02219_, _02218_);
  or (_02221_, _02220_, _02214_);
  and (_22701_, _02221_, _23049_);
  or (_02222_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_02223_, _02222_, _23049_);
  nand (_02224_, _02031_, _25332_);
  and (_22702_, _02224_, _02223_);
  not (_02225_, _25417_);
  and (_02226_, _02047_, _02225_);
  and (_02227_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_02228_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_02229_, _02228_, _02227_);
  nor (_02230_, _02229_, _02045_);
  and (_02231_, _02066_, _02205_);
  or (_02232_, _02231_, _02230_);
  or (_02233_, _02232_, _02226_);
  and (_22703_, _02233_, _23049_);
  not (_02234_, _02089_);
  or (_02235_, _02234_, _26564_);
  and (_02236_, _02235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02237_, _02236_, _02096_);
  and (_02238_, _26558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02239_, _02238_, _26557_);
  and (_02240_, _02239_, _02089_);
  or (_02242_, _02240_, _02237_);
  nand (_02243_, _02096_, _23824_);
  and (_02244_, _02243_, _23049_);
  and (_22704_, _02244_, _02242_);
  nand (_02246_, _02089_, _26524_);
  nor (_02247_, _02246_, _23729_);
  and (_02248_, _02246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_02249_, _02248_, _02096_);
  or (_02250_, _02249_, _02247_);
  nand (_02251_, _02096_, _25332_);
  and (_02252_, _02251_, _23049_);
  and (_22705_, _02252_, _02250_);
  and (_02253_, _02089_, _26136_);
  or (_02254_, _02253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_02255_, _02254_, _02098_);
  nand (_02256_, _02253_, _23729_);
  and (_02257_, _02256_, _02255_);
  nor (_02258_, _02098_, _25362_);
  or (_02259_, _02258_, _02257_);
  and (_22706_, _02259_, _23049_);
  nand (_02260_, _02089_, _23215_);
  and (_02261_, _02260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_02262_, _02261_, _02096_);
  and (_02263_, _25905_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_02264_, _02263_, _26475_);
  and (_02265_, _02264_, _02089_);
  or (_02267_, _02265_, _02262_);
  nand (_02268_, _02096_, _25160_);
  and (_02269_, _02268_, _23049_);
  and (_22707_, _02269_, _02267_);
  not (_02270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_02271_, _02050_, _02270_);
  and (_02272_, _02271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_02273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_02274_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _02273_);
  not (_02275_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02276_, _02275_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02277_, _02276_, _02274_);
  and (_02278_, _02277_, _02272_);
  and (_02279_, _02270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02281_, _02050_, _02143_);
  and (_02282_, _02281_, _02279_);
  and (_02283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02284_, _02283_, _02053_);
  nor (_02285_, _02284_, _02282_);
  nor (_02286_, _02285_, _02272_);
  or (_02287_, _02286_, _02278_);
  and (_02288_, _02050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02289_, _02288_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_02290_, _02289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02291_, _02290_, _02287_);
  nor (_02292_, _02289_, _02278_);
  or (_02293_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02294_, _02293_, _01634_);
  and (_02295_, _02294_, _02291_);
  or (_22708_, _02295_, _01633_);
  and (_02296_, _26204_, _23775_);
  not (_02297_, _02296_);
  and (_02298_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_02299_, _02296_, _26242_);
  or (_22709_, _02299_, _02298_);
  not (_02300_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_02301_, _02292_);
  nor (_02302_, _02301_, _02286_);
  nor (_02303_, _02302_, _02300_);
  or (_02304_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02306_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02300_);
  or (_02307_, _02306_, _02292_);
  and (_02308_, _02307_, _23049_);
  and (_22710_, _02308_, _02304_);
  and (_02309_, _01966_, _25927_);
  and (_02310_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_27314_, _02310_, _02309_);
  and (_02311_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02312_, _02284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not (_02313_, _02272_);
  nor (_02314_, _02277_, _02313_);
  and (_02315_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_02316_, _02272_, _02282_);
  or (_02317_, _02316_, _02315_);
  and (_02318_, _02317_, _02312_);
  not (_02319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_02320_, _02292_, _02319_);
  or (_02321_, _02320_, _02318_);
  nand (_02322_, _02289_, _02319_);
  and (_02323_, _02322_, _01634_);
  and (_02324_, _02323_, _02321_);
  or (_22711_, _02324_, _02311_);
  and (_02325_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  and (_02326_, _01996_, _26185_);
  or (_27085_, _02326_, _02325_);
  and (_02327_, _01966_, _23768_);
  and (_02328_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_22712_, _02328_, _02327_);
  and (_02329_, _26355_, _25914_);
  and (_02330_, _02329_, _26085_);
  not (_02331_, _02329_);
  and (_02332_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_22713_, _02332_, _02330_);
  not (_02333_, _02302_);
  or (_02334_, _02333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02335_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02336_, _02335_, _01634_);
  and (_02337_, _02336_, _02334_);
  or (_22714_, _02337_, _01638_);
  and (_02338_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_02339_, _01608_, _26242_);
  or (_22715_, _02339_, _02338_);
  and (_02340_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  and (_02341_, _02019_, _25886_);
  or (_22716_, _02341_, _02340_);
  not (_02342_, _00226_);
  nor (_02343_, _02342_, _25362_);
  and (_02344_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02346_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_02347_, _02346_, _00222_);
  and (_02348_, _02347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_02350_, _02349_, _00195_);
  and (_02351_, _02350_, _02348_);
  and (_02352_, _02346_, _00213_);
  and (_02353_, _02352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02354_, _02353_, _00209_);
  and (_02355_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02357_, _02356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_02358_, _02357_, _02355_);
  nor (_02359_, _02358_, _02351_);
  and (_02360_, _02359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_02361_, _02359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_02362_, _02361_, _02360_);
  nor (_02363_, _00226_, _00190_);
  and (_02364_, _02363_, _02362_);
  or (_02365_, _02364_, _02344_);
  or (_02366_, _02365_, _02343_);
  and (_22717_, _02366_, _23049_);
  and (_02367_, _02329_, _26185_);
  and (_02368_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_22718_, _02368_, _02367_);
  and (_02369_, _02277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02370_, _02369_, _02285_);
  or (_02371_, _02370_, _02302_);
  and (_02372_, _02371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02300_);
  nand (_02374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_02375_, _02374_, _02292_);
  or (_02376_, _02375_, _02373_);
  or (_02377_, _02376_, _02372_);
  and (_22719_, _02377_, _23049_);
  nor (_02379_, _02284_, _02272_);
  or (_02380_, _02379_, _02300_);
  or (_02382_, _02380_, _02275_);
  and (_02383_, _02272_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02384_, _02383_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_02385_, _02384_, _23049_);
  and (_22720_, _02385_, _02382_);
  nand (_02386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _23049_);
  nor (_02387_, _02386_, _02303_);
  or (_02388_, _02370_, _02301_);
  and (_02389_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_02390_, _02389_, _02388_);
  or (_22721_, _02390_, _02387_);
  and (_02391_, _02380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02395_, _02394_, _02392_);
  and (_02396_, _02395_, _02383_);
  or (_02397_, _02396_, _02391_);
  and (_22722_, _02397_, _23049_);
  and (_02398_, _02026_, _25927_);
  and (_02399_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_22723_, _02399_, _02398_);
  or (_02400_, _02055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_02401_, _02055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02402_, _02401_, rst);
  nand (_02403_, _02402_, _02400_);
  nor (_22724_, _02403_, _02045_);
  and (_02404_, _01568_, _26170_);
  and (_02405_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_22725_, _02405_, _02404_);
  and (_02406_, _02044_, _25226_);
  nand (_02407_, _02406_, _25160_);
  or (_02408_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_02409_, _02408_, _23049_);
  and (_22726_, _02409_, _02407_);
  and (_02410_, _02392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02411_, _02410_, _02273_);
  and (_02412_, _02383_, _02411_);
  and (_02413_, _02412_, rxd_i);
  not (_02414_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor (_02415_, _02412_, _02414_);
  or (_02416_, _02415_, _02413_);
  and (_22727_, _02416_, _23049_);
  or (_02417_, _02401_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_02418_, _02401_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02419_, _02418_, rst);
  nand (_02420_, _02419_, _02417_);
  nor (_22728_, _02420_, _02045_);
  nor (_02421_, _02418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_02422_, _02418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_02423_, _02422_, _02421_);
  nand (_02424_, _02423_, _23049_);
  nor (_22729_, _02424_, _02045_);
  and (_02425_, _02026_, _23768_);
  and (_02426_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_22730_, _02426_, _02425_);
  and (_02427_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_02428_, _01962_, _23768_);
  or (_27050_, _02428_, _02427_);
  or (_02429_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02430_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02300_);
  or (_02431_, _02430_, _02292_);
  and (_02432_, _02431_, _23049_);
  and (_22731_, _02432_, _02429_);
  and (_02433_, _02380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_02434_, _02410_, _02313_);
  or (_02435_, _02434_, _02433_);
  and (_02436_, _02392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02437_, _02436_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02438_, _02437_, _23049_);
  and (_22771_, _02438_, _02435_);
  and (_02440_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_22792_, _02440_, _02311_);
  and (_02441_, _23830_, _23231_);
  and (_02442_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_22795_, _02442_, _02441_);
  and (_02443_, _02026_, _23830_);
  and (_02444_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_22826_, _02444_, _02443_);
  and (_02446_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02447_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_22829_, _02447_, _02446_);
  nor (_26928_[7], _24222_, rst);
  and (_02448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02449_, _02448_, _02373_);
  and (_22834_, _02449_, _23049_);
  and (_02450_, _02026_, _25886_);
  and (_02451_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_22867_, _02451_, _02450_);
  and (_02452_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02453_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_22870_, _02453_, _02452_);
  and (_02454_, _02026_, _26170_);
  and (_02455_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_27299_, _02455_, _02454_);
  and (_02456_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and (_02457_, _02296_, _26170_);
  or (_27049_, _02457_, _02456_);
  or (_02458_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02459_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02300_);
  or (_02460_, _02459_, _02292_);
  and (_02461_, _02460_, _23049_);
  and (_22884_, _02461_, _02458_);
  or (_02462_, _02333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02463_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02464_, _02463_, _01634_);
  and (_02465_, _02464_, _02462_);
  or (_22887_, _02465_, _01636_);
  or (_02466_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02467_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02300_);
  or (_02468_, _02467_, _02292_);
  and (_02469_, _02468_, _23049_);
  and (_22890_, _02469_, _02466_);
  or (_02470_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02471_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _02300_);
  or (_02472_, _02471_, _02292_);
  and (_02473_, _02472_, _23049_);
  and (_22893_, _02473_, _02470_);
  and (_02474_, _26170_, _25939_);
  and (_02475_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_22930_, _02475_, _02474_);
  and (_02476_, _26170_, _23231_);
  and (_02477_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_22933_, _02477_, _02476_);
  and (_02478_, _01989_, _26085_);
  and (_02479_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_22941_, _02479_, _02478_);
  and (_02480_, _00095_, _23847_);
  and (_02481_, _02480_, _25927_);
  not (_02482_, _02480_);
  and (_02483_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_22955_, _02483_, _02481_);
  and (_02484_, _26193_, _25914_);
  and (_02485_, _02484_, _26242_);
  not (_02486_, _02484_);
  and (_02487_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_22978_, _02487_, _02485_);
  and (_02488_, _23849_, _23768_);
  and (_02489_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_27262_, _02489_, _02488_);
  and (_02490_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  and (_02492_, _01996_, _26170_);
  or (_23003_, _02492_, _02490_);
  and (_02493_, _02480_, _25886_);
  and (_02494_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_23014_, _02494_, _02493_);
  and (_02495_, _02480_, _26170_);
  and (_02496_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_23020_, _02496_, _02495_);
  and (_02497_, _01658_, _01654_);
  and (_02498_, _02497_, _00085_);
  and (_02499_, _02498_, _01664_);
  not (_02500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_02501_, _01654_, _02500_);
  or (_02502_, _00085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_02503_, _01664_);
  and (_02504_, _01670_, _02503_);
  and (_02505_, _02504_, _02502_);
  or (_02506_, _02505_, _02501_);
  or (_02507_, _02506_, _02499_);
  nand (_02508_, _02507_, _23049_);
  nor (_02509_, _02508_, _00071_);
  and (_23033_, _02509_, _00070_);
  and (_02510_, _01989_, _23830_);
  and (_02511_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_23060_, _02511_, _02510_);
  and (_02512_, _26374_, _25938_);
  and (_02513_, _02512_, _26170_);
  not (_02514_, _02512_);
  and (_02515_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_23107_, _02515_, _02513_);
  and (_02517_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_02518_, _02296_, _23830_);
  or (_23128_, _02518_, _02517_);
  and (_02519_, _26202_, _23230_);
  and (_02520_, _02519_, _23768_);
  not (_02521_, _02519_);
  and (_02522_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_23135_, _02522_, _02520_);
  and (_02523_, _02480_, _26185_);
  and (_02524_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_23141_, _02524_, _02523_);
  and (_02525_, _02480_, _26085_);
  and (_02526_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_27289_, _02526_, _02525_);
  and (_02527_, _02480_, _23830_);
  and (_02528_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_23164_, _02528_, _02527_);
  nor (_02529_, _02342_, _25279_);
  and (_02530_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_02531_, _00221_, _00213_);
  and (_02532_, _02531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_02533_, _02532_, _00209_);
  and (_02534_, _02533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_02535_, _02533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_02536_, _02535_, _02534_);
  and (_02537_, _02536_, _00195_);
  and (_02538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02539_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_02540_, _02539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_02541_, _02352_, _00209_);
  and (_02542_, _02541_, _02356_);
  and (_02543_, _02542_, _02540_);
  or (_02544_, _02543_, _02538_);
  or (_02545_, _02544_, _02537_);
  and (_02546_, _02545_, _02363_);
  or (_02547_, _02546_, _02530_);
  or (_02548_, _02547_, _02529_);
  and (_23172_, _02548_, _23049_);
  nand (_02549_, _00190_, _23824_);
  and (_02550_, _00193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_02551_, _02550_, _00209_);
  and (_02552_, _02551_, _02531_);
  not (_02553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_02554_, _01617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_02555_, _02554_, _02553_);
  nor (_02556_, _01618_, _00214_);
  and (_02557_, _02556_, _02555_);
  nor (_02558_, _02557_, _02552_);
  nor (_02559_, _02558_, _00226_);
  nor (_02560_, _01625_, _02553_);
  or (_02561_, _02560_, _02559_);
  or (_02562_, _02561_, _00190_);
  and (_02563_, _02562_, _23049_);
  and (_23188_, _02563_, _02549_);
  and (_02564_, _26213_, _26204_);
  not (_02565_, _02564_);
  and (_02566_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_02567_, _02564_, _26185_);
  or (_23206_, _02567_, _02566_);
  and (_02568_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_02569_, _02564_, _26242_);
  or (_23228_, _02569_, _02568_);
  and (_02570_, _00095_, _26258_);
  and (_02571_, _02570_, _23830_);
  not (_02572_, _02570_);
  and (_02573_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_23241_, _02573_, _02571_);
  and (_02574_, _02570_, _25886_);
  and (_02575_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_23254_, _02575_, _02574_);
  and (_02576_, _26224_, _23779_);
  not (_02577_, _02576_);
  and (_02578_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  and (_02579_, _02576_, _25886_);
  or (_23301_, _02579_, _02578_);
  and (_02580_, _25939_, _25927_);
  and (_02581_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_23310_, _02581_, _02580_);
  and (_02582_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_02583_, _02296_, _23768_);
  or (_23314_, _02583_, _02582_);
  and (_02584_, _02570_, _26242_);
  and (_02585_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_23330_, _02585_, _02584_);
  and (_02586_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  and (_02587_, _26214_, _25886_);
  or (_27065_, _02587_, _02586_);
  and (_02588_, _02570_, _26185_);
  and (_02589_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_27268_, _02589_, _02588_);
  and (_02590_, _00095_, _26374_);
  and (_02591_, _02590_, _26242_);
  not (_02592_, _02590_);
  and (_02593_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_23396_, _02593_, _02591_);
  and (_02594_, _02590_, _26185_);
  and (_02595_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_23399_, _02595_, _02594_);
  and (_02596_, _02519_, _23830_);
  and (_02598_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_23409_, _02598_, _02596_);
  and (_02599_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_02600_, _02564_, _25927_);
  or (_23413_, _02600_, _02599_);
  and (_02601_, _02570_, _25927_);
  and (_02602_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_23431_, _02602_, _02601_);
  and (_02603_, _02570_, _23768_);
  and (_02604_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_23434_, _02604_, _02603_);
  and (_02605_, _02484_, _26185_);
  and (_02606_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_23442_, _02606_, _02605_);
  and (_02607_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_02608_, _02564_, _25886_);
  or (_27048_, _02608_, _02607_);
  and (_02609_, _00095_, _23775_);
  and (_02610_, _02609_, _26242_);
  not (_02611_, _02609_);
  and (_02612_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_23477_, _02612_, _02610_);
  and (_02613_, _02590_, _23768_);
  and (_02614_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_27251_, _02614_, _02613_);
  and (_02615_, _26204_, _26190_);
  not (_02616_, _02615_);
  and (_02617_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_02618_, _02615_, _26185_);
  or (_27046_, _02618_, _02617_);
  and (_02619_, _02590_, _26170_);
  and (_02620_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_23508_, _02620_, _02619_);
  and (_02622_, _02590_, _25927_);
  and (_02623_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_23537_, _02623_, _02622_);
  nand (_02624_, _02406_, _23824_);
  or (_02625_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_02626_, _02625_, _23049_);
  and (_23593_, _02626_, _02624_);
  and (_02628_, _00226_, _25258_);
  and (_02629_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_02630_, _02347_, _00192_);
  or (_02631_, _02542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_02632_, _02631_, _02630_);
  and (_02633_, _02632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02634_, _02352_, _02356_);
  and (_02635_, _02346_, _00195_);
  and (_02636_, _02635_, _02531_);
  or (_02637_, _02636_, _02634_);
  not (_02638_, _00209_);
  nor (_02639_, _02638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02640_, _02639_, _02637_);
  or (_02641_, _02640_, _02633_);
  and (_02642_, _02641_, _02363_);
  or (_02643_, _02642_, _02629_);
  or (_02644_, _02643_, _02628_);
  and (_23596_, _02644_, _23049_);
  nand (_02645_, _02406_, _25362_);
  or (_02646_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02647_, _02646_, _23049_);
  and (_23638_, _02647_, _02645_);
  nor (_02648_, _02342_, _25160_);
  and (_02649_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_02650_, _02534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_02651_, _02650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_02652_, _02650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_02653_, _02652_, _02651_);
  and (_02654_, _02653_, _00195_);
  or (_02655_, _02354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not (_02656_, _02356_);
  nor (_02657_, _02355_, _02656_);
  and (_02658_, _02657_, _02655_);
  and (_02659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_02660_, _02659_, _02658_);
  or (_02661_, _02660_, _02654_);
  and (_02662_, _02661_, _02363_);
  or (_02663_, _02662_, _02649_);
  or (_02664_, _02663_, _02648_);
  and (_23641_, _02664_, _23049_);
  nand (_02665_, _02406_, _25332_);
  or (_02666_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_02667_, _02666_, _23049_);
  and (_23658_, _02667_, _02665_);
  and (_02668_, _22992_, _22973_);
  and (_02669_, _02668_, _22862_);
  nor (_02670_, _02669_, _25090_);
  and (_02671_, _02670_, _25089_);
  nor (_02672_, _25079_, _25068_);
  and (_02674_, _02672_, _25073_);
  and (_02675_, _25584_, _22862_);
  nor (_02676_, _24148_, _02675_);
  and (_02677_, _02676_, _25065_);
  and (_02678_, _02677_, _02674_);
  and (_02679_, _02678_, _02671_);
  nor (_02680_, _02679_, _23061_);
  nor (_02681_, _02676_, _24161_);
  nor (_02682_, _02681_, _02680_);
  nor (_26944_, _02682_, rst);
  and (_02683_, _25186_, _25225_);
  and (_02684_, _02683_, _00255_);
  and (_02685_, _02684_, _25187_);
  nand (_02686_, _02685_, _25417_);
  or (_02687_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_02688_, _02687_, _23049_);
  and (_26906_[7], _02688_, _02686_);
  and (_02689_, _02683_, _01843_);
  not (_02690_, _02689_);
  nor (_02691_, _02690_, _25417_);
  not (_02692_, _25187_);
  and (_02693_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_02694_, _02693_, _02692_);
  or (_02695_, _02694_, _02691_);
  or (_02696_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_02698_, _02696_, _23049_);
  and (_26907_[7], _02698_, _02695_);
  and (_02699_, _25131_, _23154_);
  and (_02700_, _02683_, _02699_);
  and (_02701_, _02700_, _25187_);
  nand (_02702_, _02701_, _25417_);
  or (_02703_, _02701_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_02704_, _02703_, _23049_);
  and (_26908_[7], _02704_, _02702_);
  and (_02705_, _25224_, _23154_);
  and (_02706_, _02683_, _02705_);
  and (_02707_, _02706_, _25187_);
  not (_02708_, _02707_);
  nor (_02709_, _02708_, _25417_);
  and (_02710_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_02711_, _02710_, _02709_);
  and (_26909_[7], _02711_, _23049_);
  and (_02712_, _25186_, _25134_);
  and (_02713_, _02712_, _00255_);
  and (_02714_, _02713_, _25187_);
  and (_02715_, _02714_, _02225_);
  nor (_02716_, _02689_, _02684_);
  nor (_02717_, _02706_, _02700_);
  nand (_02718_, _02717_, _02716_);
  not (_02719_, _02713_);
  and (_02720_, _02719_, _02717_);
  and (_02721_, _02720_, _02716_);
  or (_02722_, _02721_, _02692_);
  or (_02723_, _02722_, _02718_);
  and (_02724_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_02725_, _02724_, _02715_);
  and (_26910_[7], _02725_, _23049_);
  nand (_02726_, _02716_, _25187_);
  not (_02727_, _02700_);
  nand (_02728_, _02727_, _02716_);
  and (_02729_, _02712_, _01843_);
  or (_02730_, _02729_, _02713_);
  or (_02731_, _02730_, _02706_);
  nor (_02732_, _02731_, _02728_);
  or (_02733_, _02732_, _02726_);
  and (_02734_, _02733_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_02735_, _02729_, _02225_);
  not (_02736_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_02738_, _02720_, _02736_);
  or (_02739_, _02738_, _02735_);
  and (_02740_, _02739_, _25187_);
  or (_02741_, _02740_, _02734_);
  and (_26911_[7], _02741_, _23049_);
  and (_02742_, _02712_, _02699_);
  and (_02743_, _02742_, _25187_);
  not (_02744_, _02743_);
  nor (_02745_, _02744_, _25417_);
  and (_02746_, _02744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_02747_, _02746_, _02745_);
  and (_26912_[7], _02747_, _23049_);
  and (_02748_, _02712_, _02705_);
  and (_02749_, _02748_, _25187_);
  not (_02750_, _02749_);
  nor (_02751_, _02750_, _25417_);
  or (_02752_, _02742_, _02730_);
  nor (_02753_, _02752_, _02718_);
  not (_02754_, _02748_);
  and (_02755_, _02754_, _02753_);
  or (_02756_, _02718_, _02692_);
  and (_02757_, _02752_, _25187_);
  or (_02759_, _02757_, _02756_);
  or (_02760_, _02759_, _02755_);
  and (_02761_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_02762_, _02761_, _02751_);
  and (_26913_[7], _02762_, _23049_);
  and (_02763_, _02609_, _23768_);
  and (_02764_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_23778_, _02764_, _02763_);
  and (_02766_, _02609_, _26170_);
  and (_02767_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_23785_, _02767_, _02766_);
  and (_02768_, _02609_, _25927_);
  and (_02769_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_27243_, _02769_, _02768_);
  and (_02770_, _02609_, _26085_);
  and (_02771_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_23881_, _02771_, _02770_);
  and (_02772_, _02609_, _23830_);
  and (_02773_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_27244_, _02773_, _02772_);
  and (_02774_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_02775_, _02615_, _26170_);
  or (_23917_, _02775_, _02774_);
  and (_02776_, _02609_, _25886_);
  and (_02777_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_23924_, _02777_, _02776_);
  and (_02778_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_02779_, _02615_, _25927_);
  or (_23927_, _02779_, _02778_);
  and (_02780_, _00095_, _26213_);
  and (_02781_, _02780_, _23830_);
  not (_02782_, _02780_);
  and (_02783_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_23981_, _02783_, _02781_);
  and (_02784_, _02780_, _25886_);
  and (_02785_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_23984_, _02785_, _02784_);
  and (_02786_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_02787_, _02615_, _25886_);
  or (_24028_, _02787_, _02786_);
  and (_02788_, _02780_, _26242_);
  and (_02789_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_24082_, _02789_, _02788_);
  and (_02790_, _02780_, _26185_);
  and (_02791_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_24090_, _02791_, _02790_);
  and (_02792_, _26204_, _25914_);
  not (_02793_, _02792_);
  and (_02794_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_02795_, _02792_, _23830_);
  or (_27044_, _02795_, _02794_);
  and (_02796_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and (_02797_, _02792_, _26085_);
  or (_27045_, _02797_, _02796_);
  and (_02798_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_02799_, _02792_, _25886_);
  or (_24111_, _02799_, _02798_);
  and (_02800_, _00095_, _26190_);
  and (_02801_, _02800_, _26242_);
  not (_02802_, _02800_);
  and (_02803_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_24147_, _02803_, _02801_);
  and (_02804_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_02805_, _02792_, _26242_);
  or (_24181_, _02805_, _02804_);
  and (_02806_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_02807_, _02792_, _26185_);
  or (_24187_, _02807_, _02806_);
  and (_02808_, _02780_, _25927_);
  and (_02809_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_24190_, _02809_, _02808_);
  and (_02811_, _02780_, _23768_);
  and (_02812_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_24197_, _02812_, _02811_);
  and (_02813_, _02800_, _25927_);
  and (_02814_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_24215_, _02814_, _02813_);
  and (_02815_, _02800_, _23768_);
  and (_02816_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_24229_, _02816_, _02815_);
  and (_02817_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_02818_, _02792_, _25927_);
  or (_24309_, _02818_, _02817_);
  and (_02819_, _02800_, _23830_);
  and (_02820_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_24312_, _02820_, _02819_);
  and (_02821_, _02800_, _25886_);
  and (_02822_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_27117_, _02822_, _02821_);
  nand (_02823_, _02685_, _25362_);
  or (_02824_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_26947_, _02824_, _02823_);
  and (_02825_, _23777_, _23223_);
  and (_02826_, _02825_, _26202_);
  and (_02827_, _02826_, _23830_);
  not (_02828_, _02826_);
  and (_02829_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_24368_, _02829_, _02827_);
  nand (_02831_, _02685_, _23824_);
  or (_02832_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_24371_, _02832_, _02831_);
  and (_02833_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_02834_, _23780_, _23768_);
  or (_24459_, _02834_, _02833_);
  or (_02835_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_24463_, _02835_, _02686_);
  and (_02836_, _02826_, _26185_);
  and (_02837_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_24472_, _02837_, _02836_);
  and (_02838_, _02826_, _26242_);
  and (_02839_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_24488_, _02839_, _02838_);
  and (_02840_, _02685_, _25283_);
  not (_02841_, _02685_);
  and (_02842_, _02841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_24501_, _02842_, _02840_);
  and (_02843_, _02826_, _23768_);
  and (_02844_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_24511_, _02844_, _02843_);
  nand (_02845_, _02685_, _25279_);
  or (_02846_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_24563_, _02846_, _02845_);
  and (_02847_, _02826_, _25927_);
  and (_02848_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_24602_, _02848_, _02847_);
  and (_02849_, _02825_, _23220_);
  and (_02850_, _02849_, _23830_);
  not (_02851_, _02849_);
  and (_02852_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or (_24648_, _02852_, _02850_);
  and (_02853_, _02849_, _26185_);
  and (_02854_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or (_27042_, _02854_, _02853_);
  nor (_02855_, _02342_, _25417_);
  and (_02856_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02857_, _02349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02858_, _02857_, _00209_);
  and (_02859_, _02532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_02860_, _02859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02861_, _02860_, _02858_);
  and (_02862_, _02861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_02863_, _02862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02864_, _02862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02865_, _02864_, _02863_);
  and (_02866_, _02865_, _00195_);
  and (_02867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02868_, _02858_, _02353_);
  and (_02869_, _02868_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_02870_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_02871_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02872_, _02871_, _02870_);
  and (_02873_, _02872_, _02356_);
  or (_02874_, _02873_, _02867_);
  or (_02875_, _02874_, _02866_);
  and (_02876_, _02875_, _02363_);
  or (_02877_, _02876_, _02856_);
  or (_02878_, _02877_, _02855_);
  and (_24680_, _02878_, _23049_);
  and (_02879_, _26421_, _26204_);
  not (_02880_, _02879_);
  and (_02881_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and (_02882_, _02879_, _26242_);
  or (_24699_, _02882_, _02881_);
  and (_02883_, _26242_, _26073_);
  and (_02884_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_24702_, _02884_, _02883_);
  and (_02885_, _02841_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  or (_02886_, _02885_, _02840_);
  and (_26906_[0], _02886_, _23049_);
  or (_02887_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_02888_, _02887_, _23049_);
  and (_26906_[1], _02888_, _02845_);
  or (_02890_, _02841_, _25258_);
  or (_02891_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_02892_, _02891_, _23049_);
  and (_26906_[2], _02892_, _02890_);
  nand (_02893_, _02685_, _25160_);
  or (_02894_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_02895_, _02894_, _23049_);
  and (_26906_[3], _02895_, _02893_);
  or (_02896_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02897_, _02896_, _23049_);
  and (_26906_[4], _02897_, _02831_);
  or (_02898_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_02899_, _02898_, _23049_);
  and (_26906_[5], _02899_, _02823_);
  nand (_02900_, _02685_, _25332_);
  or (_02901_, _02685_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02902_, _02901_, _23049_);
  and (_26906_[6], _02902_, _02900_);
  and (_02903_, _02689_, _25187_);
  or (_02904_, _02903_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nand (_02905_, _02903_, _23761_);
  and (_02906_, _02905_, _23049_);
  and (_26907_[0], _02906_, _02904_);
  nor (_02907_, _02690_, _25279_);
  and (_02908_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_02909_, _02908_, _02692_);
  or (_02910_, _02909_, _02907_);
  or (_02911_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_02912_, _02911_, _23049_);
  and (_26907_[1], _02912_, _02910_);
  and (_02914_, _02689_, _25258_);
  and (_02915_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_02916_, _02915_, _02692_);
  or (_02917_, _02916_, _02914_);
  or (_02918_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_02919_, _02918_, _23049_);
  and (_26907_[2], _02919_, _02917_);
  nor (_02920_, _02690_, _25160_);
  and (_02921_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_02922_, _02921_, _02692_);
  or (_02923_, _02922_, _02920_);
  or (_02925_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_02926_, _02925_, _23049_);
  and (_26907_[3], _02926_, _02923_);
  nor (_02927_, _02690_, _23824_);
  and (_02928_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_02929_, _02928_, _02692_);
  or (_02930_, _02929_, _02927_);
  or (_02931_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_02932_, _02931_, _23049_);
  and (_26907_[4], _02932_, _02930_);
  nor (_02933_, _02690_, _25362_);
  and (_02934_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_02935_, _02934_, _02692_);
  or (_02936_, _02935_, _02933_);
  or (_02937_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_02938_, _02937_, _23049_);
  and (_26907_[5], _02938_, _02936_);
  nor (_02940_, _02690_, _25332_);
  and (_02941_, _02690_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_02942_, _02941_, _02692_);
  or (_02943_, _02942_, _02940_);
  or (_02944_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_02945_, _02944_, _23049_);
  and (_26907_[6], _02945_, _02943_);
  nand (_02946_, _02701_, _23761_);
  or (_02947_, _02701_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02948_, _02947_, _02946_);
  and (_26908_[0], _02948_, _23049_);
  not (_02949_, _02701_);
  nor (_02950_, _02949_, _25279_);
  and (_02951_, _02949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_02952_, _02951_, _02950_);
  and (_26908_[1], _02952_, _23049_);
  and (_02953_, _02701_, _25258_);
  and (_02954_, _02949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_02955_, _02954_, _02953_);
  and (_26908_[2], _02955_, _23049_);
  nor (_02956_, _02949_, _25160_);
  and (_02957_, _02949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_02958_, _02957_, _02956_);
  and (_26908_[3], _02958_, _23049_);
  nor (_02959_, _02949_, _23824_);
  and (_02960_, _02949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_02961_, _02960_, _02959_);
  and (_26908_[4], _02961_, _23049_);
  nand (_02962_, _02701_, _25362_);
  or (_02963_, _02701_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_02964_, _02963_, _23049_);
  and (_26908_[5], _02964_, _02962_);
  nor (_02965_, _02949_, _25332_);
  and (_02966_, _02949_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_02967_, _02966_, _02965_);
  and (_26908_[6], _02967_, _23049_);
  and (_02968_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_02969_, _02707_, _25283_);
  or (_02970_, _02969_, _02968_);
  and (_26909_[0], _02970_, _23049_);
  nor (_02971_, _02708_, _25279_);
  and (_02972_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_02973_, _02972_, _02971_);
  and (_26909_[1], _02973_, _23049_);
  and (_02974_, _02707_, _25258_);
  and (_02975_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_02976_, _02975_, _02974_);
  and (_26909_[2], _02976_, _23049_);
  nor (_02977_, _02708_, _25160_);
  and (_02978_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_02979_, _02978_, _02977_);
  and (_26909_[3], _02979_, _23049_);
  and (_02980_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_02982_, _02708_, _23824_);
  or (_02983_, _02982_, _02980_);
  and (_26909_[4], _02983_, _23049_);
  nor (_02984_, _02708_, _25362_);
  and (_02985_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_02986_, _02985_, _02984_);
  and (_26909_[5], _02986_, _23049_);
  nor (_02987_, _02708_, _25332_);
  and (_02988_, _02708_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_02989_, _02988_, _02987_);
  and (_26909_[6], _02989_, _23049_);
  and (_02991_, _02713_, _25283_);
  and (_02992_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_02993_, _02992_, _02991_);
  or (_02994_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_02995_, _02994_, _23049_);
  and (_26910_[0], _02995_, _02993_);
  or (_02996_, _02722_, _02684_);
  and (_02997_, _02996_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_02998_, _02714_, _02041_);
  nand (_02999_, _02717_, _02690_);
  and (_03000_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_03001_, _03000_, _02999_);
  or (_03002_, _03001_, _02998_);
  or (_03003_, _03002_, _02997_);
  and (_26910_[1], _03003_, _23049_);
  and (_03004_, _02714_, _25258_);
  and (_03005_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_03006_, _03005_, _03004_);
  and (_26910_[2], _03006_, _23049_);
  and (_03007_, _02714_, _02075_);
  and (_03008_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_03009_, _03008_, _03007_);
  and (_26910_[3], _03009_, _23049_);
  and (_03010_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03011_, _02714_, _02168_);
  or (_03012_, _03011_, _03010_);
  and (_26910_[4], _03012_, _23049_);
  and (_03013_, _02714_, _02171_);
  and (_03014_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_03015_, _03014_, _03013_);
  and (_26910_[5], _03015_, _23049_);
  and (_03016_, _02714_, _02205_);
  and (_03017_, _02723_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  or (_03018_, _03017_, _03016_);
  and (_26910_[6], _03018_, _23049_);
  nor (_03020_, _02720_, _02692_);
  or (_03021_, _03020_, _02733_);
  and (_03022_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_03023_, _02692_, _23761_);
  and (_03024_, _03023_, _02729_);
  or (_03025_, _03024_, _03022_);
  and (_26911_[0], _03025_, _23049_);
  and (_03026_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_03027_, _02729_, _25187_);
  and (_03028_, _03027_, _02041_);
  or (_03029_, _03028_, _03026_);
  and (_26911_[1], _03029_, _23049_);
  and (_03031_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03032_, _03027_, _25258_);
  or (_03033_, _03032_, _03031_);
  and (_26911_[2], _03033_, _23049_);
  and (_03034_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_03035_, _03027_, _02075_);
  or (_03036_, _03035_, _03034_);
  and (_26911_[3], _03036_, _23049_);
  and (_03037_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_03038_, _03027_, _02168_);
  or (_03039_, _03038_, _03037_);
  and (_26911_[4], _03039_, _23049_);
  and (_03040_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03041_, _03027_, _02171_);
  or (_03042_, _03041_, _03040_);
  and (_26911_[5], _03042_, _23049_);
  and (_03043_, _03021_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_03044_, _03027_, _02205_);
  or (_03045_, _03044_, _03043_);
  and (_26911_[6], _03045_, _23049_);
  or (_03046_, _02753_, _02692_);
  and (_03047_, _03046_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand (_03048_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_03049_, _03048_, _02732_);
  and (_03050_, _02743_, _25283_);
  or (_03051_, _03050_, _03049_);
  or (_03052_, _03051_, _03047_);
  and (_26912_[0], _03052_, _23049_);
  or (_03053_, _03046_, _02728_);
  and (_03054_, _03053_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_03055_, _02744_, _25279_);
  and (_03056_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_03057_, _03056_, _02731_);
  or (_03058_, _03057_, _03055_);
  or (_03059_, _03058_, _03054_);
  and (_26912_[1], _03059_, _23049_);
  and (_03060_, _02744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_03062_, _02743_, _25258_);
  or (_03063_, _03062_, _03060_);
  and (_26912_[2], _03063_, _23049_);
  and (_03065_, _03053_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_03066_, _02744_, _25160_);
  and (_03067_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_03068_, _03067_, _02731_);
  or (_03069_, _03068_, _03066_);
  or (_03071_, _03069_, _03065_);
  and (_26912_[3], _03071_, _23049_);
  and (_03073_, _03046_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand (_03074_, _25187_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_03075_, _03074_, _02732_);
  nor (_03077_, _02744_, _23824_);
  or (_03078_, _03077_, _03075_);
  or (_03079_, _03078_, _03073_);
  and (_26912_[4], _03079_, _23049_);
  and (_03080_, _02744_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_03082_, _02744_, _25362_);
  or (_03084_, _03082_, _03080_);
  and (_26912_[5], _03084_, _23049_);
  nor (_03085_, _02744_, _25332_);
  and (_03086_, _02731_, _25187_);
  or (_03087_, _03086_, _03053_);
  and (_03088_, _03087_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_03089_, _03088_, _03085_);
  and (_26912_[6], _03089_, _23049_);
  and (_03090_, _02749_, _25283_);
  and (_03091_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_03092_, _03091_, _03090_);
  and (_26913_[0], _03092_, _23049_);
  nor (_03093_, _02750_, _25279_);
  and (_03094_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or (_03095_, _03094_, _03093_);
  and (_26913_[1], _03095_, _23049_);
  and (_03096_, _02749_, _25258_);
  and (_03097_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_03098_, _03097_, _03096_);
  and (_26913_[2], _03098_, _23049_);
  nor (_03099_, _02750_, _25160_);
  and (_03100_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_03101_, _03100_, _03099_);
  and (_26913_[3], _03101_, _23049_);
  nor (_03102_, _02750_, _23824_);
  and (_03103_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_03104_, _03103_, _03102_);
  and (_26913_[4], _03104_, _23049_);
  nor (_03105_, _02750_, _25362_);
  and (_03106_, _02760_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or (_03107_, _03106_, _03105_);
  and (_26913_[5], _03107_, _23049_);
  and (_03108_, _02750_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_03109_, _02750_, _25332_);
  or (_03110_, _03109_, _03108_);
  and (_26913_[6], _03110_, _23049_);
  and (_03113_, _26176_, _23768_);
  and (_03114_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_25016_, _03114_, _03113_);
  and (_03115_, _25932_, _23848_);
  and (_03116_, _03115_, _26185_);
  not (_03117_, _03115_);
  and (_03118_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_25067_, _03118_, _03116_);
  and (_03120_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_03121_, _02879_, _26185_);
  or (_25229_, _03121_, _03120_);
  nor (_03122_, _02342_, _25332_);
  and (_03123_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_03124_, _02857_, _02354_);
  nor (_03125_, _00221_, _00192_);
  nor (_03126_, _03125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_03127_, _03126_, _03124_);
  nand (_03129_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_03130_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_03131_, _03130_, _03129_);
  and (_03132_, _03131_, _02363_);
  or (_03133_, _03132_, _03123_);
  or (_03135_, _03133_, _03122_);
  and (_25315_, _03135_, _23049_);
  and (_03136_, _02329_, _26242_);
  and (_03137_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_25321_, _03137_, _03136_);
  and (_03138_, _26351_, _25927_);
  and (_03139_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_25327_, _03139_, _03138_);
  and (_03140_, _26176_, _25927_);
  and (_03142_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_26970_, _03142_, _03140_);
  not (_03144_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03145_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_03146_, _03145_, _03144_);
  and (_03147_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _23049_);
  and (_27327_, _03147_, _03146_);
  nor (_03148_, _03146_, rst);
  nand (_03149_, _03145_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03151_, _03145_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03152_, _03151_, _03149_);
  and (_27328_[3], _03152_, _03148_);
  not (_03153_, _25525_);
  nor (_03154_, _03153_, _25402_);
  not (_03155_, _25485_);
  and (_03156_, _03155_, _25445_);
  and (_03157_, _03156_, _25301_);
  and (_03158_, _03157_, _03154_);
  not (_03159_, _25613_);
  nand (_03161_, _00713_, _03159_);
  and (_03162_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_03163_, _26130_, _23351_);
  nor (_03164_, _03163_, _26557_);
  and (_03165_, _25620_, _25614_);
  not (_03166_, _03165_);
  nor (_03167_, _03166_, _03164_);
  nor (_03168_, _03167_, _03162_);
  and (_03169_, _03168_, _25607_);
  nand (_03170_, _03169_, _03161_);
  nor (_03172_, _01109_, _25607_);
  not (_03173_, _03172_);
  and (_03174_, _03173_, _03170_);
  nand (_03175_, _00773_, _03159_);
  and (_03176_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_03178_, _01686_, _23729_);
  nor (_03180_, _26136_, _23319_);
  nor (_03181_, _03180_, _03178_);
  nor (_03182_, _03181_, _03166_);
  nor (_03183_, _03182_, _03176_);
  and (_03184_, _03183_, _25607_);
  and (_03185_, _03184_, _03175_);
  and (_03186_, _01160_, _25606_);
  nor (_03187_, _03186_, _03185_);
  nand (_03188_, _03187_, _03174_);
  or (_03189_, _03187_, _03174_);
  nand (_03190_, _03189_, _03188_);
  nand (_03191_, _00836_, _03159_);
  and (_03192_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_03193_, _26524_, _23573_);
  nor (_03195_, _03193_, _00244_);
  nor (_03196_, _03195_, _03166_);
  nor (_03197_, _03196_, _03192_);
  and (_03198_, _03197_, _25607_);
  nand (_03199_, _03198_, _03191_);
  or (_03200_, _01204_, _25607_);
  and (_03201_, _03200_, _03199_);
  nand (_03202_, _03159_, _25053_);
  and (_03203_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_03204_, _25536_);
  nor (_03206_, _03204_, _23729_);
  nor (_03207_, _25536_, _23284_);
  nor (_03208_, _03207_, _03206_);
  nor (_03209_, _03208_, _03166_);
  nor (_03210_, _03209_, _03203_);
  and (_03211_, _03210_, _25607_);
  nand (_03213_, _03211_, _03202_);
  or (_03214_, _25846_, _25607_);
  and (_03216_, _03214_, _03213_);
  or (_03217_, _03216_, _03201_);
  nand (_03218_, _03216_, _03201_);
  and (_03219_, _03218_, _03217_);
  nand (_03220_, _03219_, _03190_);
  or (_03221_, _03219_, _03190_);
  nand (_03222_, _03221_, _03220_);
  and (_03223_, _00500_, _03159_);
  and (_03225_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_03226_, _25131_, _23480_);
  or (_03227_, _03226_, _02142_);
  and (_03229_, _03227_, _03165_);
  or (_03230_, _03229_, _03225_);
  or (_03231_, _03230_, _25606_);
  or (_03232_, _03231_, _03223_);
  or (_03233_, _00910_, _25607_);
  and (_03234_, _03233_, _03232_);
  and (_03235_, _00557_, _03159_);
  and (_03237_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_03238_, _25224_, _23451_);
  or (_03239_, _03238_, _02177_);
  and (_03240_, _03239_, _03165_);
  or (_03241_, _03240_, _03237_);
  or (_03242_, _03241_, _25606_);
  or (_03243_, _03242_, _03235_);
  or (_03245_, _00959_, _25607_);
  and (_03246_, _03245_, _03243_);
  or (_03247_, _03246_, _03234_);
  nand (_03248_, _03246_, _03234_);
  nand (_03249_, _03248_, _03247_);
  or (_03250_, _00608_, _25613_);
  and (_03251_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_03252_, _25894_, _23416_);
  nor (_03253_, _03252_, _25896_);
  nor (_03255_, _03253_, _03166_);
  nor (_03256_, _03255_, _03251_);
  and (_03257_, _03256_, _25607_);
  and (_03258_, _03257_, _03250_);
  and (_03259_, _01012_, _25606_);
  or (_03260_, _03259_, _03258_);
  and (_03261_, _00659_, _03159_);
  and (_03262_, _25622_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_03263_, _26473_, _23381_);
  or (_03264_, _03263_, _26475_);
  and (_03265_, _03264_, _03165_);
  or (_03266_, _03265_, _03262_);
  or (_03267_, _03266_, _25606_);
  or (_03268_, _03267_, _03261_);
  or (_03269_, _01059_, _25607_);
  and (_03270_, _03269_, _03268_);
  or (_03272_, _03270_, _03260_);
  nand (_03273_, _03270_, _03260_);
  and (_03275_, _03273_, _03272_);
  nand (_03277_, _03275_, _03249_);
  or (_03278_, _03275_, _03249_);
  nand (_03279_, _03278_, _03277_);
  nand (_03281_, _03279_, _03222_);
  or (_03282_, _03279_, _03222_);
  and (_03283_, _03282_, _03281_);
  nand (_03284_, _03283_, _25707_);
  and (_03286_, _25748_, _25671_);
  or (_03287_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03288_, _03287_, _03286_);
  and (_03289_, _03288_, _03284_);
  not (_03290_, _25707_);
  not (_03291_, _25671_);
  and (_03292_, _25748_, _03291_);
  and (_03293_, _03292_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_03294_, _25748_, _25671_);
  and (_03296_, _03294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03297_, _03296_, _03293_);
  and (_03299_, _03297_, _03290_);
  nor (_03300_, _25748_, _03291_);
  nor (_03301_, _25707_, _00644_);
  and (_03302_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03304_, _03302_, _03301_);
  and (_03305_, _03304_, _03300_);
  and (_03306_, _03292_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03307_, _03294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03308_, _03307_, _03306_);
  and (_03309_, _03308_, _25707_);
  or (_03310_, _03309_, _03305_);
  or (_03311_, _03310_, _03299_);
  or (_03312_, _03311_, _03289_);
  and (_03313_, _03312_, _03158_);
  and (_03314_, _25757_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_03315_, _25301_);
  and (_03316_, _25485_, _25445_);
  and (_03317_, _03316_, _03315_);
  and (_03318_, _25525_, _25402_);
  and (_03319_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03320_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03322_, _03320_, _03319_);
  and (_03323_, _03322_, _03300_);
  nor (_03324_, _25707_, _01651_);
  and (_03325_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03326_, _03325_, _03324_);
  and (_03327_, _03326_, _03286_);
  or (_03328_, _03327_, _03323_);
  and (_03329_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_03330_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03331_, _03330_, _03329_);
  and (_03332_, _03331_, _03292_);
  and (_03333_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03334_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03335_, _03334_, _03333_);
  and (_03336_, _03335_, _03294_);
  or (_03337_, _03336_, _03332_);
  or (_03338_, _03337_, _03328_);
  and (_03339_, _03338_, _03318_);
  and (_03340_, _03153_, _25402_);
  and (_03341_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03342_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03343_, _03342_, _03341_);
  and (_03345_, _03343_, _03300_);
  nor (_03346_, _25707_, _26666_);
  and (_03347_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03349_, _03347_, _03346_);
  and (_03351_, _03349_, _03286_);
  or (_03353_, _03351_, _03345_);
  and (_03354_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03355_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_03356_, _03355_, _03354_);
  and (_03357_, _03356_, _03294_);
  nor (_03358_, _25707_, _26670_);
  and (_03359_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03360_, _03359_, _03358_);
  and (_03361_, _03360_, _03292_);
  or (_03363_, _03361_, _03357_);
  or (_03365_, _03363_, _03353_);
  and (_03367_, _03365_, _03340_);
  or (_03368_, _03367_, _03339_);
  and (_03370_, _03368_, _03317_);
  and (_03371_, _25525_, _25485_);
  not (_03372_, _25445_);
  nor (_03374_, _03372_, _25402_);
  and (_03375_, _03374_, _03371_);
  and (_03376_, _03375_, _03315_);
  and (_03377_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03378_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03379_, _03378_, _03377_);
  and (_03380_, _03379_, _03300_);
  not (_03381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_03382_, _25707_, _03381_);
  and (_03383_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_03384_, _03383_, _03382_);
  and (_03385_, _03384_, _03286_);
  or (_03386_, _03385_, _03380_);
  not (_03387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_03388_, _25707_, _03387_);
  and (_03389_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03390_, _03389_, _03388_);
  and (_03391_, _03390_, _03292_);
  and (_03392_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03393_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_03394_, _03393_, _03392_);
  and (_03395_, _03394_, _03294_);
  or (_03396_, _03395_, _03391_);
  or (_03397_, _03396_, _03386_);
  and (_03400_, _03397_, _03376_);
  and (_03401_, _25445_, _25402_);
  nor (_03402_, _25525_, _25485_);
  and (_03403_, _03402_, _03401_);
  nor (_03404_, _25707_, _26695_);
  and (_03405_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03406_, _03405_, _03404_);
  and (_03407_, _03406_, _03286_);
  nor (_03408_, _25707_, _26697_);
  and (_03409_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03410_, _03409_, _03408_);
  and (_03411_, _03410_, _03292_);
  or (_03413_, _03411_, _03407_);
  and (_03414_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03415_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_03416_, _03415_, _03414_);
  and (_03418_, _03416_, _03300_);
  and (_03419_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03421_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03422_, _03421_, _03419_);
  and (_03423_, _03422_, _03294_);
  or (_03424_, _03423_, _03418_);
  or (_03425_, _03424_, _03413_);
  and (_03427_, _03425_, _03315_);
  and (_03428_, _03427_, _03403_);
  or (_03429_, _03428_, _03400_);
  or (_03430_, _03429_, _03370_);
  nand (_03431_, _03401_, _03315_);
  not (_03432_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_03433_, _03157_, _03432_);
  and (_03434_, _03433_, _03431_);
  and (_03436_, _03316_, _25301_);
  not (_03437_, _03436_);
  nor (_03438_, _03437_, _03154_);
  nor (_03439_, _03438_, _03376_);
  and (_03440_, _03439_, _03434_);
  and (_03441_, _03318_, _03156_);
  and (_03442_, _03441_, _03315_);
  nor (_03443_, _25707_, _02136_);
  and (_03444_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03446_, _03444_, _03443_);
  and (_03447_, _03446_, _03292_);
  nor (_03448_, _25707_, _02042_);
  and (_03449_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_03450_, _03449_, _03448_);
  and (_03452_, _03450_, _03300_);
  not (_03453_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_03455_, _25707_, _03453_);
  and (_03456_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03457_, _03456_, _03455_);
  and (_03459_, _03457_, _03286_);
  or (_03461_, _03459_, _03452_);
  nor (_03462_, _25707_, _02043_);
  and (_03463_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_03464_, _03463_, _03462_);
  and (_03465_, _03464_, _03294_);
  or (_03467_, _03465_, _03461_);
  or (_03468_, _03467_, _03447_);
  and (_03469_, _03468_, _03442_);
  or (_03471_, _03469_, _03440_);
  or (_03472_, _03471_, _03430_);
  or (_03474_, _03472_, _03314_);
  nor (_03475_, _25525_, _25402_);
  and (_03476_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03477_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03478_, _03477_, _03476_);
  and (_03479_, _03478_, _03294_);
  and (_03480_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03481_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_03483_, _03481_, _03480_);
  and (_03484_, _03483_, _03286_);
  and (_03485_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_03486_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03487_, _03486_, _03485_);
  and (_03488_, _03487_, _03300_);
  or (_03489_, _03488_, _03484_);
  and (_03490_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03491_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03492_, _03491_, _03490_);
  and (_03493_, _03492_, _03292_);
  or (_03494_, _03493_, _03489_);
  or (_03495_, _03494_, _03479_);
  and (_03496_, _03495_, _03157_);
  nor (_03497_, _25707_, _23284_);
  and (_03498_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03499_, _03498_, _03497_);
  and (_03500_, _03499_, _03294_);
  nor (_03501_, _25707_, _23573_);
  and (_03502_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03504_, _03502_, _03501_);
  and (_03505_, _03504_, _03300_);
  nor (_03507_, _25707_, _23351_);
  and (_03509_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03511_, _03509_, _03507_);
  and (_03513_, _03511_, _03286_);
  or (_03514_, _03513_, _03505_);
  nor (_03515_, _25707_, _23319_);
  and (_03517_, _25707_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03518_, _03517_, _03515_);
  and (_03519_, _03518_, _03292_);
  or (_03520_, _03519_, _03514_);
  or (_03521_, _03520_, _03500_);
  and (_03522_, _03521_, _03436_);
  or (_03523_, _03522_, _03496_);
  and (_03524_, _03523_, _03475_);
  and (_03526_, _01873_, _22994_);
  not (_03527_, _03526_);
  and (_03528_, _03527_, _25081_);
  and (_03530_, _23000_, _22993_);
  not (_03532_, _03530_);
  and (_03534_, _25110_, _22939_);
  nor (_03535_, _03534_, _25099_);
  and (_03536_, _03535_, _03532_);
  not (_03537_, _25107_);
  and (_03538_, _22993_, _24143_);
  nor (_03539_, _03538_, _01900_);
  and (_03540_, _03539_, _01903_);
  and (_03541_, _03540_, _03537_);
  and (_03542_, _03541_, _03536_);
  not (_03543_, _01905_);
  nor (_03544_, _03543_, _25087_);
  and (_03545_, _03544_, _01880_);
  and (_03546_, _03545_, _03542_);
  and (_03547_, _03546_, _25078_);
  and (_03548_, _03547_, _03528_);
  nor (_03549_, _03548_, _23061_);
  or (_03550_, _03549_, p1_in[4]);
  not (_03551_, _03549_);
  or (_03552_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03554_, _03552_, _03550_);
  and (_03557_, _03554_, _03290_);
  nor (_03558_, _03549_, p1_in[0]);
  and (_03560_, _03549_, _01585_);
  nor (_03561_, _03560_, _03558_);
  and (_03562_, _03561_, _25707_);
  or (_03563_, _03562_, _03557_);
  and (_03564_, _03563_, _03286_);
  or (_03565_, _03549_, p1_in[7]);
  or (_03567_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03568_, _03567_, _03565_);
  and (_03569_, _03568_, _03290_);
  or (_03570_, _03549_, p1_in[3]);
  or (_03571_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_03572_, _03571_, _03570_);
  and (_03573_, _03572_, _25707_);
  or (_03575_, _03573_, _03569_);
  and (_03576_, _03575_, _03294_);
  or (_03578_, _03576_, _03564_);
  or (_03579_, _03549_, p1_in[5]);
  or (_03580_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03581_, _03580_, _03579_);
  and (_03582_, _03581_, _03290_);
  or (_03583_, _03549_, p1_in[1]);
  or (_03584_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03586_, _03584_, _03583_);
  and (_03588_, _03586_, _25707_);
  or (_03590_, _03588_, _03582_);
  and (_03591_, _03590_, _03292_);
  or (_03592_, _03549_, p1_in[6]);
  or (_03593_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_03596_, _03593_, _03592_);
  and (_03597_, _03596_, _03290_);
  or (_03598_, _03549_, p1_in[2]);
  or (_03599_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03601_, _03599_, _03598_);
  and (_03603_, _03601_, _25707_);
  or (_03604_, _03603_, _03597_);
  and (_03606_, _03604_, _03300_);
  or (_03607_, _03606_, _03591_);
  or (_03608_, _03607_, _03578_);
  and (_03609_, _03608_, _03157_);
  or (_03611_, _03549_, p0_in[4]);
  or (_03612_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_03614_, _03612_, _03611_);
  and (_03616_, _03614_, _03290_);
  nor (_03618_, _03549_, p0_in[0]);
  and (_03619_, _03549_, _01866_);
  nor (_03620_, _03619_, _03618_);
  and (_03621_, _03620_, _25707_);
  or (_03622_, _03621_, _03616_);
  and (_03623_, _03622_, _03286_);
  or (_03624_, _03549_, p0_in[7]);
  or (_03625_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03627_, _03625_, _03624_);
  and (_03628_, _03627_, _03290_);
  or (_03630_, _03549_, p0_in[3]);
  or (_03631_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03633_, _03631_, _03630_);
  and (_03634_, _03633_, _25707_);
  or (_03635_, _03634_, _03628_);
  and (_03636_, _03635_, _03294_);
  or (_03637_, _03636_, _03623_);
  or (_03638_, _03549_, p0_in[5]);
  or (_03639_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03640_, _03639_, _03638_);
  and (_03642_, _03640_, _03290_);
  or (_03643_, _03549_, p0_in[1]);
  or (_03644_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03645_, _03644_, _03643_);
  and (_03646_, _03645_, _25707_);
  or (_03647_, _03646_, _03642_);
  and (_03648_, _03647_, _03292_);
  or (_03649_, _03549_, p0_in[6]);
  or (_03650_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_03651_, _03650_, _03649_);
  and (_03652_, _03651_, _03290_);
  or (_03653_, _03549_, p0_in[2]);
  or (_03654_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_03655_, _03654_, _03653_);
  and (_03656_, _03655_, _25707_);
  or (_03657_, _03656_, _03652_);
  and (_03658_, _03657_, _03300_);
  or (_03659_, _03658_, _03648_);
  or (_03660_, _03659_, _03637_);
  and (_03661_, _03660_, _03436_);
  or (_03662_, _03661_, _03609_);
  and (_03663_, _03662_, _03318_);
  or (_03664_, _03549_, p3_in[4]);
  or (_03665_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_03666_, _03665_, _03664_);
  and (_03668_, _03666_, _03290_);
  nor (_03669_, _03549_, p3_in[0]);
  and (_03671_, _03549_, _00440_);
  nor (_03672_, _03671_, _03669_);
  and (_03674_, _03672_, _25707_);
  or (_03675_, _03674_, _03668_);
  and (_03677_, _03675_, _03286_);
  or (_03678_, _03549_, p3_in[7]);
  or (_03679_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03681_, _03679_, _03678_);
  and (_03683_, _03681_, _03290_);
  or (_03684_, _03549_, p3_in[3]);
  or (_03685_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03686_, _03685_, _03684_);
  and (_03687_, _03686_, _25707_);
  or (_03688_, _03687_, _03683_);
  and (_03689_, _03688_, _03294_);
  or (_03690_, _03689_, _03677_);
  or (_03691_, _03549_, p3_in[5]);
  or (_03693_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03694_, _03693_, _03691_);
  and (_03695_, _03694_, _03290_);
  or (_03696_, _03549_, p3_in[1]);
  or (_03697_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03698_, _03697_, _03696_);
  and (_03699_, _03698_, _25707_);
  or (_03700_, _03699_, _03695_);
  and (_03701_, _03700_, _03292_);
  or (_03702_, _03549_, p3_in[6]);
  or (_03703_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03704_, _03703_, _03702_);
  and (_03705_, _03704_, _03290_);
  or (_03706_, _03549_, p3_in[2]);
  or (_03707_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03708_, _03707_, _03706_);
  and (_03709_, _03708_, _25707_);
  or (_03710_, _03709_, _03705_);
  and (_03711_, _03710_, _03300_);
  or (_03712_, _03711_, _03701_);
  or (_03713_, _03712_, _03690_);
  and (_03714_, _03713_, _03157_);
  or (_03715_, _03549_, p2_in[4]);
  or (_03716_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_03717_, _03716_, _03715_);
  and (_03718_, _03717_, _03290_);
  nor (_03719_, _03549_, p2_in[0]);
  and (_03721_, _03549_, _01457_);
  nor (_03722_, _03721_, _03719_);
  and (_03723_, _03722_, _25707_);
  or (_03724_, _03723_, _03718_);
  and (_03725_, _03724_, _03286_);
  or (_03726_, _03549_, p2_in[7]);
  or (_03728_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03729_, _03728_, _03726_);
  and (_03730_, _03729_, _03290_);
  or (_03731_, _03549_, p2_in[3]);
  or (_03732_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_03733_, _03732_, _03731_);
  and (_03734_, _03733_, _25707_);
  or (_03735_, _03734_, _03730_);
  and (_03736_, _03735_, _03294_);
  or (_03737_, _03736_, _03725_);
  or (_03739_, _03549_, p2_in[5]);
  or (_03740_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03741_, _03740_, _03739_);
  and (_03742_, _03741_, _03290_);
  or (_03744_, _03549_, p2_in[1]);
  or (_03746_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_03747_, _03746_, _03744_);
  and (_03748_, _03747_, _25707_);
  or (_03750_, _03748_, _03742_);
  and (_03751_, _03750_, _03292_);
  or (_03752_, _03549_, p2_in[6]);
  or (_03753_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03754_, _03753_, _03752_);
  and (_03755_, _03754_, _03290_);
  or (_03756_, _03549_, p2_in[2]);
  or (_03757_, _03551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_03758_, _03757_, _03756_);
  and (_03759_, _03758_, _25707_);
  or (_03760_, _03759_, _03755_);
  and (_03761_, _03760_, _03300_);
  or (_03762_, _03761_, _03751_);
  or (_03764_, _03762_, _03737_);
  and (_03766_, _03764_, _03436_);
  or (_03767_, _03766_, _03714_);
  and (_03768_, _03767_, _03340_);
  or (_03769_, _03768_, _03663_);
  or (_03770_, _03769_, _03524_);
  or (_03771_, _03770_, _03474_);
  or (_03772_, _03771_, _03313_);
  and (_03773_, _03475_, _03436_);
  and (_03774_, _03773_, _25610_);
  nor (_03775_, _03774_, _25538_);
  nand (_03776_, _03314_, _23729_);
  and (_03777_, _03776_, _03775_);
  and (_03778_, _03777_, _03772_);
  nor (_03779_, _25707_, _25417_);
  and (_03780_, _25707_, _02075_);
  or (_03781_, _03780_, _03779_);
  and (_03783_, _03781_, _03294_);
  nor (_03784_, _25707_, _25332_);
  and (_03786_, _25707_, _25258_);
  or (_03787_, _03786_, _03784_);
  and (_03788_, _03787_, _03300_);
  nor (_03789_, _25707_, _23824_);
  and (_03790_, _25707_, _25283_);
  or (_03791_, _03790_, _03789_);
  and (_03792_, _03791_, _03286_);
  or (_03793_, _03792_, _03788_);
  nor (_03795_, _25707_, _25362_);
  and (_03796_, _25707_, _02041_);
  or (_03797_, _03796_, _03795_);
  and (_03798_, _03797_, _03292_);
  or (_03799_, _03798_, _03793_);
  nor (_03800_, _03799_, _03783_);
  nor (_03801_, _03800_, _03775_);
  or (_03802_, _03801_, _03778_);
  and (_27329_, _03802_, _23049_);
  nor (_03803_, _25525_, _03155_);
  and (_03804_, _25707_, _25301_);
  and (_03805_, _03804_, _03286_);
  and (_03806_, _03805_, _03374_);
  and (_03807_, _03806_, _03803_);
  and (_03808_, _03807_, _25610_);
  not (_03809_, _26470_);
  and (_03810_, _03294_, _03290_);
  nor (_03811_, _03810_, _03809_);
  and (_03812_, _03811_, _25532_);
  nor (_03813_, _03812_, _03808_);
  and (_03814_, _03813_, _25760_);
  and (_03815_, _03807_, _25606_);
  and (_03816_, _25525_, _03155_);
  and (_03817_, _03806_, _03816_);
  and (_03818_, _03817_, _25626_);
  and (_03819_, _25609_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_03820_, _03318_, _03316_);
  and (_03821_, _03820_, _03294_);
  and (_03822_, _03821_, _03804_);
  and (_03823_, _03822_, _03819_);
  or (_03824_, _03823_, _03818_);
  nor (_03825_, _03824_, _03815_);
  nor (_03827_, _03825_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_03828_, _03827_);
  and (_03829_, _03828_, _03814_);
  and (_03830_, _03820_, _03300_);
  and (_03831_, _03830_, _03804_);
  and (_03832_, _03831_, _03819_);
  or (_03833_, _03832_, rst);
  nor (_27330_, _03833_, _03829_);
  nor (_03834_, _25707_, _25301_);
  and (_03835_, _03834_, _03286_);
  and (_03836_, _03835_, _03375_);
  and (_03837_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_03838_, _25707_, _03315_);
  and (_03839_, _03838_, _03286_);
  and (_03840_, _03839_, _03375_);
  and (_03841_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_03842_, _03841_, _03837_);
  and (_03843_, _03838_, _03300_);
  and (_03845_, _03843_, _03375_);
  and (_03846_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_03847_, _03834_, _03292_);
  and (_03848_, _03847_, _03375_);
  and (_03849_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03851_, _03849_, _03846_);
  or (_03852_, _03851_, _03842_);
  and (_03853_, _03838_, _03294_);
  and (_03854_, _03853_, _03375_);
  and (_03855_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03856_, _03839_, _03820_);
  and (_03858_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03859_, _03858_, _03855_);
  and (_03860_, _03810_, _25301_);
  and (_03861_, _03860_, _03403_);
  and (_03862_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03863_, _03803_, _03401_);
  and (_03864_, _03863_, _03839_);
  and (_03865_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03867_, _03865_, _03862_);
  or (_03868_, _03867_, _03859_);
  or (_03869_, _03868_, _03852_);
  and (_03870_, _03838_, _03292_);
  and (_03871_, _03870_, _03820_);
  and (_03872_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_03873_, _03853_, _03820_);
  and (_03874_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_03875_, _03874_, _03872_);
  and (_03876_, _03843_, _03820_);
  and (_03877_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_03878_, _03847_, _03820_);
  and (_03879_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_03880_, _03879_, _03877_);
  or (_03881_, _03880_, _03875_);
  and (_03882_, _03835_, _03820_);
  and (_03884_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03885_, _03860_, _03820_);
  and (_03887_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03888_, _03887_, _03884_);
  and (_03889_, _03870_, _03441_);
  and (_03890_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03891_, _03839_, _03441_);
  and (_03892_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03893_, _03892_, _03890_);
  or (_03895_, _03893_, _03888_);
  or (_03896_, _03895_, _03881_);
  or (_03897_, _03896_, _03869_);
  and (_03898_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_03899_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_03900_, _03899_, _03898_);
  and (_03902_, _03804_, _03292_);
  and (_03904_, _03902_, _03820_);
  and (_03905_, _03904_, _25419_);
  and (_03906_, _03806_, _03402_);
  and (_03907_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_03908_, _03907_, _03905_);
  or (_03909_, _03908_, _03900_);
  and (_03910_, _03805_, _03403_);
  and (_03911_, _03910_, _03681_);
  and (_03912_, _03863_, _03805_);
  and (_03913_, _03912_, _03729_);
  or (_03914_, _03913_, _03911_);
  and (_03915_, _03805_, _03441_);
  and (_03916_, _03915_, _03568_);
  and (_03917_, _03820_, _03805_);
  and (_03918_, _03917_, _03627_);
  or (_03919_, _03918_, _03916_);
  or (_03920_, _03919_, _03914_);
  or (_03922_, _03920_, _03909_);
  and (_03924_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03925_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03926_, _03925_, _03924_);
  or (_03927_, _03926_, _03922_);
  or (_03928_, _03927_, _03897_);
  and (_03929_, _03928_, _03829_);
  not (_03930_, _03829_);
  not (_03931_, _03891_);
  not (_03932_, _03839_);
  and (_03933_, _03316_, _03153_);
  nand (_03934_, _03933_, _25402_);
  or (_03935_, _03934_, _03932_);
  and (_03936_, _03935_, _03931_);
  and (_03938_, _03821_, _25707_);
  nor (_03939_, _03938_, _03889_);
  and (_03940_, _03939_, _03936_);
  nor (_03941_, _03885_, _03861_);
  nor (_03943_, _03845_, _03904_);
  and (_03944_, _03943_, _03941_);
  not (_03945_, _03831_);
  nand (_03946_, _03805_, _03401_);
  and (_03947_, _03946_, _03945_);
  nor (_03948_, _03848_, _03882_);
  and (_03949_, _03948_, _03947_);
  and (_03950_, _03949_, _03944_);
  nor (_03951_, _03876_, _03836_);
  not (_03952_, _03371_);
  and (_03954_, _03806_, _03952_);
  nor (_03955_, _03954_, _03854_);
  and (_03956_, _03955_, _03951_);
  nor (_03957_, _03878_, _03840_);
  nor (_03958_, _03871_, _03856_);
  and (_03960_, _03958_, _03957_);
  and (_03961_, _03960_, _03956_);
  and (_03962_, _03961_, _03950_);
  and (_03963_, _03962_, _03940_);
  or (_03964_, _03963_, _03930_);
  and (_03965_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03966_, _03965_, _03929_);
  or (_03967_, _03966_, _03832_);
  not (_03968_, _03832_);
  or (_03969_, _03968_, _25053_);
  and (_03970_, _03969_, _23049_);
  and (_27331_[7], _03970_, _03967_);
  and (_26892_[4], _22968_, _23049_);
  nor (_26892_[0], _22830_, rst);
  nor (_26892_[1], _22855_, rst);
  and (_26892_[2], _22777_, _23049_);
  and (_26892_[3], _22804_, _23049_);
  nor (_26892_[5], _22883_, rst);
  and (_03974_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  and (_03975_, _00418_, _26170_);
  or (_25527_, _03975_, _03974_);
  and (_03976_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_03977_, _02879_, _23830_);
  or (_25546_, _03977_, _03976_);
  nor (_26928_[5], _24301_, rst);
  nor (_26928_[1], _24456_, rst);
  nor (_26928_[2], _24417_, rst);
  nor (_26928_[3], _24378_, rst);
  nor (_26928_[4], _24340_, rst);
  nor (_26929_[5], _24286_, rst);
  nor (_26929_[1], _24440_, rst);
  nor (_26929_[2], _24401_, rst);
  nor (_26929_[3], _24361_, rst);
  nor (_26929_[4], _24325_, rst);
  nor (_26929_[6], _24247_, rst);
  and (_03981_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_03982_, _02879_, _25927_);
  or (_25676_, _03982_, _03981_);
  and (_03983_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_03984_, _02879_, _23768_);
  or (_25690_, _03984_, _03983_);
  and (_03985_, _01871_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_03986_, _25070_, _25088_);
  and (_03987_, _23018_, _22949_);
  and (_03988_, _01898_, _23017_);
  or (_03989_, _03988_, _25100_);
  or (_03990_, _03989_, _03987_);
  or (_03991_, _03990_, _03986_);
  or (_03993_, _24152_, _22977_);
  and (_03994_, _25071_, _22989_);
  and (_03995_, _24146_, _22989_);
  or (_03997_, _03995_, _01896_);
  nor (_03999_, _03997_, _03994_);
  nand (_04000_, _03999_, _03544_);
  or (_04001_, _04000_, _03993_);
  or (_04002_, _04001_, _03991_);
  and (_04003_, _04002_, _01913_);
  or (_26902_[1], _04003_, _03985_);
  and (_04004_, _26204_, _26150_);
  not (_04005_, _04004_);
  and (_04007_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and (_04008_, _04004_, _23830_);
  or (_25726_, _04008_, _04007_);
  and (_04010_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_04012_, _04004_, _26185_);
  or (_25747_, _04012_, _04010_);
  and (_04014_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_04015_, _04004_, _26085_);
  or (_25765_, _04015_, _04014_);
  and (_04016_, _26224_, _26204_);
  not (_04017_, _04016_);
  and (_04018_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_04019_, _04016_, _23830_);
  or (_25823_, _04019_, _04018_);
  and (_04020_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_04022_, _04016_, _26085_);
  or (_25893_, _04022_, _04020_);
  and (_04024_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_04025_, _04016_, _25927_);
  or (_25929_, _04025_, _04024_);
  and (_04026_, _25126_, _23776_);
  and (_04027_, _04026_, _26072_);
  and (_04029_, _04027_, _26185_);
  not (_04030_, _04027_);
  and (_04031_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or (_27211_, _04031_, _04029_);
  and (_04032_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_04033_, _04016_, _25886_);
  or (_25954_, _04033_, _04032_);
  and (_04035_, _04026_, _25932_);
  and (_04037_, _04035_, _23768_);
  not (_04038_, _04035_);
  and (_04040_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_27209_, _04040_, _04037_);
  and (_04041_, _04026_, _26340_);
  and (_04042_, _04041_, _25886_);
  not (_04044_, _04041_);
  and (_04045_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_25968_, _04045_, _04042_);
  and (_04047_, _04026_, _26150_);
  and (_04048_, _04047_, _26185_);
  not (_04049_, _04047_);
  and (_04050_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or (_25975_, _04050_, _04048_);
  and (_04051_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_04052_, _04016_, _26170_);
  or (_25980_, _04052_, _04051_);
  and (_04053_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_04054_, _04004_, _23768_);
  or (_25986_, _04054_, _04053_);
  and (_04055_, _04026_, _23847_);
  and (_04056_, _04055_, _23768_);
  not (_04057_, _04055_);
  and (_04058_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_25993_, _04058_, _04056_);
  nor (_04059_, _02342_, _23824_);
  and (_04060_, _00190_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_04061_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_04062_, _04061_, _02638_);
  or (_04063_, _04062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_04064_, _04063_, _02656_);
  nor (_04065_, _04064_, _02657_);
  nand (_04066_, _04065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_04067_, _04065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_04068_, _04067_, _04066_);
  and (_04069_, _04068_, _02363_);
  or (_04070_, _04069_, _04060_);
  or (_04071_, _04070_, _04059_);
  and (_25995_, _04071_, _23049_);
  nand (_04072_, _00190_, _25362_);
  nor (_04074_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_04075_, _04074_, _00215_);
  and (_04076_, _04075_, _00197_);
  and (_04077_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_04078_, _04077_, _04076_);
  nor (_04079_, _04078_, _00226_);
  and (_04080_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_04081_, _04080_, _04079_);
  or (_04083_, _04081_, _00190_);
  and (_04084_, _04083_, _23049_);
  and (_26000_, _04084_, _04072_);
  and (_04085_, _04026_, _26258_);
  and (_04086_, _04085_, _26170_);
  not (_04087_, _04085_);
  and (_04089_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_26043_, _04089_, _04086_);
  and (_04090_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_04091_, _04016_, _26242_);
  or (_26064_, _04091_, _04090_);
  and (_04092_, _04026_, _23775_);
  and (_04093_, _04092_, _26085_);
  not (_04094_, _04092_);
  and (_04095_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or (_27191_, _04095_, _04093_);
  and (_04096_, _04026_, _26213_);
  and (_04097_, _04096_, _26185_);
  not (_04098_, _04096_);
  and (_04100_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_27189_, _04100_, _04097_);
  and (_04101_, _04096_, _25927_);
  and (_04103_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_27188_, _04103_, _04101_);
  and (_04105_, _26260_, _25932_);
  not (_04106_, _04105_);
  and (_04107_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_04108_, _04105_, _26185_);
  or (_26091_, _04108_, _04107_);
  and (_04111_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and (_04112_, _04004_, _26170_);
  or (_26101_, _04112_, _04111_);
  and (_04113_, _26340_, _26260_);
  not (_04114_, _04113_);
  and (_04116_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_04117_, _04113_, _25927_);
  or (_26129_, _04117_, _04116_);
  and (_04118_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and (_04119_, _04004_, _25927_);
  or (_26135_, _04119_, _04118_);
  and (_04120_, _26260_, _26224_);
  not (_04121_, _04120_);
  and (_04122_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_04123_, _04120_, _26242_);
  or (_26155_, _04123_, _04122_);
  and (_04125_, _26193_, _23847_);
  and (_04126_, _04125_, _26085_);
  not (_04127_, _04125_);
  and (_04128_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_26169_, _04128_, _04126_);
  and (_04129_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  and (_04130_, _26541_, _25886_);
  or (_27162_, _04130_, _04129_);
  and (_04131_, _04125_, _23830_);
  and (_04132_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_26187_, _04132_, _04131_);
  and (_04134_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_04135_, _26261_, _23768_);
  or (_27164_, _04135_, _04134_);
  and (_04136_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  and (_04137_, _26541_, _23830_);
  or (_26203_, _04137_, _04136_);
  and (_04139_, _04026_, _25914_);
  and (_04140_, _04139_, _23768_);
  not (_04141_, _04139_);
  and (_04142_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or (_27185_, _04142_, _04140_);
  and (_04143_, _26260_, _23220_);
  not (_04145_, _04143_);
  and (_04146_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  and (_04147_, _04143_, _26242_);
  or (_26218_, _04147_, _04146_);
  and (_04148_, _26260_, _26072_);
  not (_04149_, _04148_);
  and (_04150_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  and (_04151_, _04148_, _26185_);
  or (_26223_, _04151_, _04150_);
  and (_04152_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  and (_04153_, _04148_, _25886_);
  or (_26226_, _04153_, _04152_);
  and (_04155_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  and (_04156_, _04143_, _25886_);
  or (_26229_, _04156_, _04155_);
  and (_04157_, _25126_, _23223_);
  and (_04159_, _04157_, _26258_);
  and (_04160_, _04159_, _25927_);
  not (_04161_, _04159_);
  and (_04162_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_26232_, _04162_, _04160_);
  and (_04163_, _04157_, _26374_);
  and (_04164_, _04163_, _26170_);
  not (_04165_, _04163_);
  and (_04166_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  or (_26238_, _04166_, _04164_);
  and (_04167_, _04163_, _26242_);
  and (_04169_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or (_27142_, _04169_, _04167_);
  and (_04170_, _04159_, _23768_);
  and (_04172_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_27143_, _04172_, _04170_);
  and (_04175_, _26283_, _26193_);
  and (_04176_, _04175_, _23768_);
  not (_04177_, _04175_);
  and (_04179_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_26251_, _04179_, _04176_);
  and (_04181_, _04026_, _23220_);
  and (_04182_, _04181_, _23830_);
  not (_04184_, _04181_);
  and (_04185_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or (_26253_, _04185_, _04182_);
  and (_04187_, _04125_, _26242_);
  and (_04189_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_26259_, _04189_, _04187_);
  and (_04190_, _04035_, _26185_);
  and (_04192_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_26266_, _04192_, _04190_);
  and (_04194_, _04026_, _26224_);
  and (_04195_, _04194_, _23768_);
  not (_04196_, _04194_);
  and (_04197_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_26272_, _04197_, _04195_);
  and (_04198_, _04026_, _26374_);
  and (_04199_, _04198_, _23830_);
  not (_04200_, _04198_);
  and (_04201_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or (_26274_, _04201_, _04199_);
  and (_04202_, _04026_, _26190_);
  and (_04203_, _04202_, _23830_);
  not (_04204_, _04202_);
  and (_04205_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_26280_, _04205_, _04203_);
  not (_04206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_04207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  nor (_04208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_04209_, _04208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_04210_, _04209_, _03381_);
  and (_04211_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02042_);
  or (_04212_, _04211_, _04210_);
  nor (_04214_, _04212_, _04207_);
  nand (_04215_, _04214_, _04206_);
  nor (_04217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_04218_, _04217_, _04214_);
  nand (_04219_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_04221_, _04219_, _04218_);
  and (_04222_, _04221_, _23049_);
  and (_26282_, _04222_, _04215_);
  and (_04223_, _26258_, _26193_);
  and (_04224_, _04223_, _26242_);
  not (_04226_, _04223_);
  and (_04227_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_27113_, _04227_, _04224_);
  not (_04228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_04230_, _02058_, _04228_);
  and (_04231_, _04230_, _02124_);
  and (_04232_, _04231_, _02121_);
  nand (_04233_, _04232_, _02054_);
  not (_04234_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_04235_, _02126_, _04234_);
  and (_04236_, _04235_, _04233_);
  or (_04237_, _04236_, _02045_);
  and (_26288_, _04237_, _23049_);
  and (_26289_, _04218_, _23049_);
  and (_04240_, _04223_, _26185_);
  and (_04241_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_26300_, _04241_, _04240_);
  and (_04243_, _26260_, _26150_);
  not (_04245_, _04243_);
  and (_04246_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  and (_04247_, _04243_, _26185_);
  or (_26304_, _04247_, _04246_);
  and (_04248_, _02060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_04249_, _04248_, _02045_);
  nor (_04250_, _02046_, rst);
  and (_26306_, _04250_, _04249_);
  and (_04251_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_04252_, _04120_, _25886_);
  or (_26307_, _04252_, _04251_);
  or (_04254_, _02422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_04255_, _02422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_04256_, _04255_, _04254_);
  nand (_04257_, _04256_, _23049_);
  nor (_26309_, _04257_, _02045_);
  and (_04259_, _04223_, _26085_);
  and (_04261_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_26317_, _04261_, _04259_);
  and (_04262_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_04263_, _01608_, _25886_);
  or (_26319_, _04263_, _04262_);
  not (_04265_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_04267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_04269_, _04209_, _03387_);
  or (_04271_, _04269_, _04211_);
  nor (_04272_, _04271_, _04267_);
  nand (_04273_, _04272_, _04265_);
  nor (_04274_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_04275_, _04274_, _04272_);
  nand (_04277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_04278_, _04277_, _04275_);
  and (_04280_, _04278_, _23049_);
  and (_26325_, _04280_, _04273_);
  and (_26328_, _04275_, _23049_);
  and (_04281_, _04125_, _23768_);
  and (_04282_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_27114_, _04282_, _04281_);
  not (_04283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_04284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _03453_);
  not (_04286_, _04284_);
  nor (_04287_, _02050_, _02300_);
  and (_04288_, _04287_, _04286_);
  and (_04290_, _04288_, _02313_);
  nor (_04291_, _04290_, _04283_);
  and (_04292_, _04290_, rxd_i);
  or (_04294_, _04292_, rst);
  or (_26342_, _04294_, _04291_);
  or (_04295_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_04296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04297_, _04296_, _02050_);
  or (_04298_, _04297_, _02272_);
  nand (_04299_, _04298_, _04295_);
  nand (_26344_, _04299_, _01634_);
  and (_04300_, _26260_, _26202_);
  not (_04301_, _04300_);
  and (_04302_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_04303_, _04300_, _25886_);
  or (_26347_, _04303_, _04302_);
  and (_04304_, _04125_, _26170_);
  and (_04305_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or (_26350_, _04305_, _04304_);
  nor (_27328_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04306_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_04307_, _03145_, rst);
  and (_27328_[1], _04307_, _04306_);
  nor (_04308_, _03145_, _03144_);
  or (_04309_, _04308_, _03146_);
  and (_04311_, _03149_, _23049_);
  and (_27328_[2], _04311_, _04309_);
  and (_04313_, _04125_, _25927_);
  and (_04314_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or (_26365_, _04314_, _04313_);
  nand (_04316_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_04318_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_04319_, _04318_, _04316_);
  nand (_04321_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_04322_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_04323_, _04322_, _04321_);
  and (_04325_, _04323_, _04319_);
  nand (_04327_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_04329_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_04330_, _04329_, _04327_);
  nand (_04332_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_04333_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_04334_, _04333_, _04332_);
  and (_04335_, _04334_, _04330_);
  and (_04337_, _04335_, _04325_);
  nand (_04338_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_04339_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_04340_, _04339_, _04338_);
  nand (_04341_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_04342_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_04343_, _04342_, _04341_);
  and (_04344_, _04343_, _04340_);
  nand (_04345_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_04347_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_04348_, _04347_, _04345_);
  nand (_04349_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_04350_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_04351_, _04350_, _04349_);
  and (_04352_, _04351_, _04348_);
  and (_04353_, _04352_, _04344_);
  and (_04355_, _04353_, _04337_);
  nand (_04356_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_04357_, _03804_, _03294_);
  and (_04359_, _04357_, _03820_);
  nand (_04360_, _04359_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_04362_, _04360_, _04356_);
  nand (_04363_, _03904_, _25666_);
  nand (_04364_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_04366_, _04364_, _04363_);
  and (_04367_, _04366_, _04362_);
  nand (_04368_, _03910_, _03672_);
  nand (_04369_, _03912_, _03722_);
  and (_04370_, _04369_, _04368_);
  nand (_04372_, _03915_, _03561_);
  nand (_04373_, _03917_, _03620_);
  and (_04374_, _04373_, _04372_);
  and (_04375_, _04374_, _04370_);
  and (_04376_, _04375_, _04367_);
  not (_04377_, _03817_);
  or (_04378_, _04377_, _03283_);
  nand (_04379_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_04381_, _04379_, _04378_);
  and (_04382_, _04381_, _04376_);
  and (_04383_, _04382_, _04355_);
  nor (_04384_, _04383_, _03930_);
  and (_04385_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_04387_, _04385_, _03832_);
  or (_04388_, _04387_, _04384_);
  or (_04389_, _03968_, _00500_);
  and (_04390_, _04389_, _23049_);
  and (_27331_[0], _04390_, _04388_);
  and (_04391_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_04392_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_04394_, _04392_, _04391_);
  and (_04395_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_04397_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_04398_, _04397_, _04395_);
  or (_04399_, _04398_, _04394_);
  and (_04400_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_04401_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_04402_, _04401_, _04400_);
  and (_04403_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_04404_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_04405_, _04404_, _04403_);
  or (_04406_, _04405_, _04402_);
  or (_04407_, _04406_, _04399_);
  and (_04408_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04409_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_04410_, _04409_, _04408_);
  and (_04411_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_04412_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_04413_, _04412_, _04411_);
  or (_04414_, _04413_, _04410_);
  and (_04415_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_04416_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_04417_, _04416_, _04415_);
  and (_04418_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_04420_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_04421_, _04420_, _04418_);
  or (_04422_, _04421_, _04417_);
  or (_04424_, _04422_, _04414_);
  or (_04425_, _04424_, _04407_);
  and (_04427_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_04428_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_04430_, _04428_, _04427_);
  and (_04431_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_04432_, _03904_, _25720_);
  or (_04433_, _04432_, _04431_);
  or (_04434_, _04433_, _04430_);
  and (_04436_, _03910_, _03698_);
  and (_04437_, _03912_, _03747_);
  or (_04438_, _04437_, _04436_);
  and (_04440_, _03915_, _03586_);
  and (_04441_, _03917_, _03645_);
  or (_04443_, _04441_, _04440_);
  or (_04444_, _04443_, _04438_);
  or (_04445_, _04444_, _04434_);
  and (_04446_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_04448_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04449_, _04448_, _04446_);
  or (_04451_, _04449_, _04445_);
  or (_04453_, _04451_, _04425_);
  and (_04454_, _04453_, _03829_);
  and (_04455_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or (_04457_, _04455_, _04454_);
  or (_04458_, _04457_, _03832_);
  or (_04459_, _03968_, _00557_);
  and (_04460_, _04459_, _23049_);
  and (_27331_[1], _04460_, _04458_);
  and (_04462_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_04463_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_04464_, _04463_, _04462_);
  and (_04465_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_04467_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_04468_, _04467_, _04465_);
  or (_04470_, _04468_, _04464_);
  and (_04471_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_04472_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_04474_, _04472_, _04471_);
  and (_04475_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_04476_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_04477_, _04476_, _04475_);
  or (_04479_, _04477_, _04474_);
  or (_04480_, _04479_, _04470_);
  and (_04481_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04482_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_04483_, _04482_, _04481_);
  and (_04484_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_04485_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_04487_, _04485_, _04484_);
  or (_04488_, _04487_, _04483_);
  and (_04489_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_04490_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_04491_, _04490_, _04489_);
  and (_04492_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_04494_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_04495_, _04494_, _04492_);
  or (_04496_, _04495_, _04491_);
  or (_04497_, _04496_, _04488_);
  or (_04498_, _04497_, _04480_);
  and (_04499_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_04500_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_04502_, _04500_, _04499_);
  and (_04503_, _03904_, _25703_);
  and (_04505_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_04506_, _04505_, _04503_);
  or (_04507_, _04506_, _04502_);
  and (_04508_, _03910_, _03708_);
  and (_04509_, _03912_, _03758_);
  or (_04510_, _04509_, _04508_);
  and (_04511_, _03915_, _03601_);
  and (_04512_, _03917_, _03655_);
  or (_04513_, _04512_, _04511_);
  or (_04514_, _04513_, _04510_);
  or (_04515_, _04514_, _04507_);
  and (_04516_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_04517_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_04519_, _04517_, _04516_);
  or (_04520_, _04519_, _04515_);
  or (_04522_, _04520_, _04498_);
  and (_04523_, _04522_, _03829_);
  and (_04524_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or (_04525_, _04524_, _03832_);
  or (_04526_, _04525_, _04523_);
  nand (_04527_, _03832_, _00608_);
  and (_04529_, _04527_, _23049_);
  and (_27331_[2], _04529_, _04526_);
  and (_04531_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04532_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_04533_, _04532_, _04531_);
  and (_04534_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_04536_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_04537_, _04536_, _04534_);
  or (_04538_, _04537_, _04533_);
  and (_04539_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_04540_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_04541_, _04540_, _04539_);
  and (_04543_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_04545_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_04546_, _04545_, _04543_);
  or (_04547_, _04546_, _04541_);
  or (_04548_, _04547_, _04538_);
  and (_04550_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_04551_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_04552_, _04551_, _04550_);
  and (_04554_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_04555_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_04556_, _04555_, _04554_);
  or (_04558_, _04556_, _04552_);
  and (_04560_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_04561_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_04562_, _04561_, _04560_);
  and (_04564_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_04566_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_04567_, _04566_, _04564_);
  or (_04568_, _04567_, _04562_);
  or (_04569_, _04568_, _04558_);
  or (_04571_, _04569_, _04548_);
  and (_04572_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_04573_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_04575_, _04573_, _04572_);
  not (_04576_, _25295_);
  and (_04577_, _03904_, _04576_);
  and (_04579_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_04580_, _04579_, _04577_);
  or (_04581_, _04580_, _04575_);
  and (_04582_, _03910_, _03686_);
  and (_04584_, _03912_, _03733_);
  or (_04585_, _04584_, _04582_);
  and (_04587_, _03915_, _03572_);
  and (_04588_, _03917_, _03633_);
  or (_04590_, _04588_, _04587_);
  or (_04591_, _04590_, _04585_);
  or (_04592_, _04591_, _04581_);
  and (_04594_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_04595_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_04597_, _04595_, _04594_);
  or (_04598_, _04597_, _04592_);
  or (_04600_, _04598_, _04571_);
  and (_04601_, _04600_, _03829_);
  and (_04602_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or (_04603_, _04602_, _04601_);
  or (_04604_, _04603_, _03832_);
  or (_04605_, _03968_, _00659_);
  and (_04606_, _04605_, _23049_);
  and (_27331_[3], _04606_, _04604_);
  and (_04607_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_04608_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_04609_, _04608_, _04607_);
  and (_04610_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_04611_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_04612_, _04611_, _04610_);
  or (_04613_, _04612_, _04609_);
  and (_04614_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_04615_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_04616_, _04615_, _04614_);
  and (_04617_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_04618_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_04619_, _04618_, _04617_);
  or (_04620_, _04619_, _04616_);
  or (_04621_, _04620_, _04613_);
  and (_04622_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_04624_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_04626_, _04624_, _04622_);
  and (_04627_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_04628_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_04630_, _04628_, _04627_);
  or (_04631_, _04630_, _04626_);
  and (_04632_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_04633_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_04635_, _04633_, _04632_);
  and (_04637_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_04638_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_04640_, _04638_, _04637_);
  or (_04641_, _04640_, _04635_);
  or (_04642_, _04641_, _04631_);
  or (_04643_, _04642_, _04621_);
  and (_04644_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04645_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_04647_, _04645_, _04644_);
  not (_04648_, _25455_);
  and (_04649_, _03904_, _04648_);
  and (_04651_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_04652_, _04651_, _04649_);
  or (_04653_, _04652_, _04647_);
  and (_04654_, _03910_, _03666_);
  and (_04655_, _03912_, _03717_);
  or (_04657_, _04655_, _04654_);
  and (_04658_, _03915_, _03554_);
  and (_04659_, _03917_, _03614_);
  or (_04660_, _04659_, _04658_);
  or (_04661_, _04660_, _04657_);
  or (_04662_, _04661_, _04653_);
  and (_04663_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04664_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_04666_, _04664_, _04663_);
  or (_04667_, _04666_, _04662_);
  or (_04668_, _04667_, _04643_);
  and (_04669_, _04668_, _03829_);
  and (_04670_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_04672_, _04670_, _03832_);
  or (_04673_, _04672_, _04669_);
  or (_04674_, _03968_, _00713_);
  and (_04675_, _04674_, _23049_);
  and (_27331_[4], _04675_, _04673_);
  and (_04676_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_04677_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_04678_, _04677_, _04676_);
  and (_04679_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_04680_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_04681_, _04680_, _04679_);
  or (_04682_, _04681_, _04678_);
  and (_04683_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_04684_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_04686_, _04684_, _04683_);
  and (_04687_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_04688_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_04690_, _04688_, _04687_);
  or (_04691_, _04690_, _04686_);
  or (_04692_, _04691_, _04682_);
  and (_04693_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04694_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_04695_, _04694_, _04693_);
  and (_04696_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_04697_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04698_, _04697_, _04696_);
  or (_04699_, _04698_, _04695_);
  and (_04700_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04701_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04703_, _04701_, _04700_);
  and (_04704_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_04705_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_04706_, _04705_, _04704_);
  or (_04707_, _04706_, _04703_);
  or (_04708_, _04707_, _04699_);
  or (_04709_, _04708_, _04692_);
  and (_04710_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_04712_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_04713_, _04712_, _04710_);
  and (_04714_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_04715_, _25497_);
  and (_04716_, _03904_, _04715_);
  or (_04717_, _04716_, _04714_);
  or (_04718_, _04717_, _04713_);
  and (_04719_, _03910_, _03694_);
  and (_04720_, _03912_, _03741_);
  or (_04721_, _04720_, _04719_);
  and (_04722_, _03915_, _03581_);
  and (_04723_, _03917_, _03640_);
  or (_04724_, _04723_, _04722_);
  or (_04725_, _04724_, _04721_);
  or (_04726_, _04725_, _04718_);
  and (_04727_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_04728_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_04730_, _04728_, _04727_);
  or (_04731_, _04730_, _04726_);
  or (_04732_, _04731_, _04709_);
  and (_04733_, _04732_, _03829_);
  and (_04734_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_04735_, _04734_, _03832_);
  or (_04737_, _04735_, _04733_);
  or (_04738_, _03968_, _00773_);
  and (_04740_, _04738_, _23049_);
  and (_27331_[5], _04740_, _04737_);
  and (_04741_, _03882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_04742_, _03885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_04743_, _04742_, _04741_);
  and (_04744_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_04745_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_04746_, _04745_, _04744_);
  or (_04747_, _04746_, _04743_);
  and (_04748_, _03871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_04749_, _03873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_04750_, _04749_, _04748_);
  and (_04751_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_04752_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_04754_, _04752_, _04751_);
  or (_04755_, _04754_, _04750_);
  or (_04757_, _04755_, _04747_);
  and (_04758_, _03836_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_04760_, _03840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04761_, _04760_, _04758_);
  and (_04762_, _03845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_04763_, _03848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04764_, _04763_, _04762_);
  or (_04765_, _04764_, _04761_);
  and (_04766_, _03856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_04767_, _03854_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04768_, _04767_, _04766_);
  and (_04769_, _03861_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_04770_, _03864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_04771_, _04770_, _04769_);
  or (_04773_, _04771_, _04768_);
  or (_04774_, _04773_, _04765_);
  or (_04775_, _04774_, _04757_);
  and (_04776_, _03831_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_04777_, _03822_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_04778_, _04777_, _04776_);
  and (_04780_, _03906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_04782_, _25374_);
  and (_04783_, _03904_, _04782_);
  or (_04784_, _04783_, _04780_);
  or (_04786_, _04784_, _04778_);
  and (_04787_, _03910_, _03704_);
  and (_04789_, _03912_, _03754_);
  or (_04790_, _04789_, _04787_);
  and (_04791_, _03915_, _03596_);
  and (_04792_, _03917_, _03651_);
  or (_04793_, _04792_, _04791_);
  or (_04795_, _04793_, _04790_);
  or (_04796_, _04795_, _04786_);
  and (_04798_, _03817_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_04800_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04801_, _04800_, _04798_);
  or (_04802_, _04801_, _04796_);
  or (_04803_, _04802_, _04775_);
  and (_04804_, _04803_, _03829_);
  and (_04805_, _03964_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or (_04806_, _04805_, _04804_);
  or (_04807_, _04806_, _03832_);
  or (_04808_, _03968_, _00836_);
  and (_04809_, _04808_, _23049_);
  and (_27331_[6], _04809_, _04807_);
  and (_04810_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  and (_04811_, _04243_, _23830_);
  or (_00040_, _04811_, _04810_);
  and (_04812_, _26213_, _26193_);
  and (_04814_, _04812_, _26085_);
  not (_04815_, _04812_);
  and (_04817_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_00054_, _04817_, _04814_);
  and (_04818_, _02512_, _25886_);
  and (_04819_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_00058_, _04819_, _04818_);
  and (_04820_, _26283_, _23779_);
  not (_04821_, _04820_);
  and (_04822_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_04823_, _04820_, _23768_);
  or (_00062_, _04823_, _04822_);
  and (_04825_, _26374_, _26273_);
  and (_04826_, _04825_, _25927_);
  not (_04827_, _04825_);
  and (_04828_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or (_00075_, _04828_, _04826_);
  and (_04830_, _02329_, _25886_);
  and (_04831_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_00098_, _04831_, _04830_);
  and (_04832_, _04047_, _26242_);
  and (_04833_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or (_27202_, _04833_, _04832_);
  and (_04834_, _04055_, _25927_);
  and (_04835_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_00198_, _04835_, _04834_);
  and (_04836_, _04096_, _26242_);
  and (_04837_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_00233_, _04837_, _04836_);
  or (_04838_, _02682_, _25445_);
  or (_04840_, _04838_, _25485_);
  not (_04841_, _02682_);
  nor (_04843_, _04841_, _25748_);
  not (_04845_, _04843_);
  and (_04847_, _04845_, _04840_);
  and (_04848_, _04847_, _23139_);
  nor (_04849_, _04847_, _23139_);
  or (_04850_, _04849_, _04848_);
  and (_04851_, _04838_, _03155_);
  nor (_04852_, _04851_, _25933_);
  and (_04853_, _04838_, _25525_);
  nor (_04854_, _04853_, _25935_);
  nor (_04855_, _04854_, _04852_);
  not (_04856_, _23224_);
  not (_04857_, _04838_);
  nor (_04858_, _04857_, _25402_);
  nor (_04859_, _04858_, _04856_);
  and (_04860_, _04858_, _04856_);
  nor (_04861_, _04860_, _04859_);
  and (_04862_, _04861_, _04855_);
  and (_04863_, _04862_, _04850_);
  not (_04865_, _23217_);
  nor (_04866_, _04838_, _25525_);
  nor (_04868_, _04841_, _25707_);
  nor (_04870_, _04868_, _04866_);
  nor (_04872_, _04870_, _04865_);
  and (_04873_, _04870_, _04865_);
  nor (_04875_, _04873_, _04872_);
  not (_04876_, _04875_);
  and (_04878_, _04838_, _25301_);
  and (_04879_, _04857_, _25402_);
  nor (_04880_, _04879_, _04878_);
  and (_04881_, _04880_, _23187_);
  nor (_04882_, _04880_, _23187_);
  or (_04884_, _04882_, _04881_);
  nor (_04885_, _04884_, _04876_);
  or (_04886_, _04838_, _25301_);
  or (_04887_, _04841_, _25671_);
  nand (_04888_, _04887_, _04886_);
  and (_04889_, _04888_, _23169_);
  nor (_04890_, _04888_, _23169_);
  nor (_04892_, _04890_, _04889_);
  and (_04893_, _04853_, _25935_);
  not (_04894_, _04893_);
  and (_04895_, _04851_, _25933_);
  not (_04896_, _04895_);
  nor (_04897_, _25448_, _23101_);
  and (_04898_, _04897_, _04896_);
  and (_04899_, _04898_, _04894_);
  and (_04900_, _04899_, _04892_);
  and (_04901_, _04900_, _04885_);
  and (_04902_, _04901_, _04863_);
  and (_26942_, _04902_, _23049_);
  and (_26943_[7], _26241_, _23049_);
  and (_04903_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_04904_, _04105_, _26242_);
  or (_00240_, _04904_, _04903_);
  nor (_26945_[2], _25707_, rst);
  and (_04905_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_04906_, _26261_, _25927_);
  or (_00245_, _04906_, _04905_);
  and (_04907_, _04139_, _25927_);
  and (_04908_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or (_00248_, _04908_, _04907_);
  and (_04909_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  and (_04910_, _00418_, _23830_);
  or (_00262_, _04910_, _04909_);
  and (_04911_, _04035_, _26242_);
  and (_04912_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_27210_, _04912_, _04911_);
  and (_04913_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  and (_04914_, _00089_, _26170_);
  or (_27167_, _04914_, _04913_);
  and (_04915_, _26193_, _26150_);
  and (_04916_, _04915_, _26170_);
  not (_04917_, _04915_);
  and (_04918_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_27120_, _04918_, _04916_);
  and (_04920_, _04163_, _26185_);
  and (_04921_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  or (_00343_, _04921_, _04920_);
  and (_04922_, _04159_, _26185_);
  and (_04923_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_00346_, _04923_, _04922_);
  and (_04924_, _04159_, _25886_);
  and (_04925_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_00386_, _04925_, _04924_);
  and (_26943_[0], _23767_, _23049_);
  and (_26943_[1], _25926_, _23049_);
  and (_26943_[2], _26168_, _23049_);
  and (_26943_[3], _25885_, _23049_);
  and (_26943_[4], _23829_, _23049_);
  and (_26943_[5], _26084_, _23049_);
  and (_26943_[6], _26184_, _23049_);
  nor (_26945_[0], _25671_, rst);
  nor (_26945_[1], _25748_, rst);
  and (_04927_, _04159_, _23830_);
  and (_04928_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_00491_, _04928_, _04927_);
  nor (_04929_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_04930_, _01425_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_04931_, _04930_, _04929_);
  nor (_04932_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04933_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01425_);
  nor (_04934_, _04933_, _04932_);
  nor (_04936_, _00625_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04937_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01425_);
  nor (_04938_, _04937_, _04936_);
  nor (_04939_, _04938_, _04934_);
  not (_04940_, _04939_);
  not (_04941_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_04942_, _00676_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_04943_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01425_);
  nor (_04944_, _04943_, _04942_);
  nor (_04945_, _04944_, _04941_);
  and (_04946_, _04944_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_04948_, _04946_, _04945_);
  nor (_04949_, _04948_, _04940_);
  not (_04950_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_04951_, _04944_, _04950_);
  nor (_04952_, _04944_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04953_, _04952_, _04951_);
  not (_04954_, _04934_);
  and (_04955_, _04938_, _04954_);
  not (_04956_, _04955_);
  nor (_04957_, _04956_, _04953_);
  nor (_04958_, _04957_, _04949_);
  nor (_04959_, _04938_, _04954_);
  not (_04960_, _04959_);
  not (_04961_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_04962_, _04944_, _04961_);
  and (_04963_, _04944_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04964_, _04963_, _04962_);
  nor (_04965_, _04964_, _04960_);
  and (_04966_, _04938_, _04934_);
  not (_04967_, _04966_);
  not (_04968_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_04969_, _04944_, _04968_);
  nor (_04970_, _04944_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_04971_, _04970_, _04969_);
  nor (_04972_, _04971_, _04967_);
  nor (_04973_, _04972_, _04965_);
  and (_04974_, _04973_, _04958_);
  and (_04975_, _04974_, _04931_);
  not (_04976_, _04938_);
  and (_04977_, _04944_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not (_04978_, _04944_);
  and (_04979_, _04978_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_04980_, _04979_, _04977_);
  nor (_04981_, _04980_, _04976_);
  nor (_04982_, _04944_, _04938_);
  and (_04983_, _04982_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04984_, _04944_, _04976_);
  and (_04985_, _04984_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04986_, _04985_, _04983_);
  not (_04987_, _04986_);
  nor (_04988_, _04987_, _04981_);
  nor (_04989_, _04988_, _04934_);
  and (_04990_, _04982_, _04934_);
  and (_04991_, _04990_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_04992_, _04944_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_04993_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04994_, _04944_, _04993_);
  or (_04995_, _04994_, _04992_);
  nor (_04996_, _04995_, _04967_);
  and (_04997_, _04944_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_04998_, _04997_, _04959_);
  or (_04999_, _04998_, _04931_);
  or (_05000_, _04999_, _04996_);
  or (_05001_, _05000_, _04991_);
  nor (_05002_, _05001_, _04989_);
  nor (_05003_, _05002_, _04975_);
  not (_05004_, _05003_);
  and (_05005_, _05004_, word_in[7]);
  not (_05006_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05007_, _04931_, _05006_);
  or (_05008_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05009_, _05008_, _05007_);
  and (_05010_, _05009_, _04966_);
  not (_05011_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05012_, _04931_, _05011_);
  or (_05014_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05015_, _05014_, _05012_);
  and (_05016_, _05015_, _04959_);
  or (_05017_, _05016_, _05010_);
  not (_05018_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_05019_, _04931_, _05018_);
  or (_05020_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05021_, _05020_, _05019_);
  and (_05022_, _05021_, _04955_);
  not (_05023_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_05024_, _04931_, _05023_);
  or (_05025_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05026_, _05025_, _05024_);
  and (_05027_, _05026_, _04939_);
  or (_05028_, _05027_, _05022_);
  or (_05029_, _05028_, _05017_);
  and (_05030_, _05029_, _04944_);
  not (_05031_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_05032_, _04931_, _05031_);
  or (_05033_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05034_, _05033_, _05032_);
  and (_05035_, _05034_, _04955_);
  not (_05036_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_05037_, _04931_, _05036_);
  or (_05038_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_05039_, _05038_, _05037_);
  and (_05040_, _05039_, _04939_);
  or (_05041_, _05040_, _05035_);
  and (_05042_, _05041_, _04978_);
  and (_05044_, _04966_, _04978_);
  not (_05045_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05046_, _04931_, _05045_);
  or (_05047_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05048_, _05047_, _05046_);
  and (_05049_, _05048_, _05044_);
  not (_05051_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_05052_, _04931_, _05051_);
  or (_05053_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05055_, _05053_, _05052_);
  and (_05056_, _05055_, _04990_);
  or (_05057_, _05056_, _05049_);
  or (_05058_, _05057_, _05042_);
  or (_05059_, _05058_, _05030_);
  and (_05060_, _05059_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _05060_, _05005_);
  nor (_05063_, _04934_, _04931_);
  not (_05064_, _05063_);
  and (_05065_, _04934_, _04931_);
  and (_05066_, _05065_, _04938_);
  nor (_05067_, _05065_, _04938_);
  nor (_05068_, _05067_, _05066_);
  not (_05069_, _05068_);
  nor (_05070_, _05069_, _04953_);
  nor (_05071_, _05066_, _04978_);
  nor (_05072_, _04944_, _04976_);
  and (_05073_, _05072_, _05065_);
  nor (_05075_, _05073_, _05071_);
  nor (_05076_, _05075_, _05068_);
  and (_05077_, _05076_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05078_, _05067_, _04944_);
  nor (_05079_, _05078_, _05071_);
  and (_05080_, _05079_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05081_, _05080_, _05077_);
  nor (_05082_, _05081_, _05070_);
  nor (_05083_, _05082_, _05064_);
  nand (_05084_, _05073_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not (_05085_, _05065_);
  nor (_05086_, _05069_, _04980_);
  and (_05087_, _05079_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05088_, _05087_, _05086_);
  or (_05089_, _05088_, _05085_);
  and (_05090_, _05089_, _05084_);
  not (_05091_, _05090_);
  nor (_05092_, _05091_, _05083_);
  and (_05093_, _04954_, _04931_);
  not (_05094_, _05093_);
  and (_05095_, _05068_, _04944_);
  and (_05096_, _05095_, \oc8051_symbolic_cxrom1.regvalid [14]);
  not (_05097_, _05096_);
  and (_05098_, _05079_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05099_, _05076_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05100_, _05068_, _04978_);
  and (_05102_, _05100_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05103_, _05102_, _05099_);
  nor (_05105_, _05103_, _05098_);
  and (_05106_, _05105_, _05097_);
  nor (_05107_, _05106_, _05094_);
  not (_05108_, _04931_);
  and (_05109_, _04934_, _05108_);
  not (_05110_, _05109_);
  and (_05111_, _05100_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05112_, _05076_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05113_, _05095_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05115_, _05079_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05116_, _05115_, _05113_);
  or (_05117_, _05116_, _05112_);
  nor (_05118_, _05117_, _05111_);
  nor (_05119_, _05118_, _05110_);
  nor (_05120_, _05119_, _05107_);
  and (_05121_, _05120_, _05092_);
  or (_05122_, _05065_, _05063_);
  not (_05124_, _05122_);
  not (_05125_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05126_, _04931_, _05125_);
  or (_05127_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_05128_, _05127_, _05126_);
  and (_05129_, _05128_, _05124_);
  not (_05130_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_05131_, _04931_, _05130_);
  or (_05132_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05133_, _05132_, _05131_);
  and (_05134_, _05133_, _05122_);
  or (_05135_, _05134_, _05129_);
  and (_05136_, _05135_, _05076_);
  not (_05138_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_05139_, _04931_, _05138_);
  or (_05140_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_05141_, _05140_, _05139_);
  and (_05142_, _05141_, _05124_);
  not (_05143_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_05144_, _04931_, _05143_);
  or (_05145_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_05146_, _05145_, _05144_);
  and (_05147_, _05146_, _05122_);
  or (_05148_, _05147_, _05142_);
  and (_05149_, _05148_, _05095_);
  or (_05150_, _05149_, _05136_);
  not (_05151_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_05152_, _04931_, _05151_);
  or (_05153_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_05154_, _05153_, _05152_);
  and (_05155_, _05154_, _05122_);
  not (_05156_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_05157_, _04931_, _05156_);
  or (_05158_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_05159_, _05158_, _05157_);
  and (_05160_, _05159_, _05124_);
  or (_05161_, _05160_, _05155_);
  and (_05162_, _05161_, _05079_);
  not (_05163_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_05164_, _04931_, _05163_);
  or (_05165_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_05166_, _05165_, _05164_);
  and (_05167_, _05166_, _05122_);
  not (_05168_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_05169_, _04931_, _05168_);
  or (_05170_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_05171_, _05170_, _05169_);
  and (_05173_, _05171_, _05124_);
  or (_05174_, _05173_, _05167_);
  and (_05175_, _05174_, _05100_);
  or (_05176_, _05175_, _05162_);
  nor (_05177_, _05176_, _05150_);
  nor (_05178_, _05177_, _05121_);
  and (_05179_, _05121_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _05179_, _05178_);
  nor (_05180_, _04966_, _04939_);
  not (_05181_, _05180_);
  nor (_05182_, _05181_, _04953_);
  and (_05183_, _04966_, _04944_);
  nor (_05184_, _04966_, _04944_);
  nor (_05185_, _05184_, _05183_);
  and (_05186_, _05185_, _05181_);
  and (_05187_, _05186_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05188_, _05185_, _05180_);
  and (_05189_, _05188_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05190_, _05189_, _05187_);
  nor (_05191_, _05190_, _05182_);
  nor (_05192_, _05191_, _05085_);
  and (_05193_, _05188_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_05194_, _05193_);
  nor (_05195_, _05181_, _04971_);
  and (_05196_, _05186_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05197_, _05196_, _05195_);
  and (_05198_, _05197_, _05194_);
  nor (_05199_, _05198_, _05094_);
  nor (_05200_, _05199_, _05192_);
  nor (_05201_, _05181_, _04995_);
  and (_05202_, _05186_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05203_, _05188_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05205_, _05203_, _05202_);
  nor (_05206_, _05205_, _05201_);
  nor (_05208_, _05206_, _05064_);
  nor (_05209_, _05181_, _04980_);
  and (_05210_, _05186_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05212_, _05188_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05214_, _05212_, _05210_);
  nor (_05215_, _05214_, _05209_);
  nor (_05216_, _05215_, _05110_);
  nor (_05217_, _05216_, _05208_);
  and (_05218_, _05217_, _05200_);
  not (_05219_, _05185_);
  and (_05220_, _05048_, _04955_);
  and (_05221_, _05055_, _04939_);
  or (_05222_, _05221_, _05220_);
  and (_05223_, _05034_, _04959_);
  and (_05224_, _05039_, _04966_);
  or (_05225_, _05224_, _05223_);
  or (_05226_, _05225_, _05222_);
  and (_05227_, _05226_, _05219_);
  and (_05228_, _05021_, _04959_);
  and (_05229_, _05015_, _04939_);
  or (_05230_, _05229_, _05228_);
  and (_05232_, _05009_, _04955_);
  and (_05234_, _05026_, _04966_);
  or (_05235_, _05234_, _05232_);
  or (_05236_, _05235_, _05230_);
  and (_05237_, _05236_, _05185_);
  nor (_05238_, _05237_, _05227_);
  nor (_05239_, _05238_, _05218_);
  and (_05240_, _05218_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _05240_, _05239_);
  and (_05241_, _05064_, _04938_);
  nor (_05242_, _05064_, _04938_);
  nor (_05245_, _05242_, _05241_);
  not (_05246_, _05245_);
  and (_05247_, _05241_, _04944_);
  nor (_05248_, _05241_, _04944_);
  nor (_05249_, _05248_, _05247_);
  and (_05251_, _05249_, _05246_);
  and (_05252_, _05251_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05253_, _05249_, _05245_);
  and (_05254_, _05253_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05255_, _05246_, _04980_);
  or (_05256_, _05255_, _05254_);
  nor (_05257_, _05256_, _05252_);
  nor (_05258_, _05257_, _05094_);
  and (_05259_, _05251_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05260_, _05246_, _04953_);
  nor (_05261_, _05260_, _05259_);
  nor (_05263_, _05261_, _05110_);
  and (_05264_, _05242_, _04962_);
  or (_05265_, _05264_, _05263_);
  nor (_05266_, _05265_, _05258_);
  and (_05267_, _05251_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_05268_, _05267_);
  nor (_05269_, _04995_, _05246_);
  and (_05270_, _05253_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05271_, _05270_, _05269_);
  and (_05272_, _05271_, _05268_);
  nor (_05274_, _05272_, _05085_);
  and (_05275_, _05251_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05276_, _05246_, _04971_);
  nor (_05277_, _05276_, _05275_);
  nor (_05278_, _05277_, _05064_);
  and (_05279_, _05183_, _05108_);
  and (_05280_, _05279_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05281_, _05280_, _05278_);
  nor (_05282_, _05281_, _05274_);
  and (_05283_, _05282_, _05266_);
  and (_05284_, _05133_, _05124_);
  and (_05285_, _05128_, _05122_);
  or (_05286_, _05285_, _05284_);
  and (_05287_, _05286_, _05251_);
  and (_05288_, _05154_, _05124_);
  and (_05289_, _05159_, _05122_);
  or (_05290_, _05289_, _05288_);
  and (_05292_, _05290_, _05253_);
  and (_05293_, _05245_, _04978_);
  and (_05294_, _05166_, _05124_);
  and (_05295_, _05171_, _05122_);
  or (_05296_, _05295_, _05294_);
  and (_05297_, _05296_, _05293_);
  and (_05299_, _05245_, _04944_);
  and (_05300_, _05146_, _05124_);
  and (_05301_, _05141_, _05122_);
  or (_05302_, _05301_, _05300_);
  and (_05303_, _05302_, _05299_);
  or (_05304_, _05303_, _05297_);
  or (_05305_, _05304_, _05292_);
  nor (_05306_, _05305_, _05287_);
  nor (_05307_, _05306_, _05283_);
  and (_05309_, _05283_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _05309_, _05307_);
  and (_05310_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  and (_05312_, _02576_, _26170_);
  or (_27076_, _05312_, _05310_);
  and (_05313_, _04944_, _04938_);
  or (_05314_, _05313_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_26874_[15], _05314_, _23049_);
  and (_05315_, _05218_, _23049_);
  and (_05316_, _05315_, _05093_);
  and (_05317_, _05180_, _04944_);
  and (_05318_, _05317_, _05316_);
  not (_05319_, _05318_);
  and (_05320_, _05121_, _23049_);
  and (_05321_, _05320_, _05109_);
  and (_05322_, _05321_, _05095_);
  and (_05323_, _04975_, _23049_);
  and (_05324_, _05323_, _04934_);
  nor (_05325_, _05003_, rst);
  and (_05326_, _05325_, _05313_);
  and (_05327_, _05326_, _05324_);
  and (_05328_, _05327_, word_in[7]);
  nor (_05329_, _05327_, _05006_);
  nor (_05330_, _05329_, _05328_);
  nor (_05331_, _05330_, _05322_);
  and (_05332_, _05322_, word_in[15]);
  or (_05333_, _05332_, _05331_);
  and (_05334_, _05333_, _05319_);
  and (_05336_, _05283_, _23049_);
  and (_05337_, _05336_, _05299_);
  and (_05338_, _05337_, _05063_);
  and (_05340_, _05315_, word_in[23]);
  and (_05341_, _05340_, _05318_);
  or (_05342_, _05341_, _05338_);
  or (_05344_, _05342_, _05334_);
  not (_05346_, _05338_);
  and (_05348_, _05336_, word_in[31]);
  or (_05350_, _05348_, _05346_);
  and (_26881_[7], _05350_, _05344_);
  or (_05351_, _05253_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_26891_, _05351_, _23049_);
  and (_05352_, _05066_, _04944_);
  or (_05354_, _04944_, _04940_);
  not (_05355_, _05354_);
  nor (_05356_, _05355_, _05352_);
  nor (_05357_, _05279_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_05358_, _05357_, _05356_);
  and (_26874_[1], _05358_, _23049_);
  or (_05359_, _04944_, _04931_);
  nor (_05360_, _05359_, _04960_);
  nor (_05361_, _05360_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_05362_, _05361_, _05356_);
  and (_26874_[2], _05362_, _23049_);
  and (_05363_, _01627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_05365_, _01614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_05366_, _01618_, _01615_);
  and (_05367_, _05366_, _05365_);
  and (_05368_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_05369_, _05368_, _05367_);
  nor (_05370_, _05369_, _00226_);
  or (_05372_, _05370_, _05363_);
  and (_05373_, _05372_, _01612_);
  nor (_05374_, _01612_, _25279_);
  or (_05375_, _05374_, _05373_);
  and (_00672_, _05375_, _23049_);
  not (_05376_, _05079_);
  and (_05377_, _05065_, _04982_);
  or (_05379_, _05377_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05380_, _05379_, _05376_);
  and (_05382_, _04962_, _04939_);
  or (_05383_, _05382_, _05360_);
  or (_05384_, _05383_, _05380_);
  and (_05385_, _05384_, _05356_);
  and (_05387_, _05379_, _05352_);
  or (_05388_, _05387_, _05355_);
  or (_05389_, _05388_, _05385_);
  and (_26874_[3], _05389_, _23049_);
  and (_05390_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  and (_05392_, _01996_, _23768_);
  or (_00755_, _05392_, _05390_);
  not (_05393_, _04982_);
  and (_05394_, _05072_, _05063_);
  or (_05395_, _05394_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05396_, _05395_, _05393_);
  and (_05397_, _05242_, _04979_);
  or (_05398_, _05094_, _04938_);
  nor (_05399_, _05398_, _04944_);
  or (_05400_, _05399_, _04990_);
  or (_05401_, _05400_, _05397_);
  or (_05402_, _05401_, _05396_);
  and (_26874_[4], _05402_, _23049_);
  and (_05403_, _03115_, _26242_);
  and (_05404_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_00792_, _05404_, _05403_);
  or (_05405_, _05394_, _05377_);
  not (_05406_, _05184_);
  or (_05407_, _05406_, _05405_);
  and (_05408_, _05407_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05409_, _05360_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05410_, _05072_, _05093_);
  not (_05411_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_05412_, _05354_, _05411_);
  or (_05414_, _05412_, _05410_);
  or (_05416_, _05414_, _05409_);
  nor (_05417_, _05416_, _05408_);
  nor (_05418_, _05417_, _05248_);
  nor (_05419_, _05359_, _04940_);
  and (_05420_, _05419_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05421_, _05399_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_05422_, _05421_, _05360_);
  or (_05423_, _05422_, _05420_);
  or (_05424_, _05423_, _05394_);
  or (_05425_, _05424_, _05377_);
  or (_05427_, _05425_, _05418_);
  and (_26874_[5], _05427_, _23049_);
  and (_05428_, _01989_, _26242_);
  and (_05429_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_27260_, _05429_, _05428_);
  and (_05430_, _00249_, _25894_);
  or (_05431_, _05430_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_05432_, _05431_, _25618_);
  nand (_05434_, _05430_, _23729_);
  and (_05435_, _05434_, _05432_);
  not (_05437_, _00257_);
  or (_05438_, _05437_, _25258_);
  or (_05439_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_05441_, _05439_, _25128_);
  and (_05442_, _05441_, _05438_);
  and (_05444_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_05445_, _05444_, rst);
  or (_05447_, _05445_, _05442_);
  or (_00819_, _05447_, _05435_);
  nor (_05449_, _00404_, _01686_);
  nand (_05451_, _05449_, _23729_);
  or (_05452_, _05449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_05453_, _05452_, _25618_);
  and (_05455_, _05453_, _05451_);
  nand (_05456_, _00410_, _25362_);
  or (_05457_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_05458_, _05457_, _25128_);
  and (_05460_, _05458_, _05456_);
  and (_05461_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_05462_, _05461_, rst);
  or (_05463_, _05462_, _05460_);
  or (_00829_, _05463_, _05455_);
  and (_05465_, _02102_, _23768_);
  and (_05466_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or (_00845_, _05466_, _05465_);
  and (_05467_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  and (_05469_, _00418_, _26085_);
  or (_00865_, _05469_, _05467_);
  and (_05470_, _05241_, _04978_);
  or (_05471_, _05071_, _05470_);
  nor (_05472_, _05359_, _04967_);
  not (_05474_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_05475_, _04982_, _05474_);
  and (_05476_, _05475_, _05359_);
  or (_05477_, _05476_, _05472_);
  and (_05478_, _05477_, _05406_);
  and (_05479_, _05405_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05481_, _05479_, _05410_);
  or (_05482_, _05481_, _05478_);
  and (_05483_, _05482_, _05471_);
  or (_05485_, _05479_, _05477_);
  and (_05487_, _05485_, _05352_);
  and (_05488_, _05360_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_05489_, _05354_, _05474_);
  or (_05490_, _05489_, _05377_);
  or (_05491_, _05490_, _05488_);
  or (_05492_, _05491_, _05394_);
  or (_05493_, _05492_, _05487_);
  or (_05494_, _05493_, _05483_);
  and (_26874_[6], _05494_, _23049_);
  and (_05495_, _26341_, _26170_);
  and (_05496_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_00889_, _05496_, _05495_);
  and (_05497_, _00249_, _26473_);
  or (_05498_, _05497_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_05499_, _05498_, _25618_);
  nand (_05500_, _05497_, _23729_);
  and (_05501_, _05500_, _05499_);
  nand (_05502_, _00257_, _25160_);
  or (_05503_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_05505_, _05503_, _25128_);
  and (_05506_, _05505_, _05502_);
  and (_05507_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_05508_, _05507_, rst);
  or (_05510_, _05508_, _05506_);
  or (_00892_, _05510_, _05501_);
  and (_05511_, _00249_, _26130_);
  or (_05512_, _05511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_05513_, _05512_, _25618_);
  nand (_05514_, _05511_, _23729_);
  and (_05515_, _05514_, _05513_);
  nand (_05516_, _00257_, _23824_);
  or (_05517_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_05518_, _05517_, _25128_);
  and (_05519_, _05518_, _05516_);
  and (_05520_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_05522_, _05520_, rst);
  or (_05524_, _05522_, _05519_);
  or (_00923_, _05524_, _05515_);
  and (_05525_, _04982_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_05526_, _05525_, _05394_);
  or (_05528_, _05526_, _05472_);
  or (_05529_, _05066_, _04944_);
  or (_05530_, _05472_, _04944_);
  and (_05531_, _05530_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_05532_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_05533_, _04934_, _05532_);
  and (_05535_, _05533_, _05072_);
  or (_05536_, _05535_, _05073_);
  or (_05538_, _05536_, _05531_);
  or (_05540_, _05538_, _05525_);
  and (_05541_, _05540_, _05529_);
  or (_05542_, _05541_, _05410_);
  or (_05543_, _05542_, _05528_);
  and (_26874_[7], _05543_, _23049_);
  and (_05545_, _26194_, _26170_);
  and (_05546_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or (_00954_, _05546_, _05545_);
  and (_05547_, _26194_, _25927_);
  and (_05548_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_27103_, _05548_, _05547_);
  nor (_05549_, _22948_, _22862_);
  nand (_05550_, _01913_, _23008_);
  or (_26894_[2], _05550_, _05549_);
  and (_05551_, _23848_, _23775_);
  and (_05552_, _05551_, _26242_);
  not (_05553_, _05551_);
  and (_05554_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_27258_, _05554_, _05552_);
  and (_05555_, _01989_, _23768_);
  and (_05556_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_01003_, _05556_, _05555_);
  and (_05557_, _26273_, _25914_);
  and (_05558_, _05557_, _26085_);
  not (_05559_, _05557_);
  and (_05560_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or (_01013_, _05560_, _05558_);
  or (_05561_, _05251_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_26874_[8], _05561_, _23049_);
  not (_05562_, _26089_);
  nor (_05563_, _26138_, _26132_);
  and (_05564_, _05563_, _26104_);
  and (_05565_, _05564_, _05562_);
  or (_05566_, _05565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_05567_, _26119_);
  nand (_05568_, _05565_, _05567_);
  and (_05569_, _05568_, _23049_);
  and (_01069_, _05569_, _05566_);
  and (_01072_, t2ex_i, _23049_);
  nor (_05571_, _26133_, _25417_);
  and (_05572_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_05573_, _05572_, _26120_);
  nand (_05574_, _26110_, _26104_);
  and (_05575_, _05574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_05576_, _05574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_05578_, _05576_, _26093_);
  or (_05580_, _05578_, _05575_);
  or (_05581_, _05580_, _05573_);
  or (_05583_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_05584_, _05583_, _05563_);
  and (_05585_, _05584_, _05581_);
  and (_05586_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_05587_, _05586_, _05585_);
  or (_05588_, _05587_, _05571_);
  and (_01084_, _05588_, _23049_);
  not (_05589_, _05242_);
  and (_05590_, _05071_, _05589_);
  nor (_05591_, _05398_, _04978_);
  not (_05592_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05593_, _05184_, _05592_);
  or (_05594_, _05593_, _05591_);
  and (_05595_, _05594_, _05590_);
  and (_05596_, _05242_, _04944_);
  nor (_05597_, _04944_, _05592_);
  and (_05598_, _05597_, _04966_);
  or (_05599_, _05598_, _05596_);
  or (_05600_, _05599_, _05595_);
  and (_05601_, _05600_, _05071_);
  or (_05602_, _05410_, _05293_);
  and (_05604_, _05602_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05605_, _05594_, _05352_);
  and (_05607_, _05597_, _05242_);
  or (_05608_, _05607_, _05472_);
  or (_05610_, _05608_, _05605_);
  or (_05611_, _05610_, _05604_);
  or (_05612_, _05611_, _05073_);
  or (_05613_, _05612_, _05601_);
  and (_26874_[9], _05613_, _23049_);
  and (_01094_, t2_i, _23049_);
  and (_05615_, _02484_, _25927_);
  and (_05616_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_27100_, _05616_, _05615_);
  and (_05618_, _26118_, _26104_);
  or (_05619_, _05618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_05621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_05623_, _26096_, _05621_);
  nand (_05624_, _05623_, _26120_);
  and (_05625_, _05624_, _05619_);
  or (_05626_, _05625_, _26093_);
  nand (_05628_, _26093_, _05621_);
  and (_05630_, _05628_, _05563_);
  and (_05632_, _05630_, _05626_);
  and (_05633_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_05634_, _05633_, _05632_);
  nor (_05636_, _26142_, _25417_);
  or (_05637_, _05636_, _05634_);
  and (_01100_, _05637_, _23049_);
  not (_05639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_05640_, _05563_, _05639_);
  nor (_05641_, _26093_, _05562_);
  and (_05642_, _05641_, _26119_);
  and (_05644_, _05642_, _05564_);
  or (_05646_, _05644_, _05640_);
  and (_01104_, _05646_, _23049_);
  and (_05648_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_05650_, _26422_, _26242_);
  or (_01107_, _05650_, _05648_);
  and (_05651_, _02484_, _23768_);
  and (_05652_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_01119_, _05652_, _05651_);
  and (_05653_, _26308_, _26170_);
  and (_05654_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_01147_, _05654_, _05653_);
  and (_05655_, _05109_, _05299_);
  not (_05656_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05657_, _05122_, _05656_);
  and (_05658_, _05657_, _05293_);
  or (_05659_, _05658_, _05655_);
  and (_05660_, _05100_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_05661_, _05067_, _05398_);
  and (_05662_, _05661_, _04997_);
  or (_05663_, _05662_, _05660_);
  or (_05664_, _05663_, _05659_);
  or (_05665_, _05073_, _05596_);
  and (_05666_, _05665_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05667_, _05419_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05668_, _05667_, _05666_);
  or (_05669_, _05668_, _05664_);
  and (_05670_, _05071_, _04940_);
  and (_05671_, _05670_, _05669_);
  or (_05672_, _05666_, _05591_);
  or (_05673_, _05672_, _05671_);
  and (_05674_, _05673_, _05590_);
  and (_05675_, _05669_, _05352_);
  and (_05676_, _05180_, _04978_);
  and (_05677_, _05676_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05679_, _05472_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05680_, _05354_, _05656_);
  or (_05682_, _05680_, _05073_);
  or (_05684_, _05682_, _05679_);
  or (_05686_, _05684_, _05596_);
  or (_05687_, _05686_, _05677_);
  or (_05688_, _05687_, _05675_);
  or (_05690_, _05688_, _05674_);
  and (_26874_[10], _05690_, _23049_);
  nand (_05691_, _00069_, _23824_);
  and (_05692_, _01670_, _01667_);
  nand (_05693_, _05692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_05694_, _01654_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_05695_, _05694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_05696_, _05695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_05697_, _05696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not (_05698_, _02497_);
  nand (_05699_, _05698_, _05697_);
  and (_05700_, _05699_, _05693_);
  nor (_05701_, _05700_, _00071_);
  or (_05702_, _05698_, _00071_);
  and (_05703_, _05702_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_05704_, _05703_, _05701_);
  or (_05705_, _05704_, _00069_);
  and (_05706_, _05705_, _23049_);
  and (_01225_, _05706_, _05691_);
  and (_05708_, _26308_, _25927_);
  and (_05709_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_01245_, _05709_, _05708_);
  and (_05711_, _26308_, _23768_);
  and (_05712_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_01254_, _05712_, _05711_);
  and (_05714_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  and (_05715_, _02576_, _25927_);
  or (_01259_, _05715_, _05714_);
  or (_05717_, _05655_, _04960_);
  and (_05718_, _05717_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05719_, _05065_, _05299_);
  and (_05720_, _04990_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05721_, _05720_, _05719_);
  or (_05722_, _05721_, _05718_);
  and (_05723_, _05722_, _05095_);
  and (_05724_, _05124_, _04982_);
  or (_05726_, _05724_, _05078_);
  and (_05727_, _05726_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05728_, _04944_, _04939_);
  and (_05729_, _05728_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05731_, _05729_, _05655_);
  or (_05732_, _05731_, _05727_);
  or (_05733_, _05732_, _05723_);
  and (_05734_, _05733_, _05670_);
  and (_05735_, _05722_, _05352_);
  or (_05736_, _04944_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05738_, _05727_, _05242_);
  and (_05739_, _05738_, _05736_);
  or (_05740_, _05739_, _05735_);
  or (_05741_, _05740_, _05591_);
  or (_05742_, _05741_, _05734_);
  and (_26874_[11], _05742_, _23049_);
  and (_05743_, _01604_, _26170_);
  and (_05744_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_01271_, _05744_, _05743_);
  and (_05745_, _04812_, _26242_);
  and (_05746_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_01325_, _05746_, _05745_);
  and (_05747_, _05247_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05748_, _05072_, _04939_);
  or (_05750_, _05748_, _04990_);
  and (_05751_, _05750_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05752_, _05751_, _05299_);
  or (_05753_, _05752_, _05747_);
  and (_26874_[12], _05753_, _23049_);
  and (_05755_, _26340_, _23848_);
  and (_05757_, _05755_, _26242_);
  not (_05758_, _05755_);
  and (_05759_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_01377_, _05759_, _05757_);
  and (_05761_, _05755_, _26185_);
  and (_05762_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_01382_, _05762_, _05761_);
  and (_05764_, _05755_, _26085_);
  and (_05765_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_01385_, _05765_, _05764_);
  or (_05766_, _05317_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_26874_[13], _05766_, _23049_);
  and (_05768_, _01989_, _26170_);
  and (_05770_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_01412_, _05770_, _05768_);
  and (_05771_, _04157_, _26421_);
  and (_05772_, _05771_, _23830_);
  not (_05773_, _05771_);
  and (_05774_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  or (_27150_, _05774_, _05772_);
  and (_05776_, _03115_, _26170_);
  and (_05777_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_27269_, _05777_, _05776_);
  and (_05779_, _03115_, _25927_);
  and (_05780_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_01434_, _05780_, _05779_);
  or (_05781_, _05095_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_26874_[14], _05781_, _23049_);
  and (_05783_, _02089_, _25536_);
  or (_05784_, _05783_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_05786_, _05784_, _02098_);
  nand (_05787_, _05783_, _23729_);
  and (_05788_, _05787_, _05786_);
  nor (_05790_, _02098_, _25417_);
  or (_05791_, _05790_, _05788_);
  and (_01502_, _05791_, _23049_);
  or (_05792_, _02434_, _02380_);
  and (_05793_, _05792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_05794_, _05793_, _02412_);
  and (_01504_, _05794_, _23049_);
  nor (_01505_, _04208_, rst);
  and (_05795_, _03115_, _23768_);
  and (_05796_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_01508_, _05796_, _05795_);
  and (_05797_, _05771_, _23768_);
  and (_05798_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  or (_01510_, _05798_, _05797_);
  and (_05799_, _26273_, _26213_);
  and (_05800_, _05799_, _23830_);
  not (_05801_, _05799_);
  and (_05802_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_26978_, _05802_, _05800_);
  and (_05804_, _01632_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_05806_, _01634_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01520_, _05806_, _05804_);
  and (_05808_, _05771_, _26170_);
  and (_05809_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or (_01524_, _05809_, _05808_);
  or (_05811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_05812_, _05811_, _23049_);
  and (_05813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_05814_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_05815_, _05814_, rxd_i);
  or (_05816_, _05815_, _05813_);
  and (_05818_, _05816_, _02278_);
  and (_05819_, _02302_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_05820_, _05819_, _05818_);
  and (_05822_, _02289_, rxd_i);
  or (_05823_, _05822_, _02300_);
  or (_05824_, _05823_, _05820_);
  and (_01529_, _05824_, _05812_);
  and (_05826_, _04157_, _23847_);
  and (_05827_, _05826_, _26170_);
  not (_05829_, _05826_);
  and (_05831_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_27144_, _05831_, _05827_);
  and (_05833_, _04159_, _26242_);
  and (_05835_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_01623_, _05835_, _05833_);
  and (_05837_, _05826_, _23768_);
  and (_05838_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_01626_, _05838_, _05837_);
  and (_05839_, _05315_, _05279_);
  not (_05840_, _05839_);
  and (_05841_, _05320_, _05352_);
  not (_05842_, _05841_);
  and (_05843_, _05325_, _04934_);
  nor (_05844_, _05843_, _05323_);
  and (_05846_, _05325_, _04982_);
  and (_05847_, _05846_, _05844_);
  and (_05849_, _05847_, word_in[0]);
  not (_05850_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_05852_, _05847_, _05850_);
  or (_05854_, _05852_, _05849_);
  and (_05855_, _05854_, _05842_);
  and (_05856_, _05841_, word_in[8]);
  or (_05857_, _05856_, _05855_);
  and (_05859_, _05857_, _05840_);
  and (_05860_, _05093_, _05313_);
  and (_05861_, _05336_, _05860_);
  and (_05862_, _05315_, word_in[16]);
  and (_05863_, _05862_, _05279_);
  or (_05864_, _05863_, _05861_);
  or (_05866_, _05864_, _05859_);
  not (_05867_, _05861_);
  or (_05869_, _05867_, word_in[24]);
  and (_26875_[0], _05869_, _05866_);
  and (_05870_, _05336_, word_in[25]);
  and (_05871_, _05870_, _05861_);
  not (_05872_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_05874_, _05847_, _05872_);
  and (_05875_, _05325_, word_in[1]);
  and (_05876_, _05875_, _05847_);
  or (_05878_, _05876_, _05874_);
  or (_05879_, _05878_, _05841_);
  or (_05880_, _05842_, word_in[9]);
  and (_05882_, _05880_, _05879_);
  or (_05883_, _05882_, _05839_);
  or (_05885_, _05840_, word_in[17]);
  and (_05886_, _05885_, _05867_);
  and (_05887_, _05886_, _05883_);
  or (_26875_[1], _05887_, _05871_);
  not (_05889_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_05891_, _05847_, _05889_);
  and (_05892_, _05325_, word_in[2]);
  and (_05893_, _05892_, _05847_);
  or (_05895_, _05893_, _05891_);
  or (_05896_, _05895_, _05841_);
  or (_05897_, _05842_, word_in[10]);
  and (_05898_, _05897_, _05896_);
  or (_05899_, _05898_, _05839_);
  or (_05900_, _05840_, word_in[18]);
  and (_05901_, _05900_, _05867_);
  and (_05902_, _05901_, _05899_);
  and (_05903_, _05336_, word_in[26]);
  and (_05904_, _05903_, _05861_);
  or (_26875_[2], _05904_, _05902_);
  not (_05905_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_05906_, _05847_, _05905_);
  and (_05907_, _05325_, word_in[3]);
  and (_05908_, _05907_, _05847_);
  or (_05909_, _05908_, _05906_);
  or (_05910_, _05909_, _05841_);
  or (_05911_, _05842_, word_in[11]);
  and (_05912_, _05911_, _05910_);
  or (_05913_, _05912_, _05839_);
  or (_05915_, _05840_, word_in[19]);
  and (_05917_, _05915_, _05867_);
  and (_05918_, _05917_, _05913_);
  and (_05919_, _05336_, word_in[27]);
  and (_05920_, _05919_, _05861_);
  or (_26875_[3], _05920_, _05918_);
  and (_05922_, _05839_, word_in[20]);
  and (_05923_, _05847_, word_in[4]);
  not (_05925_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_05926_, _05847_, _05925_);
  or (_05927_, _05926_, _05923_);
  or (_05928_, _05927_, _05841_);
  or (_05929_, _05842_, word_in[12]);
  and (_05930_, _05929_, _05840_);
  and (_05932_, _05930_, _05928_);
  or (_05934_, _05932_, _05922_);
  and (_05935_, _05934_, _05867_);
  and (_05936_, _05861_, word_in[28]);
  or (_26875_[4], _05936_, _05935_);
  not (_05937_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_05938_, _05847_, _05937_);
  and (_05939_, _05325_, word_in[5]);
  and (_05940_, _05939_, _05847_);
  or (_05942_, _05940_, _05938_);
  or (_05943_, _05942_, _05841_);
  or (_05944_, _05842_, word_in[13]);
  and (_05945_, _05944_, _05943_);
  or (_05946_, _05945_, _05839_);
  or (_05947_, _05840_, word_in[21]);
  and (_05948_, _05947_, _05867_);
  and (_05949_, _05948_, _05946_);
  and (_05950_, _05336_, word_in[29]);
  and (_05951_, _05950_, _05861_);
  or (_26875_[5], _05951_, _05949_);
  not (_05953_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_05954_, _05847_, _05953_);
  and (_05955_, _05325_, word_in[6]);
  and (_05957_, _05955_, _05847_);
  or (_05958_, _05957_, _05954_);
  or (_05960_, _05958_, _05841_);
  or (_05961_, _05842_, word_in[14]);
  and (_05963_, _05961_, _05960_);
  or (_05964_, _05963_, _05839_);
  or (_05965_, _05840_, word_in[22]);
  and (_05966_, _05965_, _05867_);
  and (_05967_, _05966_, _05964_);
  and (_05968_, _05336_, word_in[30]);
  and (_05969_, _05968_, _05861_);
  or (_26875_[6], _05969_, _05967_);
  nor (_05970_, _05847_, _05151_);
  and (_05971_, _05325_, word_in[7]);
  and (_05972_, _05847_, _05971_);
  or (_05974_, _05972_, _05970_);
  or (_05975_, _05974_, _05841_);
  or (_05976_, _05842_, word_in[15]);
  and (_05977_, _05976_, _05975_);
  or (_05978_, _05977_, _05839_);
  or (_05980_, _05840_, word_in[23]);
  and (_05981_, _05980_, _05867_);
  and (_05982_, _05981_, _05978_);
  and (_05983_, _05861_, word_in[31]);
  or (_26875_[7], _05983_, _05982_);
  and (_05984_, _01989_, _25927_);
  and (_05985_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_01762_, _05985_, _05984_);
  and (_05988_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_05989_, _04120_, _23830_);
  or (_01766_, _05989_, _05988_);
  and (_05991_, _05336_, _05279_);
  not (_05992_, _05991_);
  and (_05993_, _05315_, _05065_);
  and (_05994_, _05993_, _05188_);
  and (_05995_, _05994_, word_in[16]);
  not (_05996_, _05994_);
  and (_05998_, _05320_, _05063_);
  and (_06000_, _05998_, _05079_);
  and (_06002_, _05325_, word_in[0]);
  and (_06003_, _05325_, _05393_);
  and (_06004_, _05323_, _04954_);
  not (_06005_, _06004_);
  nor (_06006_, _06005_, _06003_);
  and (_06007_, _06006_, _06002_);
  not (_06009_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_06010_, _06006_, _06009_);
  nor (_06011_, _06010_, _06007_);
  nor (_06012_, _06011_, _06000_);
  and (_06013_, _06000_, word_in[8]);
  or (_06014_, _06013_, _06012_);
  and (_06015_, _06014_, _05996_);
  or (_06016_, _06015_, _05995_);
  and (_06017_, _06016_, _05992_);
  and (_06019_, _05991_, word_in[24]);
  or (_26882_[0], _06019_, _06017_);
  not (_06020_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_06021_, _06006_, _06020_);
  and (_06022_, _06006_, _05875_);
  or (_06023_, _06022_, _06021_);
  or (_06024_, _06023_, _06000_);
  not (_06025_, _06000_);
  or (_06026_, _06025_, word_in[9]);
  and (_06027_, _06026_, _06024_);
  or (_06028_, _06027_, _05994_);
  or (_06029_, _05996_, word_in[17]);
  and (_06030_, _06029_, _05992_);
  and (_06032_, _06030_, _06028_);
  and (_06033_, _05991_, word_in[25]);
  or (_26882_[1], _06033_, _06032_);
  and (_06034_, _05994_, word_in[18]);
  and (_06035_, _06006_, _05892_);
  not (_06036_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_06037_, _06006_, _06036_);
  nor (_06038_, _06037_, _06035_);
  nor (_06039_, _06038_, _06000_);
  and (_06040_, _06000_, word_in[10]);
  or (_06041_, _06040_, _06039_);
  and (_06042_, _06041_, _05996_);
  or (_06043_, _06042_, _06034_);
  and (_06044_, _06043_, _05992_);
  and (_06045_, _05991_, word_in[26]);
  or (_26882_[2], _06045_, _06044_);
  and (_06046_, _05994_, word_in[19]);
  and (_06047_, _06006_, _05907_);
  not (_06048_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_06049_, _06006_, _06048_);
  nor (_06051_, _06049_, _06047_);
  nor (_06052_, _06051_, _06000_);
  and (_06054_, _06000_, word_in[11]);
  or (_06055_, _06054_, _06052_);
  and (_06056_, _06055_, _05996_);
  or (_06057_, _06056_, _06046_);
  and (_06058_, _06057_, _05992_);
  and (_06059_, _05991_, word_in[27]);
  or (_26882_[3], _06059_, _06058_);
  and (_06060_, _05994_, word_in[20]);
  and (_06061_, _05325_, word_in[4]);
  and (_06062_, _06006_, _06061_);
  not (_06063_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_06064_, _06006_, _06063_);
  nor (_06066_, _06064_, _06062_);
  nor (_06067_, _06066_, _06000_);
  and (_06069_, _06000_, word_in[12]);
  or (_06070_, _06069_, _06067_);
  and (_06071_, _06070_, _05996_);
  or (_06072_, _06071_, _06060_);
  and (_06073_, _06072_, _05992_);
  and (_06074_, _05991_, word_in[28]);
  or (_26882_[4], _06074_, _06073_);
  and (_06076_, _05994_, word_in[21]);
  and (_06077_, _06006_, _05939_);
  not (_06078_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_06080_, _06006_, _06078_);
  nor (_06081_, _06080_, _06077_);
  nor (_06083_, _06081_, _06000_);
  and (_06084_, _06000_, word_in[13]);
  or (_06085_, _06084_, _06083_);
  and (_06086_, _06085_, _05996_);
  or (_06087_, _06086_, _06076_);
  and (_06088_, _06087_, _05992_);
  and (_06089_, _05991_, word_in[29]);
  or (_26882_[5], _06089_, _06088_);
  not (_06091_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_06092_, _06006_, _06091_);
  and (_06093_, _06006_, _05955_);
  or (_06095_, _06093_, _06092_);
  or (_06096_, _06095_, _06000_);
  or (_06097_, _06025_, word_in[14]);
  and (_06098_, _06097_, _06096_);
  or (_06099_, _06098_, _05994_);
  or (_06101_, _05996_, word_in[22]);
  and (_06102_, _06101_, _05992_);
  and (_06103_, _06102_, _06099_);
  and (_06104_, _05991_, word_in[30]);
  or (_26882_[6], _06104_, _06103_);
  nor (_06106_, _06006_, _05036_);
  and (_06107_, _06006_, _05971_);
  or (_06109_, _06107_, _06106_);
  or (_06110_, _06109_, _06000_);
  or (_06111_, _06025_, word_in[15]);
  and (_06112_, _06111_, _06110_);
  or (_06113_, _06112_, _05994_);
  or (_06114_, _05996_, word_in[23]);
  and (_06115_, _06114_, _05992_);
  and (_06117_, _06115_, _06113_);
  and (_06118_, _05991_, word_in[31]);
  or (_26882_[7], _06118_, _06117_);
  and (_06119_, _05336_, _05352_);
  not (_06120_, _06119_);
  and (_06121_, _05315_, _05063_);
  and (_06122_, _06121_, _05188_);
  and (_06124_, _06122_, word_in[16]);
  not (_06125_, _06122_);
  and (_06127_, _05320_, _05093_);
  and (_06129_, _06127_, _05079_);
  not (_06130_, _05323_);
  and (_06131_, _05843_, _06130_);
  and (_06132_, _06131_, _04982_);
  and (_06133_, _06132_, _06002_);
  not (_06134_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_06135_, _06132_, _06134_);
  nor (_06136_, _06135_, _06133_);
  nor (_06137_, _06136_, _06129_);
  and (_06138_, _06129_, word_in[8]);
  or (_06139_, _06138_, _06137_);
  and (_06140_, _06139_, _06125_);
  or (_06141_, _06140_, _06124_);
  and (_06142_, _06141_, _06120_);
  and (_06143_, _06119_, word_in[24]);
  or (_26883_[0], _06143_, _06142_);
  and (_06144_, _06122_, word_in[17]);
  and (_06146_, _06132_, _05875_);
  not (_06147_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_06148_, _06132_, _06147_);
  nor (_06149_, _06148_, _06146_);
  nor (_06150_, _06149_, _06129_);
  and (_06151_, _06129_, word_in[9]);
  or (_06152_, _06151_, _06150_);
  and (_06153_, _06152_, _06125_);
  or (_06154_, _06153_, _06144_);
  and (_06155_, _06154_, _06120_);
  and (_06156_, _06119_, word_in[25]);
  or (_26883_[1], _06156_, _06155_);
  and (_06157_, _06132_, _05892_);
  not (_06158_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_06159_, _06132_, _06158_);
  nor (_06160_, _06159_, _06157_);
  nor (_06161_, _06160_, _06129_);
  and (_06162_, _06129_, word_in[10]);
  or (_06163_, _06162_, _06161_);
  and (_06164_, _06163_, _06125_);
  and (_06165_, _06122_, word_in[18]);
  or (_06166_, _06165_, _06119_);
  or (_06167_, _06166_, _06164_);
  or (_06168_, _06120_, word_in[26]);
  and (_26883_[2], _06168_, _06167_);
  and (_06169_, _06119_, word_in[27]);
  not (_06170_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_06171_, _06132_, _06170_);
  and (_06172_, _06132_, _05907_);
  or (_06173_, _06172_, _06171_);
  or (_06174_, _06173_, _06129_);
  not (_06175_, _06129_);
  or (_06176_, _06175_, word_in[11]);
  and (_06178_, _06176_, _06174_);
  or (_06179_, _06178_, _06122_);
  or (_06180_, _06125_, word_in[19]);
  and (_06181_, _06180_, _06120_);
  and (_06182_, _06181_, _06179_);
  or (_26883_[3], _06182_, _06169_);
  and (_06184_, _06132_, _06061_);
  not (_06185_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_06187_, _06132_, _06185_);
  nor (_06189_, _06187_, _06184_);
  nor (_06190_, _06189_, _06129_);
  and (_06191_, _06129_, word_in[12]);
  or (_06193_, _06191_, _06190_);
  and (_06194_, _06193_, _06125_);
  and (_06195_, _06122_, word_in[20]);
  or (_06196_, _06195_, _06119_);
  or (_06198_, _06196_, _06194_);
  or (_06199_, _06120_, word_in[28]);
  and (_26883_[4], _06199_, _06198_);
  and (_06200_, _06132_, _05939_);
  not (_06201_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_06202_, _06132_, _06201_);
  nor (_06203_, _06202_, _06200_);
  nor (_06204_, _06203_, _06129_);
  and (_06206_, _06129_, word_in[13]);
  or (_06207_, _06206_, _06204_);
  and (_06208_, _06207_, _06125_);
  and (_06209_, _06122_, word_in[21]);
  or (_06210_, _06209_, _06119_);
  or (_06212_, _06210_, _06208_);
  or (_06213_, _06120_, word_in[29]);
  and (_26883_[5], _06213_, _06212_);
  not (_06214_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_06215_, _06132_, _06214_);
  and (_06216_, _06132_, _05955_);
  or (_06217_, _06216_, _06215_);
  or (_06218_, _06217_, _06129_);
  or (_06219_, _06175_, word_in[14]);
  and (_06221_, _06219_, _06218_);
  or (_06222_, _06221_, _06122_);
  or (_06223_, _06125_, word_in[22]);
  and (_06224_, _06223_, _06120_);
  and (_06225_, _06224_, _06222_);
  and (_06226_, _06119_, word_in[30]);
  or (_26883_[6], _06226_, _06225_);
  and (_06228_, _06132_, _05971_);
  nor (_06229_, _06132_, _05156_);
  nor (_06230_, _06229_, _06228_);
  nor (_06231_, _06230_, _06129_);
  and (_06232_, _06129_, word_in[15]);
  or (_06233_, _06232_, _06231_);
  and (_06234_, _06233_, _06125_);
  and (_06235_, _06122_, word_in[23]);
  or (_06236_, _06235_, _06119_);
  or (_06237_, _06236_, _06234_);
  or (_06238_, _06120_, word_in[31]);
  and (_26883_[7], _06238_, _06237_);
  and (_06239_, _26176_, _25886_);
  and (_06240_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_01867_, _06240_, _06239_);
  and (_06242_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  and (_06243_, _04148_, _23830_);
  or (_01890_, _06243_, _06242_);
  and (_06244_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_06245_, _04300_, _26170_);
  or (_01906_, _06245_, _06244_);
  and (_06246_, _05336_, _05419_);
  not (_06247_, _06246_);
  and (_06248_, _05316_, _05188_);
  and (_06249_, _06248_, word_in[16]);
  not (_06250_, _06248_);
  and (_06251_, _05321_, _05079_);
  not (_06252_, _05324_);
  nor (_06253_, _06003_, _06252_);
  and (_06254_, _06253_, _06002_);
  not (_06255_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_06256_, _06253_, _06255_);
  nor (_06257_, _06256_, _06254_);
  nor (_06258_, _06257_, _06251_);
  and (_06259_, _06251_, word_in[8]);
  or (_06260_, _06259_, _06258_);
  and (_06261_, _06260_, _06250_);
  or (_06262_, _06261_, _06249_);
  and (_06263_, _06262_, _06247_);
  and (_06264_, _06246_, word_in[24]);
  or (_26884_[0], _06264_, _06263_);
  and (_06265_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_06266_, _04300_, _26085_);
  or (_27181_, _06266_, _06265_);
  and (_06267_, _06248_, word_in[17]);
  and (_06268_, _06253_, _05875_);
  not (_06269_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_06270_, _06253_, _06269_);
  nor (_06271_, _06270_, _06268_);
  nor (_06272_, _06271_, _06251_);
  and (_06273_, _06251_, word_in[9]);
  or (_06274_, _06273_, _06272_);
  and (_06275_, _06274_, _06250_);
  or (_06276_, _06275_, _06267_);
  and (_06277_, _06276_, _06247_);
  and (_06279_, _06246_, word_in[25]);
  or (_26884_[1], _06279_, _06277_);
  and (_06280_, _06253_, _05892_);
  not (_06281_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_06283_, _06253_, _06281_);
  nor (_06285_, _06283_, _06280_);
  nor (_06286_, _06285_, _06251_);
  and (_06287_, _06251_, word_in[10]);
  or (_06289_, _06287_, _06286_);
  and (_06290_, _06289_, _06250_);
  and (_06292_, _06248_, word_in[18]);
  or (_06293_, _06292_, _06246_);
  or (_06296_, _06293_, _06290_);
  or (_06297_, _06247_, word_in[26]);
  and (_26884_[2], _06297_, _06296_);
  and (_06298_, _06253_, _05907_);
  not (_06299_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_06300_, _06253_, _06299_);
  nor (_06301_, _06300_, _06298_);
  nor (_06302_, _06301_, _06251_);
  and (_06303_, _06251_, word_in[11]);
  or (_06304_, _06303_, _06302_);
  and (_06305_, _06304_, _06250_);
  and (_06306_, _06248_, word_in[19]);
  or (_06307_, _06306_, _06246_);
  or (_06308_, _06307_, _06305_);
  or (_06309_, _06247_, word_in[27]);
  and (_26884_[3], _06309_, _06308_);
  and (_06311_, _06253_, _06061_);
  not (_06312_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_06313_, _06253_, _06312_);
  nor (_06314_, _06313_, _06311_);
  nor (_06315_, _06314_, _06251_);
  and (_06316_, _06251_, word_in[12]);
  or (_06317_, _06316_, _06315_);
  and (_06318_, _06317_, _06250_);
  and (_06319_, _06248_, word_in[20]);
  or (_06320_, _06319_, _06246_);
  or (_06322_, _06320_, _06318_);
  or (_06323_, _06247_, word_in[28]);
  and (_26884_[4], _06323_, _06322_);
  and (_06324_, _06253_, _05939_);
  not (_06325_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_06326_, _06253_, _06325_);
  nor (_06327_, _06326_, _06324_);
  nor (_06328_, _06327_, _06251_);
  and (_06329_, _06251_, word_in[13]);
  or (_06330_, _06329_, _06328_);
  and (_06332_, _06330_, _06250_);
  and (_06333_, _06248_, word_in[21]);
  or (_06334_, _06333_, _06246_);
  or (_06335_, _06334_, _06332_);
  or (_06336_, _06247_, word_in[29]);
  and (_26884_[5], _06336_, _06335_);
  and (_06337_, _06253_, _05955_);
  not (_06338_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_06339_, _06253_, _06338_);
  nor (_06340_, _06339_, _06337_);
  nor (_06341_, _06340_, _06251_);
  and (_06342_, _06251_, word_in[14]);
  or (_06343_, _06342_, _06341_);
  and (_06344_, _06343_, _06250_);
  and (_06345_, _06248_, word_in[22]);
  or (_06346_, _06345_, _06246_);
  or (_06347_, _06346_, _06344_);
  or (_06349_, _06247_, word_in[30]);
  and (_26884_[6], _06349_, _06347_);
  and (_06352_, _06253_, _05971_);
  nor (_06353_, _06253_, _05051_);
  nor (_06354_, _06353_, _06352_);
  nor (_06355_, _06354_, _06251_);
  and (_06356_, _06251_, word_in[15]);
  or (_06357_, _06356_, _06355_);
  and (_06359_, _06357_, _06250_);
  and (_06360_, _06248_, word_in[23]);
  or (_06361_, _06360_, _06246_);
  or (_06362_, _06361_, _06359_);
  or (_06363_, _06247_, word_in[31]);
  and (_26884_[7], _06363_, _06362_);
  and (_06364_, _05771_, _26185_);
  and (_06365_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  or (_01945_, _06365_, _06364_);
  and (_06367_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  and (_06368_, _26541_, _26242_);
  or (_01955_, _06368_, _06367_);
  and (_06369_, _26374_, _26260_);
  not (_06370_, _06369_);
  and (_06371_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  and (_06372_, _06369_, _23830_);
  or (_27163_, _06372_, _06371_);
  and (_06373_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  and (_06374_, _06369_, _26185_);
  or (_01974_, _06374_, _06373_);
  and (_06376_, _05336_, _05293_);
  and (_06377_, _06376_, _05093_);
  not (_06378_, _06377_);
  and (_06380_, _05315_, _05180_);
  and (_06382_, _06380_, _05219_);
  and (_06383_, _06382_, _05109_);
  and (_06384_, _06383_, _05862_);
  not (_06385_, _06383_);
  and (_06386_, _05320_, _05377_);
  not (_06387_, _06386_);
  not (_06388_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_06389_, _05325_, _05072_);
  and (_06390_, _06389_, _05844_);
  nor (_06392_, _06390_, _06388_);
  and (_06393_, _06390_, word_in[0]);
  or (_06394_, _06393_, _06392_);
  and (_06395_, _06394_, _06387_);
  and (_06396_, _06386_, word_in[8]);
  or (_06397_, _06396_, _06395_);
  and (_06399_, _06397_, _06385_);
  or (_06400_, _06399_, _06384_);
  and (_06401_, _06400_, _06378_);
  and (_06402_, _06377_, word_in[24]);
  or (_26885_[0], _06402_, _06401_);
  and (_06403_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_06404_, _26261_, _23830_);
  or (_01983_, _06404_, _06403_);
  not (_06405_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_06407_, _06390_, _06405_);
  and (_06408_, _06390_, word_in[1]);
  or (_06410_, _06408_, _06407_);
  and (_06411_, _06410_, _06387_);
  and (_06412_, _06386_, word_in[9]);
  or (_06413_, _06412_, _06411_);
  and (_06414_, _06413_, _06385_);
  and (_06415_, _05315_, word_in[17]);
  and (_06416_, _06383_, _06415_);
  or (_06417_, _06416_, _06377_);
  or (_06418_, _06417_, _06414_);
  or (_06419_, _06378_, _05870_);
  and (_26885_[1], _06419_, _06418_);
  not (_06420_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_06422_, _06390_, _06420_);
  and (_06424_, _06390_, word_in[2]);
  or (_06425_, _06424_, _06422_);
  and (_06427_, _06425_, _06387_);
  and (_06428_, _06386_, word_in[10]);
  or (_06429_, _06428_, _06427_);
  and (_06430_, _06429_, _06385_);
  and (_06431_, _05315_, word_in[18]);
  and (_06432_, _06383_, _06431_);
  or (_06434_, _06432_, _06377_);
  or (_06435_, _06434_, _06430_);
  or (_06436_, _06378_, _05903_);
  and (_26885_[2], _06436_, _06435_);
  and (_06437_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_06438_, _01608_, _26170_);
  or (_01986_, _06438_, _06437_);
  and (_06439_, _05315_, word_in[19]);
  and (_06441_, _06383_, _06439_);
  not (_06442_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_06443_, _06390_, _06442_);
  and (_06444_, _06390_, word_in[3]);
  or (_06445_, _06444_, _06443_);
  and (_06446_, _06445_, _06387_);
  and (_06447_, _06386_, word_in[11]);
  or (_06448_, _06447_, _06446_);
  and (_06449_, _06448_, _06385_);
  or (_06450_, _06449_, _06441_);
  and (_06451_, _06450_, _06378_);
  and (_06452_, _06377_, word_in[27]);
  or (_26885_[3], _06452_, _06451_);
  not (_06453_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_06454_, _06390_, _06453_);
  and (_06455_, _06390_, word_in[4]);
  or (_06456_, _06455_, _06454_);
  and (_06457_, _06456_, _06387_);
  and (_06458_, _06386_, word_in[12]);
  or (_06459_, _06458_, _06457_);
  and (_06460_, _06459_, _06385_);
  and (_06461_, _05315_, word_in[20]);
  and (_06462_, _06383_, _06461_);
  or (_06463_, _06462_, _06377_);
  or (_06464_, _06463_, _06460_);
  and (_06465_, _05336_, word_in[28]);
  or (_06466_, _06378_, _06465_);
  and (_26885_[4], _06466_, _06464_);
  not (_06467_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_06468_, _06390_, _06467_);
  and (_06469_, _06390_, word_in[5]);
  or (_06470_, _06469_, _06468_);
  and (_06471_, _06470_, _06387_);
  and (_06473_, _06386_, word_in[13]);
  or (_06474_, _06473_, _06471_);
  and (_06475_, _06474_, _06385_);
  and (_06477_, _05315_, word_in[21]);
  and (_06478_, _06383_, _06477_);
  or (_06479_, _06478_, _06377_);
  or (_06480_, _06479_, _06475_);
  or (_06481_, _06378_, _05950_);
  and (_26885_[5], _06481_, _06480_);
  not (_06483_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_06484_, _06390_, _06483_);
  and (_06485_, _06390_, word_in[6]);
  or (_06486_, _06485_, _06484_);
  and (_06487_, _06486_, _06387_);
  and (_06488_, _06386_, word_in[14]);
  or (_06489_, _06488_, _06487_);
  and (_06490_, _06489_, _06385_);
  and (_06492_, _05315_, word_in[22]);
  and (_06493_, _06383_, _06492_);
  or (_06494_, _06493_, _06377_);
  or (_06495_, _06494_, _06490_);
  or (_06496_, _06378_, _05968_);
  and (_26885_[6], _06496_, _06495_);
  nor (_06497_, _06390_, _05163_);
  and (_06498_, _06390_, word_in[7]);
  or (_06499_, _06498_, _06497_);
  and (_06500_, _06499_, _06387_);
  and (_06501_, _06386_, word_in[15]);
  or (_06502_, _06501_, _06500_);
  and (_06503_, _06502_, _06385_);
  and (_06505_, _06383_, _05340_);
  or (_06506_, _06505_, _06377_);
  or (_06507_, _06506_, _06503_);
  or (_06508_, _06378_, _05348_);
  and (_26885_[7], _06508_, _06507_);
  and (_06509_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_06510_, _01608_, _26185_);
  or (_01995_, _06510_, _06509_);
  and (_06512_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_06513_, _01608_, _26085_);
  or (_02000_, _06513_, _06512_);
  and (_06514_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  and (_06515_, _00089_, _25927_);
  or (_02005_, _06515_, _06514_);
  and (_06516_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  and (_06517_, _00089_, _26185_);
  or (_02016_, _06517_, _06516_);
  and (_06518_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_06519_, _04120_, _26170_);
  or (_02022_, _06519_, _06518_);
  and (_06520_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_06521_, _04120_, _23768_);
  or (_02027_, _06521_, _06520_);
  and (_06524_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_06526_, _04120_, _26085_);
  or (_02033_, _06526_, _06524_);
  and (_06527_, _06382_, _05065_);
  and (_06528_, _05998_, _05100_);
  and (_06529_, _06389_, _06004_);
  and (_06531_, _06529_, word_in[0]);
  not (_06532_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_06533_, _06529_, _06532_);
  nor (_06534_, _06533_, _06531_);
  nor (_06535_, _06534_, _06528_);
  and (_06537_, _06528_, word_in[8]);
  or (_06538_, _06537_, _06535_);
  or (_06539_, _06538_, _06527_);
  and (_06541_, _06376_, _05109_);
  not (_06542_, _06541_);
  not (_06544_, _06527_);
  or (_06545_, _06544_, _05862_);
  and (_06546_, _06545_, _06542_);
  and (_06548_, _06546_, _06539_);
  and (_06550_, _06541_, word_in[24]);
  or (_26886_[0], _06550_, _06548_);
  and (_06551_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  and (_06552_, _04243_, _26085_);
  or (_02039_, _06552_, _06551_);
  not (_06554_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_06555_, _06529_, _06554_);
  and (_06556_, _06529_, _05875_);
  or (_06557_, _06556_, _06555_);
  or (_06558_, _06557_, _06528_);
  not (_06559_, _06528_);
  or (_06560_, _06559_, word_in[9]);
  and (_06562_, _06560_, _06558_);
  or (_06564_, _06562_, _06527_);
  or (_06566_, _06544_, _06415_);
  and (_06567_, _06566_, _06564_);
  or (_06569_, _06567_, _06541_);
  or (_06570_, _06542_, word_in[25]);
  and (_26886_[1], _06570_, _06569_);
  not (_06572_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_06573_, _06529_, _06572_);
  and (_06574_, _06529_, _05892_);
  or (_06575_, _06574_, _06573_);
  or (_06576_, _06575_, _06528_);
  or (_06577_, _06559_, word_in[10]);
  and (_06578_, _06577_, _06576_);
  or (_06580_, _06578_, _06527_);
  or (_06581_, _06544_, _06431_);
  and (_06583_, _06581_, _06542_);
  and (_06585_, _06583_, _06580_);
  and (_06586_, _06541_, _05903_);
  or (_26886_[2], _06586_, _06585_);
  and (_06587_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  and (_06588_, _04243_, _26170_);
  or (_27169_, _06588_, _06587_);
  and (_06589_, _06529_, word_in[3]);
  not (_06590_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_06591_, _06529_, _06590_);
  nor (_06592_, _06591_, _06589_);
  nor (_06593_, _06592_, _06528_);
  and (_06595_, _06528_, word_in[11]);
  or (_06597_, _06595_, _06593_);
  and (_06599_, _06597_, _06544_);
  and (_06600_, _06527_, _06439_);
  or (_06601_, _06600_, _06599_);
  and (_06602_, _06601_, _06542_);
  and (_06604_, _06541_, word_in[27]);
  or (_26886_[3], _06604_, _06602_);
  or (_06605_, _06559_, word_in[12]);
  not (_06606_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_06607_, _06529_, _06606_);
  and (_06608_, _06529_, _06061_);
  or (_06609_, _06608_, _06607_);
  or (_06610_, _06609_, _06528_);
  and (_06611_, _06610_, _06544_);
  and (_06612_, _06611_, _06605_);
  and (_06613_, _06527_, _06461_);
  or (_06614_, _06613_, _06541_);
  or (_06615_, _06614_, _06612_);
  or (_06616_, _06542_, word_in[28]);
  and (_26886_[4], _06616_, _06615_);
  and (_06617_, _26421_, _26260_);
  not (_06618_, _06617_);
  and (_06619_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  and (_06620_, _06617_, _25886_);
  or (_02048_, _06620_, _06619_);
  not (_06621_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_06622_, _06529_, _06621_);
  and (_06623_, _06529_, _05939_);
  or (_06624_, _06623_, _06622_);
  or (_06625_, _06624_, _06528_);
  or (_06626_, _06559_, word_in[13]);
  and (_06627_, _06626_, _06625_);
  or (_06628_, _06627_, _06527_);
  or (_06630_, _06544_, _06477_);
  and (_06631_, _06630_, _06628_);
  or (_06633_, _06631_, _06541_);
  or (_06634_, _06542_, word_in[29]);
  and (_26886_[5], _06634_, _06633_);
  not (_06636_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_06637_, _06529_, _06636_);
  and (_06638_, _06529_, _05955_);
  or (_06640_, _06638_, _06637_);
  or (_06641_, _06640_, _06528_);
  or (_06642_, _06559_, word_in[14]);
  and (_06643_, _06642_, _06641_);
  or (_06644_, _06643_, _06527_);
  or (_06645_, _06544_, _06492_);
  and (_06646_, _06645_, _06542_);
  and (_06647_, _06646_, _06644_);
  and (_06649_, _06541_, _05968_);
  or (_26886_[6], _06649_, _06647_);
  and (_06650_, _06529_, word_in[7]);
  nor (_06651_, _06529_, _05031_);
  nor (_06652_, _06651_, _06650_);
  nor (_06653_, _06652_, _06528_);
  and (_06655_, _06528_, word_in[15]);
  or (_06656_, _06655_, _06653_);
  and (_06657_, _06656_, _06544_);
  and (_06659_, _06527_, _05340_);
  or (_06661_, _06659_, _06541_);
  or (_06662_, _06661_, _06657_);
  or (_06663_, _06542_, _05348_);
  and (_26886_[7], _06663_, _06662_);
  and (_06664_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_06665_, _04113_, _26242_);
  or (_02077_, _06665_, _06664_);
  and (_06666_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_06667_, _04113_, _23830_);
  or (_02080_, _06667_, _06666_);
  and (_06668_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_06670_, _04105_, _26170_);
  or (_02086_, _06670_, _06668_);
  and (_06672_, _04139_, _26185_);
  and (_06673_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or (_02094_, _06673_, _06672_);
  and (_06674_, _04139_, _23830_);
  and (_06675_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or (_02099_, _06675_, _06674_);
  and (_06676_, _04202_, _25886_);
  and (_06677_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_27187_, _06677_, _06676_);
  and (_06679_, _06376_, _05065_);
  not (_06680_, _06679_);
  and (_06681_, _06382_, _05063_);
  and (_06682_, _06681_, _05862_);
  not (_06683_, _06681_);
  and (_06684_, _06127_, _05100_);
  and (_06685_, _06131_, _05072_);
  and (_06686_, _06685_, word_in[0]);
  not (_06687_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_06689_, _06685_, _06687_);
  nor (_06690_, _06689_, _06686_);
  nor (_06691_, _06690_, _06684_);
  and (_06692_, _06684_, word_in[8]);
  or (_06693_, _06692_, _06691_);
  and (_06694_, _06693_, _06683_);
  or (_06695_, _06694_, _06682_);
  and (_06697_, _06695_, _06680_);
  and (_06698_, _06679_, word_in[24]);
  or (_26887_[0], _06698_, _06697_);
  not (_06699_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_06700_, _06685_, _06699_);
  and (_06702_, _06685_, word_in[1]);
  or (_06704_, _06702_, _06700_);
  or (_06705_, _06704_, _06684_);
  not (_06706_, _06684_);
  or (_06707_, _06706_, word_in[9]);
  and (_06708_, _06707_, _06705_);
  or (_06709_, _06708_, _06681_);
  or (_06710_, _06683_, _06415_);
  and (_06711_, _06710_, _06709_);
  or (_06712_, _06711_, _06679_);
  or (_06713_, _06680_, word_in[25]);
  and (_26887_[1], _06713_, _06712_);
  not (_06714_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_06715_, _06685_, _06714_);
  and (_06716_, _06685_, word_in[2]);
  nor (_06717_, _06716_, _06715_);
  nor (_06718_, _06717_, _06684_);
  and (_06719_, _06684_, word_in[10]);
  or (_06720_, _06719_, _06718_);
  and (_06721_, _06720_, _06683_);
  and (_06722_, _06681_, _06431_);
  or (_06724_, _06722_, _06679_);
  or (_06725_, _06724_, _06721_);
  or (_06727_, _06680_, _05903_);
  and (_26887_[2], _06727_, _06725_);
  or (_06729_, _06706_, word_in[11]);
  not (_06731_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_06732_, _06685_, _06731_);
  and (_06733_, _06685_, word_in[3]);
  or (_06734_, _06733_, _06732_);
  or (_06735_, _06734_, _06684_);
  and (_06736_, _06735_, _06683_);
  and (_06738_, _06736_, _06729_);
  and (_06739_, _06681_, _06439_);
  or (_06740_, _06739_, _06679_);
  or (_06741_, _06740_, _06738_);
  or (_06743_, _06680_, word_in[27]);
  and (_26887_[3], _06743_, _06741_);
  and (_06745_, _06685_, word_in[4]);
  not (_06746_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_06747_, _06685_, _06746_);
  nor (_06748_, _06747_, _06745_);
  nor (_06749_, _06748_, _06684_);
  and (_06750_, _06684_, word_in[12]);
  or (_06751_, _06750_, _06749_);
  and (_06753_, _06751_, _06683_);
  and (_06755_, _06681_, _06461_);
  or (_06757_, _06755_, _06753_);
  and (_06758_, _06757_, _06680_);
  and (_06759_, _06679_, word_in[28]);
  or (_26887_[4], _06759_, _06758_);
  and (_06760_, _04202_, _26185_);
  and (_06761_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_02115_, _06761_, _06760_);
  not (_06763_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_06764_, _06685_, _06763_);
  and (_06766_, _06685_, word_in[5]);
  or (_06767_, _06766_, _06764_);
  or (_06768_, _06767_, _06684_);
  or (_06770_, _06706_, word_in[13]);
  and (_06771_, _06770_, _06768_);
  or (_06772_, _06771_, _06681_);
  or (_06773_, _06683_, _06477_);
  and (_06774_, _06773_, _06680_);
  and (_06775_, _06774_, _06772_);
  and (_06777_, _06679_, _05950_);
  or (_26887_[5], _06777_, _06775_);
  not (_06778_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_06780_, _06685_, _06778_);
  and (_06781_, _06685_, word_in[6]);
  nor (_06782_, _06781_, _06780_);
  nor (_06783_, _06782_, _06684_);
  and (_06784_, _06684_, word_in[14]);
  or (_06785_, _06784_, _06783_);
  and (_06786_, _06785_, _06683_);
  and (_06787_, _06681_, _06492_);
  or (_06789_, _06787_, _06679_);
  or (_06791_, _06789_, _06786_);
  or (_06792_, _06680_, _05968_);
  and (_26887_[6], _06792_, _06791_);
  and (_06793_, _06681_, _05340_);
  nor (_06794_, _06685_, _05168_);
  and (_06796_, _06685_, word_in[7]);
  nor (_06797_, _06796_, _06794_);
  nor (_06798_, _06797_, _06684_);
  and (_06799_, _06684_, word_in[15]);
  or (_06800_, _06799_, _06798_);
  and (_06802_, _06800_, _06683_);
  or (_06803_, _06802_, _06793_);
  and (_06804_, _06803_, _06680_);
  and (_06805_, _06679_, word_in[31]);
  or (_26887_[7], _06805_, _06804_);
  and (_06806_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  and (_06808_, _26541_, _26170_);
  or (_02133_, _06808_, _06806_);
  and (_06809_, _04092_, _26170_);
  and (_06810_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or (_27190_, _06810_, _06809_);
  and (_06811_, _04198_, _25886_);
  and (_06812_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or (_02145_, _06812_, _06811_);
  and (_06813_, _04198_, _23768_);
  and (_06814_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or (_02150_, _06814_, _06813_);
  and (_06815_, _06376_, _05063_);
  not (_06816_, _06815_);
  and (_06817_, _06382_, _05093_);
  and (_06818_, _06817_, _05862_);
  not (_06819_, _06817_);
  and (_06821_, _05321_, _05100_);
  not (_06822_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_06823_, _06389_, _05324_);
  nor (_06824_, _06823_, _06822_);
  and (_06826_, _06823_, word_in[0]);
  nor (_06828_, _06826_, _06824_);
  nor (_06829_, _06828_, _06821_);
  and (_06830_, _06821_, word_in[8]);
  or (_06831_, _06830_, _06829_);
  and (_06832_, _06831_, _06819_);
  or (_06833_, _06832_, _06818_);
  and (_06834_, _06833_, _06816_);
  and (_06835_, _06815_, word_in[24]);
  or (_26888_[0], _06835_, _06834_);
  and (_06836_, _04026_, _26283_);
  and (_06837_, _06836_, _25927_);
  not (_06838_, _06836_);
  and (_06839_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or (_02174_, _06839_, _06837_);
  not (_06840_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_06841_, _06823_, _06840_);
  and (_06842_, _06823_, _05875_);
  or (_06843_, _06842_, _06841_);
  or (_06844_, _06843_, _06821_);
  not (_06845_, _06821_);
  or (_06847_, _06845_, word_in[9]);
  and (_06848_, _06847_, _06844_);
  or (_06849_, _06848_, _06817_);
  or (_06850_, _06819_, _06415_);
  and (_06852_, _06850_, _06816_);
  and (_06853_, _06852_, _06849_);
  and (_06854_, _06815_, _05870_);
  or (_26888_[1], _06854_, _06853_);
  or (_06855_, _06819_, _06431_);
  not (_06857_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_06859_, _06823_, _06857_);
  and (_06860_, _06823_, _05892_);
  or (_06861_, _06860_, _06859_);
  or (_06862_, _06861_, _06821_);
  or (_06863_, _06845_, word_in[10]);
  and (_06864_, _06863_, _06862_);
  or (_06865_, _06864_, _06817_);
  and (_06866_, _06865_, _06855_);
  or (_06867_, _06866_, _06815_);
  or (_06868_, _06816_, word_in[26]);
  and (_26888_[2], _06868_, _06867_);
  not (_06869_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_06871_, _06823_, _06869_);
  and (_06872_, _06823_, word_in[3]);
  nor (_06873_, _06872_, _06871_);
  nor (_06874_, _06873_, _06821_);
  and (_06875_, _06821_, word_in[11]);
  or (_06877_, _06875_, _06874_);
  and (_06878_, _06877_, _06819_);
  and (_06879_, _06817_, _06439_);
  or (_06881_, _06879_, _06878_);
  and (_06882_, _06881_, _06816_);
  and (_06884_, _06815_, word_in[27]);
  or (_26888_[3], _06884_, _06882_);
  not (_06885_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_06886_, _06823_, _06885_);
  and (_06888_, _06823_, word_in[4]);
  nor (_06889_, _06888_, _06886_);
  nor (_06890_, _06889_, _06821_);
  and (_06892_, _06821_, word_in[12]);
  or (_06894_, _06892_, _06890_);
  and (_06895_, _06894_, _06819_);
  and (_06896_, _06817_, _06461_);
  or (_06898_, _06896_, _06895_);
  and (_06899_, _06898_, _06816_);
  and (_06901_, _06815_, word_in[28]);
  or (_26888_[4], _06901_, _06899_);
  and (_06902_, _06817_, _06477_);
  not (_06903_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_06905_, _06823_, _06903_);
  and (_06906_, _06823_, word_in[5]);
  nor (_06907_, _06906_, _06905_);
  nor (_06908_, _06907_, _06821_);
  and (_06909_, _06821_, word_in[13]);
  or (_06911_, _06909_, _06908_);
  and (_06912_, _06911_, _06819_);
  or (_06913_, _06912_, _06902_);
  and (_06915_, _06913_, _06816_);
  and (_06916_, _06815_, word_in[29]);
  or (_26888_[5], _06916_, _06915_);
  and (_06917_, _06817_, _06492_);
  not (_06918_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_06919_, _06823_, _06918_);
  and (_06920_, _06823_, word_in[6]);
  nor (_06921_, _06920_, _06919_);
  nor (_06922_, _06921_, _06821_);
  and (_06923_, _06821_, word_in[14]);
  or (_06924_, _06923_, _06922_);
  and (_06925_, _06924_, _06819_);
  or (_06926_, _06925_, _06917_);
  and (_06927_, _06926_, _06816_);
  and (_06928_, _06815_, word_in[30]);
  or (_26888_[6], _06928_, _06927_);
  nor (_06929_, _06823_, _05045_);
  and (_06930_, _06823_, _05971_);
  or (_06931_, _06930_, _06929_);
  or (_06932_, _06931_, _06821_);
  or (_06933_, _06845_, word_in[15]);
  and (_06934_, _06933_, _06932_);
  or (_06936_, _06934_, _06817_);
  or (_06937_, _06819_, _05340_);
  and (_06938_, _06937_, _06936_);
  or (_06940_, _06938_, _06815_);
  or (_06941_, _06816_, word_in[31]);
  and (_26888_[7], _06941_, _06940_);
  and (_06942_, _04194_, _26242_);
  and (_06943_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_02194_, _06943_, _06942_);
  nor (_26929_[7], _24205_, rst);
  and (_06946_, _04026_, _26421_);
  and (_06947_, _06946_, _26185_);
  not (_06948_, _06946_);
  and (_06949_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or (_27206_, _06949_, _06947_);
  and (_06951_, _05336_, _05251_);
  and (_06953_, _06951_, _05093_);
  and (_06954_, _05315_, _05472_);
  and (_06955_, _05320_, _05073_);
  not (_06956_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_06957_, _05325_, _04984_);
  and (_06958_, _06957_, _05844_);
  nor (_06959_, _06958_, _06956_);
  and (_06961_, _06958_, word_in[0]);
  or (_06962_, _06961_, _06959_);
  or (_06964_, _06962_, _06955_);
  not (_06965_, _06955_);
  or (_06967_, _06965_, word_in[8]);
  and (_06968_, _06967_, _06964_);
  or (_06970_, _06968_, _06954_);
  not (_06971_, _06954_);
  or (_06973_, _06971_, word_in[16]);
  and (_06974_, _06973_, _06970_);
  or (_06976_, _06974_, _06953_);
  not (_06978_, _06953_);
  or (_06979_, _06978_, word_in[24]);
  and (_26889_[0], _06979_, _06976_);
  not (_06980_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_06982_, _06958_, _06980_);
  and (_06983_, _06958_, word_in[1]);
  or (_06984_, _06983_, _06982_);
  and (_06985_, _06984_, _06965_);
  and (_06986_, _06955_, word_in[9]);
  or (_06987_, _06986_, _06985_);
  and (_06988_, _06987_, _06971_);
  and (_06989_, _06954_, word_in[17]);
  or (_06990_, _06989_, _06988_);
  and (_06991_, _06990_, _06978_);
  and (_06993_, _06953_, word_in[25]);
  or (_26889_[1], _06993_, _06991_);
  and (_06995_, _06954_, word_in[18]);
  not (_06997_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_06999_, _06958_, _06997_);
  and (_07001_, _06958_, word_in[2]);
  or (_07003_, _07001_, _06999_);
  and (_07004_, _07003_, _06965_);
  and (_07005_, _06955_, word_in[10]);
  or (_07006_, _07005_, _07004_);
  and (_07008_, _07006_, _06971_);
  or (_07009_, _07008_, _06995_);
  and (_07010_, _07009_, _06978_);
  and (_07012_, _06953_, word_in[26]);
  or (_26889_[2], _07012_, _07010_);
  and (_07014_, _04035_, _26085_);
  and (_07015_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_02241_, _07015_, _07014_);
  not (_07016_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_07017_, _06958_, _07016_);
  and (_07019_, _06958_, word_in[3]);
  or (_07021_, _07019_, _07017_);
  and (_07023_, _07021_, _06965_);
  and (_07024_, _06955_, word_in[11]);
  or (_07025_, _07024_, _07023_);
  and (_07026_, _07025_, _06971_);
  and (_07027_, _06954_, word_in[19]);
  or (_07028_, _07027_, _07026_);
  and (_07029_, _07028_, _06978_);
  and (_07030_, _06953_, word_in[27]);
  or (_26889_[3], _07030_, _07029_);
  and (_07031_, _06954_, word_in[20]);
  not (_07032_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_07033_, _06958_, _07032_);
  and (_07034_, _06958_, word_in[4]);
  or (_07035_, _07034_, _07033_);
  and (_07036_, _07035_, _06965_);
  and (_07037_, _06955_, word_in[12]);
  or (_07038_, _07037_, _07036_);
  and (_07039_, _07038_, _06971_);
  or (_07041_, _07039_, _07031_);
  and (_07043_, _07041_, _06978_);
  and (_07044_, _06953_, word_in[28]);
  or (_26889_[4], _07044_, _07043_);
  and (_07046_, _04035_, _25886_);
  and (_07048_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_02245_, _07048_, _07046_);
  not (_07051_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_07053_, _06958_, _07051_);
  and (_07054_, _06958_, word_in[5]);
  or (_07056_, _07054_, _07053_);
  and (_07058_, _07056_, _06965_);
  and (_07060_, _06955_, word_in[13]);
  or (_07061_, _07060_, _07058_);
  and (_07062_, _07061_, _06971_);
  and (_07064_, _06954_, word_in[21]);
  or (_07066_, _07064_, _07062_);
  and (_07068_, _07066_, _06978_);
  and (_07070_, _06953_, word_in[29]);
  or (_26889_[5], _07070_, _07068_);
  not (_07073_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_07074_, _06958_, _07073_);
  and (_07075_, _06958_, word_in[6]);
  or (_07076_, _07075_, _07074_);
  and (_07077_, _07076_, _06965_);
  and (_07079_, _06955_, word_in[14]);
  or (_07080_, _07079_, _07077_);
  and (_07081_, _07080_, _06971_);
  and (_07082_, _06954_, word_in[22]);
  or (_07083_, _07082_, _07081_);
  and (_07084_, _07083_, _06978_);
  and (_07085_, _06953_, word_in[30]);
  or (_26889_[6], _07085_, _07084_);
  and (_07087_, _06954_, word_in[23]);
  nor (_07088_, _06958_, _05130_);
  and (_07089_, _06958_, word_in[7]);
  or (_07091_, _07089_, _07088_);
  and (_07092_, _07091_, _06965_);
  and (_07094_, _06955_, word_in[15]);
  or (_07095_, _07094_, _07092_);
  and (_07096_, _07095_, _06971_);
  or (_07097_, _07096_, _07087_);
  and (_07098_, _07097_, _06978_);
  and (_07099_, _06953_, word_in[31]);
  or (_26889_[7], _07099_, _07098_);
  and (_07102_, _04181_, _25886_);
  and (_07103_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or (_02266_, _07103_, _07102_);
  and (_07104_, _04026_, _26202_);
  and (_07105_, _07104_, _25927_);
  not (_07106_, _07104_);
  and (_07107_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_02280_, _07107_, _07105_);
  and (_07108_, _06951_, _05109_);
  not (_07109_, _07108_);
  and (_07110_, _05993_, _05186_);
  and (_07111_, _07110_, _05862_);
  not (_07112_, _07110_);
  and (_07113_, _05998_, _05076_);
  and (_07114_, _06957_, _06004_);
  and (_07115_, _07114_, word_in[0]);
  not (_07116_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_07117_, _07114_, _07116_);
  nor (_07118_, _07117_, _07115_);
  nor (_07119_, _07118_, _07113_);
  and (_07120_, _07113_, word_in[8]);
  or (_07121_, _07120_, _07119_);
  and (_07122_, _07121_, _07112_);
  or (_07123_, _07122_, _07111_);
  and (_07124_, _07123_, _07109_);
  and (_07125_, _07108_, word_in[24]);
  or (_26890_[0], _07125_, _07124_);
  not (_07126_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_07127_, _07114_, _07126_);
  and (_07128_, _07114_, _05875_);
  or (_07129_, _07128_, _07127_);
  or (_07130_, _07129_, _07113_);
  not (_07131_, _07113_);
  or (_07132_, _07131_, word_in[9]);
  and (_07133_, _07132_, _07130_);
  or (_07134_, _07133_, _07110_);
  or (_07136_, _07112_, _06415_);
  and (_07137_, _07136_, _07109_);
  and (_07138_, _07137_, _07134_);
  and (_07139_, _07108_, word_in[25]);
  or (_26890_[1], _07139_, _07138_);
  and (_07141_, _07110_, _06431_);
  and (_07142_, _07114_, word_in[2]);
  not (_07143_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_07144_, _07114_, _07143_);
  nor (_07145_, _07144_, _07142_);
  nor (_07146_, _07145_, _07113_);
  and (_07147_, _07113_, word_in[10]);
  or (_07148_, _07147_, _07146_);
  and (_07149_, _07148_, _07112_);
  or (_07150_, _07149_, _07141_);
  and (_07152_, _07150_, _07109_);
  and (_07154_, _07108_, word_in[26]);
  or (_26890_[2], _07154_, _07152_);
  and (_07155_, _07110_, _06439_);
  and (_07157_, _07114_, word_in[3]);
  not (_07158_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_07159_, _07114_, _07158_);
  nor (_07160_, _07159_, _07157_);
  nor (_07161_, _07160_, _07113_);
  and (_07162_, _07113_, word_in[11]);
  or (_07164_, _07162_, _07161_);
  and (_07165_, _07164_, _07112_);
  or (_07166_, _07165_, _07155_);
  and (_07168_, _07166_, _07109_);
  and (_07171_, _07108_, word_in[27]);
  or (_26890_[3], _07171_, _07168_);
  not (_07172_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_07173_, _07114_, _07172_);
  and (_07174_, _07114_, _06061_);
  or (_07175_, _07174_, _07173_);
  or (_07176_, _07175_, _07113_);
  or (_07178_, _07131_, word_in[12]);
  and (_07180_, _07178_, _07176_);
  or (_07181_, _07180_, _07110_);
  or (_07182_, _07112_, _06461_);
  and (_07183_, _07182_, _07109_);
  and (_07184_, _07183_, _07181_);
  and (_07185_, _07108_, word_in[28]);
  or (_26890_[4], _07185_, _07184_);
  and (_07186_, _07114_, word_in[5]);
  not (_07188_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_07190_, _07114_, _07188_);
  nor (_07191_, _07190_, _07186_);
  nor (_07192_, _07191_, _07113_);
  and (_07193_, _07113_, word_in[13]);
  or (_07194_, _07193_, _07192_);
  and (_07195_, _07194_, _07112_);
  and (_07196_, _07110_, _06477_);
  or (_07197_, _07196_, _07108_);
  or (_07199_, _07197_, _07195_);
  or (_07200_, _07109_, word_in[29]);
  and (_26890_[5], _07200_, _07199_);
  and (_07201_, _07110_, _06492_);
  and (_07202_, _07114_, word_in[6]);
  not (_07204_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_07205_, _07114_, _07204_);
  nor (_07206_, _07205_, _07202_);
  nor (_07207_, _07206_, _07113_);
  and (_07208_, _07113_, word_in[14]);
  or (_07209_, _07208_, _07207_);
  and (_07210_, _07209_, _07112_);
  or (_07211_, _07210_, _07201_);
  and (_07212_, _07211_, _07109_);
  and (_07213_, _07108_, word_in[30]);
  or (_26890_[6], _07213_, _07212_);
  not (_07215_, rxd_i);
  and (_07216_, _02394_, _02274_);
  and (_07217_, _02383_, _07216_);
  nand (_07218_, _07217_, _07215_);
  or (_07219_, _07217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_07220_, _07219_, _23049_);
  and (_02305_, _07220_, _07218_);
  and (_07221_, _07110_, _05340_);
  and (_07222_, _07114_, word_in[7]);
  nor (_07223_, _07114_, _05023_);
  nor (_07224_, _07223_, _07222_);
  nor (_07225_, _07224_, _07113_);
  and (_07226_, _07113_, word_in[15]);
  or (_07227_, _07226_, _07225_);
  and (_07228_, _07227_, _07112_);
  or (_07229_, _07228_, _07221_);
  and (_07230_, _07229_, _07109_);
  and (_07231_, _07108_, word_in[31]);
  or (_26890_[7], _07231_, _07230_);
  and (_07232_, _06121_, _05186_);
  not (_07233_, _07232_);
  and (_07234_, _06127_, _05076_);
  and (_07235_, _06131_, _04984_);
  and (_07236_, _07235_, word_in[0]);
  not (_07238_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_07239_, _07235_, _07238_);
  nor (_07241_, _07239_, _07236_);
  nor (_07242_, _07241_, _07234_);
  and (_07243_, _07234_, word_in[8]);
  or (_07245_, _07243_, _07242_);
  and (_07246_, _07245_, _07233_);
  and (_07248_, _06951_, _05065_);
  and (_07249_, _07232_, _05862_);
  or (_07250_, _07249_, _07248_);
  or (_07251_, _07250_, _07246_);
  not (_07252_, _07248_);
  or (_07253_, _07252_, word_in[24]);
  and (_26876_[0], _07253_, _07251_);
  and (_07256_, _07232_, _06415_);
  and (_07258_, _07235_, word_in[1]);
  not (_07259_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_07260_, _07235_, _07259_);
  nor (_07261_, _07260_, _07258_);
  nor (_07262_, _07261_, _07234_);
  and (_07263_, _07234_, word_in[9]);
  or (_07264_, _07263_, _07262_);
  and (_07265_, _07264_, _07233_);
  or (_07266_, _07265_, _07256_);
  and (_07268_, _07266_, _07252_);
  and (_07270_, _07248_, word_in[25]);
  or (_26876_[1], _07270_, _07268_);
  not (_07271_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_07273_, _07235_, _07271_);
  and (_07274_, _07235_, word_in[2]);
  or (_07276_, _07274_, _07273_);
  or (_07278_, _07276_, _07234_);
  not (_07280_, _07234_);
  or (_07281_, _07280_, word_in[10]);
  and (_07283_, _07281_, _07278_);
  or (_07285_, _07283_, _07232_);
  or (_07286_, _07233_, _06431_);
  and (_07287_, _07286_, _07285_);
  or (_07288_, _07287_, _07248_);
  or (_07289_, _07252_, word_in[26]);
  and (_26876_[2], _07289_, _07288_);
  not (_07291_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_07292_, _07235_, _07291_);
  and (_07293_, _07235_, word_in[3]);
  or (_07294_, _07293_, _07292_);
  or (_07295_, _07294_, _07234_);
  or (_07297_, _07280_, word_in[11]);
  and (_07298_, _07297_, _07295_);
  or (_07299_, _07298_, _07232_);
  or (_07300_, _07233_, _06439_);
  and (_07301_, _07300_, _07252_);
  and (_07302_, _07301_, _07299_);
  and (_07303_, _07248_, word_in[27]);
  or (_26876_[3], _07303_, _07302_);
  not (_07305_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_07306_, _07235_, _07305_);
  and (_07308_, _07235_, word_in[4]);
  or (_07309_, _07308_, _07306_);
  or (_07310_, _07309_, _07234_);
  or (_07311_, _07280_, word_in[12]);
  and (_07312_, _07311_, _07310_);
  or (_07313_, _07312_, _07232_);
  or (_07315_, _07233_, _06461_);
  and (_07316_, _07315_, _07252_);
  and (_07317_, _07316_, _07313_);
  and (_07320_, _07248_, word_in[28]);
  or (_26876_[4], _07320_, _07317_);
  not (_07321_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_07322_, _07235_, _07321_);
  and (_07323_, _07235_, word_in[5]);
  or (_07324_, _07323_, _07322_);
  or (_07325_, _07324_, _07234_);
  or (_07326_, _07280_, word_in[13]);
  and (_07328_, _07326_, _07325_);
  or (_07329_, _07328_, _07232_);
  or (_07330_, _07233_, _06477_);
  and (_07332_, _07330_, _07252_);
  and (_07333_, _07332_, _07329_);
  and (_07335_, _07248_, word_in[29]);
  or (_26876_[5], _07335_, _07333_);
  and (_07337_, _07232_, _06492_);
  and (_07338_, _07235_, word_in[6]);
  not (_07339_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_07340_, _07235_, _07339_);
  nor (_07341_, _07340_, _07338_);
  nor (_07342_, _07341_, _07234_);
  and (_07343_, _07234_, word_in[14]);
  or (_07344_, _07343_, _07342_);
  and (_07345_, _07344_, _07233_);
  or (_07346_, _07345_, _07337_);
  and (_07347_, _07346_, _07252_);
  and (_07348_, _07248_, word_in[30]);
  or (_26876_[6], _07348_, _07347_);
  or (_07349_, _04283_, rxd_i);
  nand (_07350_, _07349_, _02283_);
  or (_07351_, _02284_, _02271_);
  and (_07352_, _07351_, _07350_);
  or (_07353_, _02288_, _02282_);
  or (_07354_, _07353_, _02272_);
  or (_07355_, _07354_, _07352_);
  and (_02345_, _07355_, _01634_);
  or (_07356_, _07233_, _05340_);
  nor (_07358_, _07235_, _05125_);
  and (_07360_, _07235_, word_in[7]);
  or (_07361_, _07360_, _07358_);
  or (_07362_, _07361_, _07234_);
  or (_07363_, _07280_, word_in[15]);
  and (_07365_, _07363_, _07362_);
  or (_07366_, _07365_, _07232_);
  and (_07368_, _07366_, _07356_);
  or (_07370_, _07368_, _07248_);
  or (_07371_, _07252_, word_in[31]);
  and (_26876_[7], _07371_, _07370_);
  or (_07372_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_07373_, _07372_, _23049_);
  nand (_07375_, _02031_, _25417_);
  and (_02378_, _07375_, _07373_);
  not (_07376_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_07377_, _02058_, _07376_);
  or (_07378_, _07377_, _04232_);
  and (_07379_, _07378_, _02055_);
  nand (_07380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_07381_, _07380_, _02054_);
  nor (_07383_, _07381_, _07379_);
  nor (_07384_, _07383_, _02052_);
  or (_07385_, _07384_, _02126_);
  nand (_07386_, _07385_, _23049_);
  nor (_02381_, _07386_, _02045_);
  and (_07387_, _05316_, _05186_);
  not (_07388_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_07389_, _06957_, _05324_);
  nor (_07390_, _07389_, _07388_);
  and (_07391_, _07389_, _06002_);
  or (_07393_, _07391_, _07390_);
  and (_07394_, _05321_, _05076_);
  or (_07395_, _07394_, _07393_);
  not (_07396_, _07394_);
  or (_07398_, _07396_, word_in[8]);
  and (_07399_, _07398_, _07395_);
  or (_07400_, _07399_, _07387_);
  and (_07401_, _06951_, _05063_);
  not (_07402_, _07401_);
  not (_07403_, _07387_);
  or (_07404_, _07403_, _05862_);
  and (_07405_, _07404_, _07402_);
  and (_07406_, _07405_, _07400_);
  and (_07407_, _05336_, word_in[24]);
  and (_07408_, _07401_, _07407_);
  or (_26877_[0], _07408_, _07406_);
  and (_07409_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  and (_07411_, _06369_, _26085_);
  or (_02393_, _07411_, _07409_);
  and (_07412_, _07389_, word_in[1]);
  not (_07413_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_07415_, _07389_, _07413_);
  nor (_07417_, _07415_, _07412_);
  nor (_07418_, _07417_, _07394_);
  and (_07419_, _07394_, word_in[9]);
  or (_07420_, _07419_, _07418_);
  and (_07421_, _07420_, _07403_);
  and (_07423_, _07387_, _06415_);
  or (_07424_, _07423_, _07401_);
  or (_07425_, _07424_, _07421_);
  or (_07426_, _07402_, _05870_);
  and (_26877_[1], _07426_, _07425_);
  and (_07428_, _07389_, word_in[2]);
  not (_07430_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_07432_, _07389_, _07430_);
  nor (_07434_, _07432_, _07428_);
  nor (_07435_, _07434_, _07394_);
  and (_07436_, _07394_, word_in[10]);
  or (_07437_, _07436_, _07435_);
  and (_07439_, _07437_, _07403_);
  and (_07440_, _07387_, _06431_);
  or (_07441_, _07440_, _07401_);
  or (_07442_, _07441_, _07439_);
  or (_07443_, _07402_, _05903_);
  and (_26877_[2], _07443_, _07442_);
  not (_07444_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_07445_, _07389_, _07444_);
  and (_07446_, _07389_, _05907_);
  or (_07447_, _07446_, _07445_);
  or (_07448_, _07447_, _07394_);
  or (_07449_, _07396_, word_in[11]);
  and (_07450_, _07449_, _07448_);
  or (_07451_, _07450_, _07387_);
  or (_07452_, _07403_, _06439_);
  and (_07453_, _07452_, _07402_);
  and (_07454_, _07453_, _07451_);
  and (_07455_, _07401_, _05919_);
  or (_26877_[3], _07455_, _07454_);
  and (_07456_, _07389_, word_in[4]);
  not (_07457_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_07459_, _07389_, _07457_);
  nor (_07460_, _07459_, _07456_);
  nor (_07461_, _07460_, _07394_);
  and (_07462_, _07394_, word_in[12]);
  or (_07464_, _07462_, _07461_);
  and (_07466_, _07464_, _07403_);
  and (_07467_, _07387_, _06461_);
  or (_07468_, _07467_, _07401_);
  or (_07470_, _07468_, _07466_);
  or (_07471_, _07402_, _06465_);
  and (_26877_[4], _07471_, _07470_);
  and (_07473_, _07389_, word_in[5]);
  not (_07475_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_07476_, _07389_, _07475_);
  nor (_07478_, _07476_, _07473_);
  nor (_07479_, _07478_, _07394_);
  and (_07481_, _07394_, word_in[13]);
  or (_07482_, _07481_, _07479_);
  and (_07483_, _07482_, _07403_);
  and (_07484_, _07387_, _06477_);
  or (_07485_, _07484_, _07401_);
  or (_07486_, _07485_, _07483_);
  or (_07488_, _07402_, _05950_);
  and (_26877_[5], _07488_, _07486_);
  and (_07490_, _07387_, _06492_);
  and (_07491_, _07389_, word_in[6]);
  not (_07492_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_07494_, _07389_, _07492_);
  nor (_07495_, _07494_, _07491_);
  nor (_07496_, _07495_, _07394_);
  and (_07498_, _07394_, word_in[14]);
  or (_07500_, _07498_, _07496_);
  and (_07501_, _07500_, _07403_);
  or (_07503_, _07501_, _07490_);
  and (_07505_, _07503_, _07402_);
  and (_07506_, _07401_, word_in[30]);
  or (_26877_[6], _07506_, _07505_);
  nor (_07508_, _07389_, _05011_);
  and (_07509_, _07389_, _05971_);
  or (_07510_, _07509_, _07508_);
  or (_07511_, _07510_, _07394_);
  or (_07512_, _07396_, word_in[15]);
  and (_07515_, _07512_, _07511_);
  or (_07517_, _07515_, _07387_);
  or (_07518_, _07403_, _05340_);
  and (_07520_, _07518_, _07402_);
  and (_07522_, _07520_, _07517_);
  and (_07523_, _07401_, _05348_);
  or (_26877_[7], _07523_, _07522_);
  and (_07525_, _05771_, _26242_);
  and (_07526_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  or (_02439_, _07526_, _07525_);
  and (_07527_, _06380_, _05185_);
  and (_07528_, _07527_, _05109_);
  not (_07529_, _07528_);
  and (_07531_, _05320_, _05719_);
  not (_07533_, _07531_);
  not (_07534_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_07536_, _05844_, _05326_);
  nor (_07537_, _07536_, _07534_);
  and (_07538_, _07536_, word_in[0]);
  or (_07539_, _07538_, _07537_);
  and (_07540_, _07539_, _07533_);
  and (_07541_, _07531_, word_in[8]);
  or (_07542_, _07541_, _07540_);
  and (_07543_, _07542_, _07529_);
  and (_07544_, _05337_, _05093_);
  and (_07545_, _07528_, _05862_);
  or (_07546_, _07545_, _07544_);
  or (_07548_, _07546_, _07543_);
  not (_07550_, _07544_);
  or (_07552_, _07550_, _07407_);
  and (_26878_[0], _07552_, _07548_);
  and (_07553_, _07528_, _06415_);
  not (_07555_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_07556_, _07536_, _07555_);
  and (_07557_, _07536_, word_in[1]);
  or (_07558_, _07557_, _07556_);
  and (_07559_, _07558_, _07533_);
  and (_07560_, _07531_, word_in[9]);
  or (_07561_, _07560_, _07559_);
  and (_07562_, _07561_, _07529_);
  or (_07563_, _07562_, _07553_);
  and (_07564_, _07563_, _07550_);
  and (_07565_, _07544_, _05870_);
  or (_26878_[1], _07565_, _07564_);
  and (_07566_, _07528_, _06431_);
  not (_07567_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_07568_, _07536_, _07567_);
  and (_07569_, _07536_, word_in[2]);
  or (_07570_, _07569_, _07568_);
  and (_07571_, _07570_, _07533_);
  and (_07572_, _07531_, word_in[10]);
  or (_07573_, _07572_, _07571_);
  and (_07574_, _07573_, _07529_);
  or (_07575_, _07574_, _07566_);
  and (_07576_, _07575_, _07550_);
  and (_07577_, _07544_, _05903_);
  or (_26878_[2], _07577_, _07576_);
  not (_07578_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_07579_, _07536_, _07578_);
  and (_07580_, _07536_, word_in[3]);
  or (_07582_, _07580_, _07579_);
  and (_07584_, _07582_, _07533_);
  and (_07585_, _07531_, word_in[11]);
  or (_07586_, _07585_, _07584_);
  and (_07587_, _07586_, _07529_);
  and (_07588_, _07528_, _06439_);
  or (_07589_, _07588_, _07587_);
  and (_07590_, _07589_, _07550_);
  and (_07591_, _07544_, _05919_);
  or (_26878_[3], _07591_, _07590_);
  and (_07592_, _07528_, _06461_);
  not (_07593_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_07594_, _07536_, _07593_);
  and (_07595_, _07536_, word_in[4]);
  or (_07596_, _07595_, _07594_);
  and (_07598_, _07596_, _07533_);
  and (_07599_, _07531_, word_in[12]);
  or (_07601_, _07599_, _07598_);
  and (_07603_, _07601_, _07529_);
  or (_07604_, _07603_, _07592_);
  and (_07605_, _07604_, _07550_);
  and (_07606_, _07544_, _06465_);
  or (_26878_[4], _07606_, _07605_);
  and (_07607_, _07528_, _06477_);
  not (_07608_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_07609_, _07536_, _07608_);
  and (_07610_, _07536_, word_in[5]);
  or (_07611_, _07610_, _07609_);
  and (_07612_, _07611_, _07533_);
  and (_07613_, _07531_, word_in[13]);
  or (_07614_, _07613_, _07612_);
  and (_07615_, _07614_, _07529_);
  or (_07616_, _07615_, _07607_);
  and (_07617_, _07616_, _07550_);
  and (_07618_, _07544_, _05950_);
  or (_26878_[5], _07618_, _07617_);
  and (_07619_, _07528_, _06492_);
  not (_07620_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_07621_, _07536_, _07620_);
  and (_07622_, _07536_, word_in[6]);
  or (_07623_, _07622_, _07621_);
  and (_07624_, _07623_, _07533_);
  and (_07625_, _07531_, word_in[14]);
  or (_07626_, _07625_, _07624_);
  and (_07627_, _07626_, _07529_);
  or (_07628_, _07627_, _07619_);
  and (_07629_, _07628_, _07550_);
  and (_07630_, _07544_, _05968_);
  or (_26878_[6], _07630_, _07629_);
  and (_07631_, _07528_, _05340_);
  nor (_07633_, _07536_, _05143_);
  and (_07634_, _07536_, word_in[7]);
  or (_07635_, _07634_, _07633_);
  and (_07636_, _07635_, _07533_);
  and (_07637_, _07531_, word_in[15]);
  or (_07638_, _07637_, _07636_);
  and (_07639_, _07638_, _07529_);
  or (_07640_, _07639_, _07631_);
  and (_07641_, _07640_, _07550_);
  and (_07642_, _07544_, _05348_);
  or (_26878_[7], _07642_, _07641_);
  and (_07643_, _05799_, _25886_);
  and (_07644_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_26977_, _07644_, _07643_);
  and (_07645_, _04157_, _26340_);
  and (_07646_, _07645_, _25927_);
  not (_07647_, _07645_);
  and (_07648_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_02491_, _07648_, _07646_);
  and (_07649_, _05337_, _05109_);
  and (_07650_, _07527_, _05065_);
  not (_07651_, _07650_);
  or (_07652_, _07651_, _05862_);
  and (_07653_, _05998_, _05095_);
  not (_07654_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_07655_, _06004_, _05326_);
  nor (_07656_, _07655_, _07654_);
  and (_07657_, _07655_, word_in[0]);
  or (_07658_, _07657_, _07656_);
  or (_07659_, _07658_, _07653_);
  not (_07660_, _07653_);
  or (_07661_, _07660_, word_in[8]);
  and (_07662_, _07661_, _07659_);
  or (_07663_, _07662_, _07650_);
  and (_07664_, _07663_, _07652_);
  or (_07665_, _07664_, _07649_);
  not (_07666_, _07649_);
  or (_07667_, _07666_, _07407_);
  and (_26879_[0], _07667_, _07665_);
  not (_07668_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_07669_, _07655_, _07668_);
  and (_07670_, _07655_, word_in[1]);
  or (_07671_, _07670_, _07669_);
  or (_07672_, _07671_, _07653_);
  or (_07673_, _07660_, word_in[9]);
  and (_07674_, _07673_, _07672_);
  or (_07675_, _07674_, _07650_);
  or (_07676_, _07651_, _06415_);
  and (_07677_, _07676_, _07675_);
  or (_07678_, _07677_, _07649_);
  or (_07679_, _07666_, _05870_);
  and (_26879_[1], _07679_, _07678_);
  and (_07680_, _07650_, _06431_);
  not (_07681_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_07682_, _07655_, _07681_);
  and (_07683_, _07655_, word_in[2]);
  nor (_07684_, _07683_, _07682_);
  nor (_07685_, _07684_, _07653_);
  and (_07686_, _07653_, word_in[10]);
  or (_07687_, _07686_, _07685_);
  and (_07689_, _07687_, _07651_);
  or (_07690_, _07689_, _07680_);
  and (_07691_, _07690_, _07666_);
  and (_07692_, _07649_, _05903_);
  or (_26879_[2], _07692_, _07691_);
  not (_07693_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_07694_, _07655_, _07693_);
  and (_07695_, _07655_, word_in[3]);
  or (_07696_, _07695_, _07694_);
  or (_07697_, _07696_, _07653_);
  or (_07698_, _07660_, word_in[11]);
  and (_07699_, _07698_, _07697_);
  or (_07700_, _07699_, _07650_);
  or (_07701_, _07651_, _06439_);
  and (_07702_, _07701_, _07700_);
  or (_07703_, _07702_, _07649_);
  or (_07704_, _07666_, _05919_);
  and (_26879_[3], _07704_, _07703_);
  not (_07705_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_07706_, _07655_, _07705_);
  and (_07708_, _07655_, word_in[4]);
  or (_07709_, _07708_, _07706_);
  or (_07710_, _07709_, _07653_);
  or (_07711_, _07660_, word_in[12]);
  and (_07712_, _07711_, _07710_);
  or (_07713_, _07712_, _07650_);
  or (_07714_, _07651_, _06461_);
  and (_07715_, _07714_, _07713_);
  or (_07716_, _07715_, _07649_);
  or (_07717_, _07666_, _06465_);
  and (_26879_[4], _07717_, _07716_);
  or (_07718_, _07660_, word_in[13]);
  not (_07719_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_07720_, _07655_, _07719_);
  and (_07721_, _07655_, word_in[5]);
  or (_07722_, _07721_, _07720_);
  or (_07723_, _07722_, _07653_);
  and (_07724_, _07723_, _07651_);
  and (_07725_, _07724_, _07718_);
  and (_07726_, _07650_, _06477_);
  or (_07727_, _07726_, _07649_);
  or (_07728_, _07727_, _07725_);
  or (_07729_, _07666_, _05950_);
  and (_26879_[5], _07729_, _07728_);
  and (_07730_, _05551_, _26170_);
  and (_07731_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_02516_, _07731_, _07730_);
  and (_07732_, _07650_, _06492_);
  and (_07733_, _07655_, word_in[6]);
  not (_07734_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_07735_, _07655_, _07734_);
  nor (_07736_, _07735_, _07733_);
  nor (_07737_, _07736_, _07653_);
  and (_07738_, _07653_, word_in[14]);
  or (_07739_, _07738_, _07737_);
  and (_07740_, _07739_, _07651_);
  or (_07741_, _07740_, _07732_);
  and (_07742_, _07741_, _07666_);
  and (_07743_, _07649_, _05968_);
  or (_26879_[6], _07743_, _07742_);
  and (_07744_, _07650_, _05340_);
  and (_07745_, _07655_, word_in[7]);
  nor (_07746_, _07655_, _05018_);
  nor (_07747_, _07746_, _07745_);
  nor (_07748_, _07747_, _07653_);
  and (_07749_, _07653_, word_in[15]);
  or (_07750_, _07749_, _07748_);
  and (_07751_, _07750_, _07651_);
  or (_07752_, _07751_, _07744_);
  and (_07753_, _07752_, _07666_);
  and (_07754_, _07649_, _05348_);
  or (_26879_[7], _07754_, _07753_);
  and (_07755_, _05337_, _05065_);
  not (_07756_, _07755_);
  and (_07757_, _07527_, _05063_);
  and (_07758_, _07757_, _05862_);
  not (_07759_, _07757_);
  and (_07760_, _06127_, _05095_);
  and (_07761_, _06131_, _05313_);
  and (_07762_, _07761_, word_in[0]);
  not (_07763_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_07764_, _07761_, _07763_);
  nor (_07765_, _07764_, _07762_);
  nor (_07766_, _07765_, _07760_);
  and (_07767_, _07760_, word_in[8]);
  or (_07768_, _07767_, _07766_);
  and (_07769_, _07768_, _07759_);
  or (_07770_, _07769_, _07758_);
  and (_07771_, _07770_, _07756_);
  and (_07772_, _07755_, _07407_);
  or (_26880_[0], _07772_, _07771_);
  and (_07773_, _07757_, _06415_);
  not (_07774_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_07775_, _07761_, _07774_);
  and (_07776_, _07761_, word_in[1]);
  nor (_07777_, _07776_, _07775_);
  nor (_07778_, _07777_, _07760_);
  and (_07779_, _07760_, word_in[9]);
  or (_07780_, _07779_, _07778_);
  and (_07781_, _07780_, _07759_);
  or (_07782_, _07781_, _07773_);
  and (_07783_, _07782_, _07756_);
  and (_07784_, _07755_, _05870_);
  or (_26880_[1], _07784_, _07783_);
  and (_07785_, _07757_, _06431_);
  not (_07786_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_07787_, _07761_, _07786_);
  and (_07788_, _07761_, word_in[2]);
  nor (_07789_, _07788_, _07787_);
  nor (_07790_, _07789_, _07760_);
  and (_07791_, _07760_, word_in[10]);
  or (_07792_, _07791_, _07790_);
  and (_07793_, _07792_, _07759_);
  or (_07794_, _07793_, _07785_);
  and (_07795_, _07794_, _07756_);
  and (_07796_, _07755_, _05903_);
  or (_26880_[2], _07796_, _07795_);
  and (_07797_, _07757_, _06439_);
  not (_07798_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_07799_, _07761_, _07798_);
  and (_07800_, _07761_, word_in[3]);
  nor (_07801_, _07800_, _07799_);
  nor (_07802_, _07801_, _07760_);
  and (_07803_, _07760_, word_in[11]);
  or (_07804_, _07803_, _07802_);
  and (_07805_, _07804_, _07759_);
  or (_07806_, _07805_, _07797_);
  and (_07807_, _07806_, _07756_);
  and (_07808_, _07755_, _05919_);
  or (_26880_[3], _07808_, _07807_);
  and (_07809_, _07757_, _06461_);
  not (_07810_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_07811_, _07761_, _07810_);
  and (_07812_, _07761_, word_in[4]);
  nor (_07813_, _07812_, _07811_);
  nor (_07814_, _07813_, _07760_);
  and (_07815_, _07760_, word_in[12]);
  or (_07816_, _07815_, _07814_);
  and (_07817_, _07816_, _07759_);
  or (_07818_, _07817_, _07809_);
  and (_07819_, _07818_, _07756_);
  and (_07820_, _07755_, _06465_);
  or (_26880_[4], _07820_, _07819_);
  and (_07821_, _07757_, _06477_);
  not (_07822_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_07823_, _07761_, _07822_);
  and (_07824_, _07761_, word_in[5]);
  nor (_07825_, _07824_, _07823_);
  nor (_07826_, _07825_, _07760_);
  and (_07827_, _07760_, word_in[13]);
  or (_07829_, _07827_, _07826_);
  and (_07830_, _07829_, _07759_);
  or (_07831_, _07830_, _07821_);
  and (_07833_, _07831_, _07756_);
  and (_07834_, _07755_, _05950_);
  or (_26880_[5], _07834_, _07833_);
  or (_07835_, _07759_, _06492_);
  not (_07836_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_07837_, _07761_, _07836_);
  and (_07838_, _07761_, word_in[6]);
  or (_07839_, _07838_, _07837_);
  or (_07840_, _07839_, _07760_);
  not (_07841_, _07760_);
  or (_07842_, _07841_, word_in[14]);
  and (_07843_, _07842_, _07840_);
  or (_07845_, _07843_, _07757_);
  and (_07847_, _07845_, _07835_);
  or (_07848_, _07847_, _07755_);
  or (_07850_, _07756_, _05968_);
  and (_26880_[6], _07850_, _07848_);
  and (_07852_, _07757_, _05340_);
  nor (_07853_, _07761_, _05138_);
  and (_07855_, _07761_, word_in[7]);
  nor (_07856_, _07855_, _07853_);
  nor (_07858_, _07856_, _07760_);
  and (_07859_, _07760_, word_in[15]);
  or (_07860_, _07859_, _07858_);
  and (_07861_, _07860_, _07759_);
  or (_07862_, _07861_, _07852_);
  and (_07863_, _07862_, _07756_);
  and (_07864_, _07755_, _05348_);
  or (_26880_[7], _07864_, _07863_);
  and (_07865_, _05755_, _23768_);
  and (_07866_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_02597_, _07866_, _07865_);
  and (_07867_, _26341_, _26085_);
  and (_07868_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_02621_, _07868_, _07867_);
  and (_07869_, _26341_, _23830_);
  and (_07870_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_02627_, _07870_, _07869_);
  and (_07871_, _05862_, _05318_);
  not (_07872_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_07873_, _05327_, _07872_);
  and (_07874_, _05327_, word_in[0]);
  nor (_07875_, _07874_, _07873_);
  nor (_07876_, _07875_, _05322_);
  and (_07877_, _05322_, word_in[8]);
  or (_07878_, _07877_, _07876_);
  and (_07879_, _07878_, _05319_);
  or (_07880_, _07879_, _07871_);
  and (_07881_, _07880_, _05346_);
  and (_07882_, _07407_, _05338_);
  or (_26881_[0], _07882_, _07881_);
  not (_07883_, _05322_);
  or (_07884_, _07883_, word_in[9]);
  not (_07885_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_07886_, _05327_, _07885_);
  and (_07887_, _05875_, _05327_);
  or (_07888_, _07887_, _07886_);
  or (_07889_, _07888_, _05322_);
  and (_07890_, _07889_, _07884_);
  or (_07891_, _07890_, _05318_);
  or (_07892_, _06415_, _05319_);
  and (_07893_, _07892_, _07891_);
  or (_07894_, _07893_, _05338_);
  or (_07895_, _05870_, _05346_);
  and (_26881_[1], _07895_, _07894_);
  or (_07897_, _07883_, word_in[10]);
  not (_07898_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_07899_, _05327_, _07898_);
  and (_07900_, _05892_, _05327_);
  or (_07901_, _07900_, _07899_);
  or (_07902_, _07901_, _05322_);
  and (_07903_, _07902_, _07897_);
  or (_07905_, _07903_, _05318_);
  or (_07907_, _06431_, _05319_);
  and (_07908_, _07907_, _07905_);
  or (_07910_, _07908_, _05338_);
  or (_07911_, _05903_, _05346_);
  and (_26881_[2], _07911_, _07910_);
  and (_07914_, _06439_, _05318_);
  not (_07916_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_07917_, _05327_, _07916_);
  and (_07918_, _05327_, word_in[3]);
  nor (_07920_, _07918_, _07917_);
  nor (_07921_, _07920_, _05322_);
  and (_07922_, _05322_, word_in[11]);
  or (_07923_, _07922_, _07921_);
  and (_07924_, _07923_, _05319_);
  or (_07926_, _07924_, _07914_);
  and (_07927_, _07926_, _05346_);
  and (_07928_, _05919_, _05338_);
  or (_26881_[3], _07928_, _07927_);
  or (_07930_, _07883_, word_in[12]);
  not (_07931_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_07933_, _05327_, _07931_);
  and (_07934_, _06061_, _05327_);
  or (_07935_, _07934_, _07933_);
  or (_07937_, _07935_, _05322_);
  and (_07938_, _07937_, _07930_);
  or (_07940_, _07938_, _05318_);
  or (_07941_, _06461_, _05319_);
  and (_07943_, _07941_, _07940_);
  or (_07944_, _07943_, _05338_);
  or (_07945_, _06465_, _05346_);
  and (_26881_[4], _07945_, _07944_);
  or (_07948_, _07883_, word_in[13]);
  not (_07950_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_07951_, _05327_, _07950_);
  and (_07953_, _05939_, _05327_);
  or (_07954_, _07953_, _07951_);
  or (_07955_, _07954_, _05322_);
  and (_07956_, _07955_, _07948_);
  or (_07957_, _07956_, _05318_);
  or (_07958_, _06477_, _05319_);
  and (_07959_, _07958_, _07957_);
  or (_07960_, _07959_, _05338_);
  or (_07961_, _05950_, _05346_);
  and (_26881_[5], _07961_, _07960_);
  and (_07962_, _06492_, _05318_);
  not (_07963_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_07964_, _05327_, _07963_);
  and (_07965_, _05327_, word_in[6]);
  nor (_07966_, _07965_, _07964_);
  nor (_07967_, _07966_, _05322_);
  and (_07968_, _05322_, word_in[14]);
  or (_07969_, _07968_, _07967_);
  and (_07970_, _07969_, _05319_);
  or (_07971_, _07970_, _07962_);
  and (_07972_, _07971_, _05346_);
  and (_07973_, _05968_, _05338_);
  or (_26881_[6], _07973_, _07972_);
  and (_07974_, _04159_, _26170_);
  and (_07975_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_02697_, _07975_, _07974_);
  and (_07976_, _05004_, word_in[0]);
  nand (_07977_, _04931_, _06822_);
  or (_07978_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_07979_, _07978_, _07977_);
  and (_07980_, _07979_, _04966_);
  nand (_07981_, _04931_, _06009_);
  or (_07982_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_07983_, _07982_, _07981_);
  and (_07984_, _07983_, _04939_);
  or (_07985_, _07984_, _07980_);
  nand (_07986_, _04931_, _06532_);
  or (_07987_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_07988_, _07987_, _07986_);
  and (_07989_, _07988_, _04955_);
  nand (_07990_, _04931_, _06255_);
  or (_07991_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_07992_, _07991_, _07990_);
  and (_07993_, _07992_, _04959_);
  or (_07994_, _07993_, _07989_);
  or (_07995_, _07994_, _07985_);
  and (_07996_, _07995_, _04978_);
  nand (_07997_, _04931_, _07654_);
  or (_07998_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_07999_, _07998_, _07997_);
  and (_08001_, _07999_, _04955_);
  nand (_08002_, _04931_, _07116_);
  or (_08003_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_08004_, _08003_, _08002_);
  and (_08005_, _08004_, _04939_);
  or (_08006_, _08005_, _08001_);
  and (_08007_, _08006_, _04944_);
  and (_08008_, _04944_, _04959_);
  nand (_08009_, _04931_, _07388_);
  or (_08010_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_08011_, _08010_, _08009_);
  and (_08012_, _08011_, _08008_);
  or (_08013_, _08012_, _08007_);
  nand (_08014_, _04931_, _07872_);
  or (_08015_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08016_, _08015_, _08014_);
  and (_08017_, _08016_, _05183_);
  or (_08018_, _08017_, _08013_);
  or (_08019_, _08018_, _07996_);
  and (_08020_, _08019_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08020_, _07976_);
  and (_08021_, _05004_, word_in[1]);
  nand (_08022_, _04931_, _06840_);
  or (_08023_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_08024_, _08023_, _08022_);
  and (_08025_, _08024_, _04966_);
  nand (_08026_, _04931_, _06269_);
  or (_08027_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_08028_, _08027_, _08026_);
  and (_08029_, _08028_, _04959_);
  or (_08030_, _08029_, _08025_);
  nand (_08031_, _04931_, _06554_);
  or (_08032_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_08033_, _08032_, _08031_);
  and (_08034_, _08033_, _04955_);
  nand (_08035_, _04931_, _06020_);
  or (_08036_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_08037_, _08036_, _08035_);
  and (_08038_, _08037_, _04939_);
  or (_08039_, _08038_, _08034_);
  or (_08040_, _08039_, _08030_);
  and (_08041_, _08040_, _04978_);
  nand (_08042_, _04931_, _07668_);
  or (_08043_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_08044_, _08043_, _08042_);
  and (_08045_, _08044_, _04955_);
  nand (_08046_, _04931_, _07413_);
  or (_08047_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_08048_, _08047_, _08046_);
  and (_08049_, _08048_, _04959_);
  or (_08050_, _08049_, _08045_);
  and (_08051_, _08050_, _04944_);
  nand (_08052_, _04931_, _07126_);
  or (_08053_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_08054_, _08053_, _08052_);
  and (_08055_, _08054_, _05728_);
  or (_08056_, _08055_, _08051_);
  nand (_08057_, _04931_, _07885_);
  or (_08058_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_08059_, _08058_, _08057_);
  and (_08060_, _08059_, _05183_);
  or (_08061_, _08060_, _08056_);
  or (_08062_, _08061_, _08041_);
  and (_08063_, _08062_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08063_, _08021_);
  and (_08064_, _05004_, word_in[2]);
  nand (_08065_, _04931_, _06857_);
  or (_08066_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_08067_, _08066_, _08065_);
  and (_08068_, _08067_, _04966_);
  nand (_08069_, _04931_, _06281_);
  or (_08070_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_08071_, _08070_, _08069_);
  and (_08072_, _08071_, _04959_);
  or (_08073_, _08072_, _08068_);
  nand (_08074_, _04931_, _06572_);
  or (_08075_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_08076_, _08075_, _08074_);
  and (_08077_, _08076_, _04955_);
  nand (_08078_, _04931_, _06036_);
  or (_08079_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_08080_, _08079_, _08078_);
  and (_08081_, _08080_, _04939_);
  or (_08082_, _08081_, _08077_);
  or (_08083_, _08082_, _08073_);
  and (_08084_, _08083_, _04978_);
  nand (_08085_, _04931_, _07681_);
  or (_08086_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_08087_, _08086_, _08085_);
  and (_08088_, _08087_, _04955_);
  nand (_08089_, _04931_, _07143_);
  or (_08090_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_08091_, _08090_, _08089_);
  and (_08092_, _08091_, _04939_);
  or (_08093_, _08092_, _08088_);
  and (_08094_, _08093_, _04944_);
  nand (_08095_, _04931_, _07430_);
  or (_08096_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_08097_, _08096_, _08095_);
  and (_08098_, _08097_, _08008_);
  or (_08100_, _08098_, _08094_);
  nand (_08101_, _04931_, _07898_);
  or (_08102_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_08103_, _08102_, _08101_);
  and (_08104_, _08103_, _05183_);
  or (_08105_, _08104_, _08100_);
  or (_08106_, _08105_, _08084_);
  and (_08107_, _08106_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08107_, _08064_);
  and (_08108_, _05004_, word_in[3]);
  nand (_08109_, _04931_, _06869_);
  or (_08110_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_08111_, _08110_, _08109_);
  and (_08112_, _08111_, _04966_);
  nand (_08113_, _04931_, _06299_);
  or (_08114_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_08115_, _08114_, _08113_);
  and (_08116_, _08115_, _04959_);
  or (_08117_, _08116_, _08112_);
  nand (_08118_, _04931_, _06590_);
  or (_08119_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_08120_, _08119_, _08118_);
  and (_08121_, _08120_, _04955_);
  nand (_08122_, _04931_, _06048_);
  or (_08123_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_08124_, _08123_, _08122_);
  and (_08125_, _08124_, _04939_);
  or (_08126_, _08125_, _08121_);
  or (_08127_, _08126_, _08117_);
  and (_08128_, _08127_, _04978_);
  nand (_08129_, _04931_, _07693_);
  or (_08130_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_08131_, _08130_, _08129_);
  and (_08132_, _08131_, _04955_);
  nand (_08133_, _04931_, _07158_);
  or (_08134_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_08135_, _08134_, _08133_);
  and (_08136_, _08135_, _04939_);
  or (_08137_, _08136_, _08132_);
  and (_08138_, _08137_, _04944_);
  nand (_08139_, _04931_, _07444_);
  or (_08140_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_08141_, _08140_, _08139_);
  and (_08142_, _08141_, _08008_);
  or (_08143_, _08142_, _08138_);
  nand (_08144_, _04931_, _07916_);
  or (_08145_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_08146_, _08145_, _08144_);
  and (_08147_, _08146_, _05183_);
  or (_08148_, _08147_, _08143_);
  or (_08149_, _08148_, _08128_);
  and (_08150_, _08149_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08150_, _08108_);
  and (_08151_, _05004_, word_in[4]);
  nand (_08152_, _04931_, _06606_);
  or (_08153_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_08154_, _08153_, _08152_);
  and (_08155_, _08154_, _04955_);
  nand (_08156_, _04931_, _06063_);
  or (_08157_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_08158_, _08157_, _08156_);
  and (_08159_, _08158_, _04939_);
  or (_08160_, _08159_, _08155_);
  nand (_08161_, _04931_, _06885_);
  or (_08162_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_08163_, _08162_, _08161_);
  and (_08164_, _08163_, _04966_);
  nand (_08165_, _04931_, _06312_);
  or (_08166_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_08167_, _08166_, _08165_);
  and (_08168_, _08167_, _04959_);
  or (_08169_, _08168_, _08164_);
  or (_08170_, _08169_, _08160_);
  and (_08171_, _08170_, _04978_);
  nand (_08172_, _04931_, _07705_);
  or (_08173_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_08174_, _08173_, _08172_);
  and (_08175_, _08174_, _04955_);
  nand (_08176_, _04931_, _07172_);
  or (_08177_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_08178_, _08177_, _08176_);
  and (_08179_, _08178_, _04939_);
  or (_08180_, _08179_, _08175_);
  and (_08181_, _08180_, _04944_);
  nand (_08182_, _04931_, _07931_);
  or (_08183_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _05183_);
  nand (_08186_, _04931_, _07457_);
  or (_08187_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_08189_, _08187_, _08186_);
  and (_08190_, _08189_, _08008_);
  or (_08191_, _08190_, _08185_);
  or (_08192_, _08191_, _08181_);
  or (_08193_, _08192_, _08171_);
  and (_08194_, _08193_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08194_, _08151_);
  and (_08196_, _05004_, word_in[5]);
  nand (_08197_, _04931_, _06903_);
  or (_08199_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_08202_, _08199_, _08197_);
  and (_08203_, _08202_, _04966_);
  nand (_08204_, _04931_, _06325_);
  or (_08205_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_08206_, _08205_, _08204_);
  and (_08208_, _08206_, _04959_);
  or (_08210_, _08208_, _08203_);
  nand (_08211_, _04931_, _06621_);
  or (_08212_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_08214_, _08212_, _08211_);
  and (_08215_, _08214_, _04955_);
  nand (_08216_, _04931_, _06078_);
  or (_08217_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_08218_, _08217_, _08216_);
  and (_08219_, _08218_, _04939_);
  or (_08220_, _08219_, _08215_);
  or (_08222_, _08220_, _08210_);
  and (_08223_, _08222_, _04978_);
  nand (_08224_, _04931_, _07719_);
  or (_08225_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_08226_, _08225_, _08224_);
  and (_08227_, _08226_, _04955_);
  nand (_08228_, _04931_, _07188_);
  or (_08229_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_08230_, _08229_, _08228_);
  and (_08231_, _08230_, _04939_);
  or (_08232_, _08231_, _08227_);
  and (_08233_, _08232_, _04944_);
  nand (_08234_, _04931_, _07475_);
  or (_08235_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_08236_, _08235_, _08234_);
  and (_08237_, _08236_, _08008_);
  or (_08238_, _08237_, _08233_);
  nand (_08239_, _04931_, _07950_);
  or (_08240_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_08241_, _08240_, _08239_);
  and (_08242_, _08241_, _05183_);
  or (_08243_, _08242_, _08238_);
  or (_08244_, _08243_, _08223_);
  and (_08245_, _08244_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08245_, _08196_);
  and (_08246_, _05004_, word_in[6]);
  nand (_08247_, _04931_, _06918_);
  or (_08248_, _04931_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_08249_, _08248_, _08247_);
  and (_08250_, _08249_, _04966_);
  nand (_08251_, _04931_, _06091_);
  or (_08252_, _04931_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_08253_, _08252_, _08251_);
  and (_08254_, _08253_, _04939_);
  or (_08255_, _08254_, _08250_);
  nand (_08256_, _04931_, _06636_);
  or (_08257_, _04931_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_08258_, _08257_, _08256_);
  and (_08259_, _08258_, _04955_);
  nand (_08260_, _04931_, _06338_);
  or (_08261_, _04931_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_08262_, _08261_, _08260_);
  and (_08263_, _08262_, _04959_);
  or (_08264_, _08263_, _08259_);
  or (_08265_, _08264_, _08255_);
  and (_08266_, _08265_, _04978_);
  nand (_08267_, _04931_, _07734_);
  or (_08268_, _04931_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_08269_, _08268_, _08267_);
  and (_08270_, _08269_, _04955_);
  nand (_08271_, _04931_, _07204_);
  or (_08272_, _04931_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_08273_, _08272_, _08271_);
  and (_08274_, _08273_, _04939_);
  or (_08275_, _08274_, _08270_);
  and (_08276_, _08275_, _04944_);
  nand (_08277_, _04931_, _07492_);
  or (_08278_, _04931_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_08279_, _08278_, _08277_);
  and (_08280_, _08279_, _08008_);
  or (_08281_, _08280_, _08276_);
  nand (_08282_, _04931_, _07963_);
  or (_08283_, _04931_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_08284_, _08283_, _08282_);
  and (_08285_, _08284_, _05183_);
  or (_08286_, _08285_, _08281_);
  or (_08287_, _08286_, _08266_);
  and (_08288_, _08287_, _05003_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08288_, _08246_);
  and (_08289_, _26224_, _26193_);
  and (_08290_, _08289_, _26085_);
  not (_08291_, _08289_);
  and (_08292_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_02737_, _08292_, _08290_);
  and (_08294_, _05121_, word_in[8]);
  nand (_08295_, _04931_, _07238_);
  or (_08296_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_08297_, _08296_, _08295_);
  and (_08298_, _08297_, _05124_);
  nand (_08299_, _04931_, _06956_);
  or (_08300_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_08301_, _08300_, _08299_);
  and (_08302_, _08301_, _05122_);
  or (_08303_, _08302_, _08298_);
  and (_08304_, _08303_, _05076_);
  nand (_08305_, _04931_, _06134_);
  or (_08306_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_08307_, _08306_, _08305_);
  and (_08309_, _08307_, _05124_);
  nand (_08311_, _04931_, _05850_);
  or (_08312_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_08314_, _08312_, _08311_);
  and (_08315_, _08314_, _05122_);
  or (_08317_, _08315_, _08309_);
  and (_08318_, _08317_, _05079_);
  nand (_08319_, _04931_, _06687_);
  or (_08320_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_08321_, _08320_, _08319_);
  and (_08322_, _08321_, _05124_);
  nand (_08323_, _04931_, _06388_);
  or (_08324_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_08325_, _08324_, _08323_);
  and (_08326_, _08325_, _05122_);
  or (_08327_, _08326_, _08322_);
  and (_08329_, _08327_, _05100_);
  or (_08330_, _08329_, _08318_);
  nand (_08331_, _04931_, _07763_);
  or (_08332_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_08333_, _08332_, _08331_);
  and (_08334_, _08333_, _05124_);
  nand (_08335_, _04931_, _07534_);
  or (_08336_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_08337_, _08336_, _08335_);
  and (_08338_, _08337_, _05122_);
  or (_08339_, _08338_, _08334_);
  and (_08340_, _08339_, _05095_);
  or (_08341_, _08340_, _08330_);
  nor (_08342_, _08341_, _08304_);
  nor (_08343_, _08342_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08343_, _08294_);
  and (_08344_, _05121_, word_in[9]);
  nand (_08345_, _04931_, _07259_);
  or (_08346_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_08347_, _08346_, _08345_);
  and (_08349_, _08347_, _05124_);
  nand (_08350_, _04931_, _06980_);
  or (_08351_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_08352_, _08351_, _08350_);
  and (_08353_, _08352_, _05122_);
  or (_08354_, _08353_, _08349_);
  and (_08355_, _08354_, _05076_);
  nand (_08356_, _04931_, _07774_);
  or (_08357_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_08358_, _08357_, _08356_);
  and (_08359_, _08358_, _05124_);
  nand (_08361_, _04931_, _07555_);
  or (_08362_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_08363_, _08362_, _08361_);
  and (_08364_, _08363_, _05122_);
  or (_08365_, _08364_, _08359_);
  and (_08366_, _08365_, _05095_);
  nand (_08367_, _04931_, _06699_);
  or (_08368_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_08369_, _08368_, _08367_);
  and (_08370_, _08369_, _05124_);
  nand (_08371_, _04931_, _06405_);
  or (_08372_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_08373_, _08372_, _08371_);
  and (_08374_, _08373_, _05122_);
  or (_08375_, _08374_, _08370_);
  and (_08376_, _08375_, _05100_);
  nand (_08377_, _04931_, _06147_);
  or (_08378_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_08379_, _08378_, _08377_);
  and (_08380_, _08379_, _05124_);
  nand (_08381_, _04931_, _05872_);
  or (_08382_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_08383_, _08382_, _08381_);
  and (_08384_, _08383_, _05122_);
  or (_08385_, _08384_, _08380_);
  and (_08386_, _08385_, _05079_);
  or (_08387_, _08386_, _08376_);
  or (_08388_, _08387_, _08366_);
  nor (_08390_, _08388_, _08355_);
  nor (_08391_, _08390_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _08391_, _08344_);
  and (_08392_, _05121_, word_in[10]);
  nand (_08393_, _04931_, _07271_);
  or (_08394_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_08395_, _08394_, _08393_);
  and (_08396_, _08395_, _05124_);
  nand (_08397_, _04931_, _06997_);
  or (_08398_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_08399_, _08398_, _08397_);
  and (_08401_, _08399_, _05122_);
  or (_08402_, _08401_, _08396_);
  and (_08403_, _08402_, _05076_);
  nand (_08404_, _04931_, _06158_);
  or (_08405_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_08406_, _08405_, _08404_);
  and (_08407_, _08406_, _05124_);
  nand (_08408_, _04931_, _05889_);
  or (_08409_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_08410_, _08409_, _08408_);
  and (_08412_, _08410_, _05122_);
  or (_08413_, _08412_, _08407_);
  and (_08414_, _08413_, _05079_);
  nand (_08415_, _04931_, _06714_);
  or (_08416_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_08417_, _08416_, _08415_);
  and (_08418_, _08417_, _05124_);
  nand (_08419_, _04931_, _06420_);
  or (_08420_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_08421_, _08420_, _08419_);
  and (_08422_, _08421_, _05122_);
  or (_08423_, _08422_, _08418_);
  and (_08424_, _08423_, _05100_);
  or (_08425_, _08424_, _08414_);
  nand (_08426_, _04931_, _07786_);
  or (_08427_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_08428_, _08427_, _08426_);
  and (_08429_, _08428_, _05124_);
  nand (_08430_, _04931_, _07567_);
  or (_08431_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_08432_, _08431_, _08430_);
  and (_08433_, _08432_, _05122_);
  or (_08434_, _08433_, _08429_);
  and (_08435_, _08434_, _05095_);
  or (_08436_, _08435_, _08425_);
  nor (_08437_, _08436_, _08403_);
  nor (_08438_, _08437_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _08438_, _08392_);
  and (_08439_, _05121_, word_in[11]);
  nand (_08440_, _04931_, _07291_);
  or (_08441_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_08442_, _08441_, _08440_);
  and (_08443_, _08442_, _05124_);
  nand (_08444_, _04931_, _07016_);
  or (_08445_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_08446_, _08445_, _08444_);
  and (_08447_, _08446_, _05122_);
  or (_08448_, _08447_, _08443_);
  and (_08449_, _08448_, _05076_);
  nand (_08450_, _04931_, _06170_);
  or (_08451_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_08452_, _08451_, _08450_);
  and (_08453_, _08452_, _05124_);
  nand (_08454_, _04931_, _05905_);
  or (_08455_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_08456_, _08455_, _08454_);
  and (_08457_, _08456_, _05122_);
  or (_08458_, _08457_, _08453_);
  and (_08459_, _08458_, _05079_);
  nand (_08460_, _04931_, _06731_);
  or (_08461_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_08462_, _08461_, _08460_);
  and (_08464_, _08462_, _05124_);
  nand (_08465_, _04931_, _06442_);
  or (_08466_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_08467_, _08466_, _08465_);
  and (_08468_, _08467_, _05122_);
  or (_08469_, _08468_, _08464_);
  and (_08470_, _08469_, _05100_);
  or (_08471_, _08470_, _08459_);
  nand (_08472_, _04931_, _07798_);
  or (_08473_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_08474_, _08473_, _08472_);
  and (_08475_, _08474_, _05124_);
  nand (_08476_, _04931_, _07578_);
  or (_08477_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_08479_, _08477_, _08476_);
  and (_08480_, _08479_, _05122_);
  or (_08482_, _08480_, _08475_);
  and (_08483_, _08482_, _05095_);
  or (_08484_, _08483_, _08471_);
  nor (_08485_, _08484_, _08449_);
  nor (_08486_, _08485_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _08486_, _08439_);
  and (_08487_, _05121_, word_in[12]);
  nand (_08488_, _04931_, _07305_);
  or (_08489_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_08490_, _08489_, _08488_);
  and (_08491_, _08490_, _05124_);
  nand (_08492_, _04931_, _07032_);
  or (_08493_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_08494_, _08493_, _08492_);
  and (_08495_, _08494_, _05122_);
  or (_08496_, _08495_, _08491_);
  and (_08497_, _08496_, _05076_);
  nand (_08498_, _04931_, _06185_);
  or (_08499_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_08500_, _08499_, _08498_);
  and (_08501_, _08500_, _05124_);
  nand (_08502_, _04931_, _05925_);
  or (_08503_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_08504_, _08503_, _08502_);
  and (_08505_, _08504_, _05122_);
  or (_08506_, _08505_, _08501_);
  and (_08508_, _08506_, _05079_);
  nand (_08509_, _04931_, _06746_);
  or (_08510_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_08512_, _08510_, _08509_);
  and (_08514_, _08512_, _05124_);
  nand (_08515_, _04931_, _06453_);
  or (_08516_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_08517_, _08516_, _08515_);
  and (_08518_, _08517_, _05122_);
  or (_08519_, _08518_, _08514_);
  and (_08520_, _08519_, _05100_);
  or (_08521_, _08520_, _08508_);
  nand (_08522_, _04931_, _07810_);
  or (_08523_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_08525_, _08523_, _08522_);
  and (_08526_, _08525_, _05124_);
  nand (_08528_, _04931_, _07593_);
  or (_08529_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _05122_);
  or (_08532_, _08531_, _08526_);
  and (_08533_, _08532_, _05095_);
  or (_08534_, _08533_, _08521_);
  nor (_08535_, _08534_, _08497_);
  nor (_08536_, _08535_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _08536_, _08487_);
  and (_08538_, _05121_, word_in[13]);
  nand (_08539_, _04931_, _07321_);
  or (_08540_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_08541_, _08540_, _08539_);
  and (_08542_, _08541_, _05124_);
  nand (_08543_, _04931_, _07051_);
  or (_08544_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_08545_, _08544_, _08543_);
  and (_08546_, _08545_, _05122_);
  or (_08547_, _08546_, _08542_);
  and (_08548_, _08547_, _05076_);
  nand (_08549_, _04931_, _06201_);
  or (_08550_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_08551_, _08550_, _08549_);
  and (_08552_, _08551_, _05124_);
  nand (_08553_, _04931_, _05937_);
  or (_08554_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_08555_, _08554_, _08553_);
  and (_08556_, _08555_, _05122_);
  or (_08558_, _08556_, _08552_);
  and (_08559_, _08558_, _05079_);
  nand (_08560_, _04931_, _06763_);
  or (_08561_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_08562_, _08561_, _08560_);
  and (_08563_, _08562_, _05124_);
  nand (_08564_, _04931_, _06467_);
  or (_08565_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_08566_, _08565_, _08564_);
  and (_08567_, _08566_, _05122_);
  or (_08568_, _08567_, _08563_);
  and (_08570_, _08568_, _05100_);
  or (_08571_, _08570_, _08559_);
  nand (_08572_, _04931_, _07822_);
  or (_08573_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_08574_, _08573_, _08572_);
  and (_08575_, _08574_, _05124_);
  nand (_08576_, _04931_, _07608_);
  or (_08577_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_08578_, _08577_, _08576_);
  and (_08579_, _08578_, _05122_);
  or (_08580_, _08579_, _08575_);
  and (_08581_, _08580_, _05095_);
  or (_08583_, _08581_, _08571_);
  nor (_08584_, _08583_, _08548_);
  nor (_08585_, _08584_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _08585_, _08538_);
  and (_08586_, _05121_, word_in[14]);
  nand (_08587_, _04931_, _07339_);
  or (_08589_, _04931_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_08590_, _08589_, _08587_);
  and (_08592_, _08590_, _05124_);
  nand (_08593_, _04931_, _07073_);
  or (_08594_, _04931_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_08595_, _08594_, _08593_);
  and (_08596_, _08595_, _05122_);
  or (_08597_, _08596_, _08592_);
  and (_08598_, _08597_, _05076_);
  nand (_08599_, _04931_, _07836_);
  or (_08600_, _04931_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_08601_, _08600_, _08599_);
  and (_08602_, _08601_, _05124_);
  nand (_08603_, _04931_, _07620_);
  or (_08604_, _04931_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_08605_, _08604_, _08603_);
  and (_08606_, _08605_, _05122_);
  or (_08607_, _08606_, _08602_);
  and (_08608_, _08607_, _05095_);
  nand (_08610_, _04931_, _06778_);
  or (_08611_, _04931_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_08613_, _08611_, _08610_);
  and (_08614_, _08613_, _05124_);
  nand (_08616_, _04931_, _06483_);
  or (_08617_, _04931_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_08618_, _08617_, _08616_);
  and (_08619_, _08618_, _05122_);
  or (_08620_, _08619_, _08614_);
  and (_08621_, _08620_, _05100_);
  nand (_08623_, _04931_, _06214_);
  or (_08624_, _04931_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_08625_, _08624_, _08623_);
  and (_08627_, _08625_, _05124_);
  nand (_08628_, _04931_, _05953_);
  or (_08629_, _04931_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_08630_, _08629_, _08628_);
  and (_08631_, _08630_, _05122_);
  or (_08632_, _08631_, _08627_);
  and (_08633_, _08632_, _05079_);
  or (_08634_, _08633_, _08621_);
  or (_08635_, _08634_, _08608_);
  nor (_08636_, _08635_, _08598_);
  nor (_08637_, _08636_, _05121_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _08637_, _08586_);
  and (_08638_, _23030_, _22949_);
  and (_08639_, _24146_, _23027_);
  and (_08640_, _24176_, _22972_);
  or (_08641_, _08640_, _08639_);
  or (_08642_, _08641_, _08638_);
  and (_08643_, _08641_, _22944_);
  or (_08644_, _08643_, _23040_);
  and (_08645_, _08644_, _08642_);
  not (_08646_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_08647_, _23041_, _08646_);
  not (_08648_, _23009_);
  or (_08649_, _05549_, _08648_);
  and (_08650_, _23022_, _22949_);
  not (_08651_, _08650_);
  and (_08652_, _08651_, _08649_);
  not (_08653_, _08652_);
  and (_08654_, _08653_, _08647_);
  or (_08655_, _08654_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_08656_, _08655_, _08645_);
  or (_08657_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _22734_);
  and (_08658_, _08657_, _23049_);
  and (_26901_[2], _08658_, _08656_);
  and (_08659_, _08289_, _23830_);
  and (_08660_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_02765_, _08660_, _08659_);
  and (_08662_, _05218_, word_in[16]);
  and (_08663_, _08016_, _04955_);
  and (_08664_, _07999_, _04959_);
  or (_08666_, _08664_, _08663_);
  and (_08668_, _08004_, _04966_);
  and (_08670_, _08011_, _04939_);
  or (_08671_, _08670_, _08668_);
  or (_08673_, _08671_, _08666_);
  or (_08674_, _08673_, _05219_);
  and (_08676_, _07988_, _04959_);
  and (_08678_, _07992_, _04939_);
  or (_08679_, _08678_, _08676_);
  and (_08681_, _07979_, _04955_);
  and (_08683_, _07983_, _04966_);
  or (_08685_, _08683_, _08681_);
  or (_08687_, _08685_, _08679_);
  or (_08689_, _08687_, _05185_);
  nand (_08690_, _08689_, _08674_);
  nor (_08692_, _08690_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _08692_, _08662_);
  and (_08695_, _05218_, word_in[17]);
  and (_08697_, _08024_, _04955_);
  and (_08698_, _08033_, _04959_);
  or (_08700_, _08698_, _08697_);
  and (_08702_, _08037_, _04966_);
  and (_08703_, _08028_, _04939_);
  or (_08704_, _08703_, _08702_);
  or (_08706_, _08704_, _08700_);
  or (_08708_, _08706_, _05185_);
  and (_08710_, _08044_, _04959_);
  and (_08711_, _08048_, _04939_);
  or (_08712_, _08711_, _08710_);
  and (_08714_, _08059_, _04955_);
  and (_08716_, _08054_, _04966_);
  or (_08717_, _08716_, _08714_);
  or (_08718_, _08717_, _08712_);
  or (_08719_, _08718_, _05219_);
  nand (_08720_, _08719_, _08708_);
  nor (_08722_, _08720_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _08722_, _08695_);
  and (_08723_, _05218_, word_in[18]);
  and (_08725_, _08067_, _04955_);
  and (_08726_, _08076_, _04959_);
  or (_08727_, _08726_, _08725_);
  and (_08728_, _08080_, _04966_);
  and (_08729_, _08071_, _04939_);
  or (_08730_, _08729_, _08728_);
  or (_08731_, _08730_, _08727_);
  or (_08732_, _08731_, _05185_);
  and (_08734_, _08087_, _04959_);
  and (_08736_, _08097_, _04939_);
  or (_08737_, _08736_, _08734_);
  and (_08738_, _08103_, _04955_);
  and (_08740_, _08091_, _04966_);
  or (_08742_, _08740_, _08738_);
  or (_08744_, _08742_, _08737_);
  or (_08745_, _08744_, _05219_);
  nand (_08747_, _08745_, _08732_);
  nor (_08749_, _08747_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _08749_, _08723_);
  and (_08750_, _05218_, word_in[19]);
  and (_08752_, _08111_, _04955_);
  and (_08754_, _08120_, _04959_);
  or (_08756_, _08754_, _08752_);
  and (_08758_, _08124_, _04966_);
  and (_08760_, _08115_, _04939_);
  or (_08762_, _08760_, _08758_);
  or (_08763_, _08762_, _08756_);
  or (_08764_, _08763_, _05185_);
  and (_08765_, _08131_, _04959_);
  and (_08766_, _08141_, _04939_);
  or (_08767_, _08766_, _08765_);
  and (_08769_, _08146_, _04955_);
  and (_08771_, _08135_, _04966_);
  or (_08772_, _08771_, _08769_);
  or (_08773_, _08772_, _08767_);
  or (_08774_, _08773_, _05219_);
  nand (_08775_, _08774_, _08764_);
  nor (_08776_, _08775_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _08776_, _08750_);
  and (_08778_, _05218_, word_in[20]);
  and (_08779_, _08184_, _04955_);
  and (_08780_, _08174_, _04959_);
  or (_08782_, _08780_, _08779_);
  and (_08783_, _08178_, _04966_);
  and (_08784_, _08189_, _04939_);
  or (_08786_, _08784_, _08783_);
  or (_08787_, _08786_, _08782_);
  or (_08788_, _08787_, _05219_);
  and (_08790_, _08154_, _04959_);
  and (_08792_, _08167_, _04939_);
  or (_08793_, _08792_, _08790_);
  and (_08794_, _08163_, _04955_);
  and (_08795_, _08158_, _04966_);
  or (_08796_, _08795_, _08794_);
  or (_08798_, _08796_, _08793_);
  or (_08799_, _08798_, _05185_);
  nand (_08800_, _08799_, _08788_);
  nor (_08801_, _08800_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _08801_, _08778_);
  and (_08802_, _05218_, word_in[21]);
  and (_08803_, _08214_, _04959_);
  and (_08804_, _08206_, _04939_);
  or (_08805_, _08804_, _08803_);
  and (_08806_, _08202_, _04955_);
  and (_08807_, _08218_, _04966_);
  or (_08808_, _08807_, _08806_);
  or (_08809_, _08808_, _08805_);
  or (_08810_, _08809_, _05185_);
  and (_08811_, _08226_, _04959_);
  and (_08812_, _08236_, _04939_);
  or (_08813_, _08812_, _08811_);
  and (_08814_, _08241_, _04955_);
  and (_08815_, _08230_, _04966_);
  or (_08816_, _08815_, _08814_);
  or (_08817_, _08816_, _08813_);
  or (_08818_, _08817_, _05219_);
  nand (_08819_, _08818_, _08810_);
  nor (_08820_, _08819_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _08820_, _08802_);
  and (_08822_, _05218_, word_in[22]);
  and (_08823_, _08258_, _04959_);
  and (_08824_, _08262_, _04939_);
  or (_08826_, _08824_, _08823_);
  and (_08827_, _08249_, _04955_);
  and (_08828_, _08253_, _04966_);
  or (_08829_, _08828_, _08827_);
  or (_08830_, _08829_, _08826_);
  or (_08831_, _08830_, _05185_);
  and (_08832_, _08269_, _04959_);
  and (_08833_, _08279_, _04939_);
  or (_08834_, _08833_, _08832_);
  and (_08835_, _08284_, _04955_);
  and (_08836_, _08273_, _04966_);
  or (_08837_, _08836_, _08835_);
  or (_08838_, _08837_, _08834_);
  or (_08839_, _08838_, _05219_);
  nand (_08840_, _08839_, _08831_);
  nor (_08841_, _08840_, _05218_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _08841_, _08822_);
  and (_08842_, _05283_, word_in[24]);
  and (_08843_, _08301_, _05124_);
  and (_08845_, _08297_, _05122_);
  or (_08846_, _08845_, _08843_);
  and (_08847_, _08846_, _05251_);
  and (_08848_, _08314_, _05124_);
  and (_08849_, _08307_, _05122_);
  or (_08850_, _08849_, _08848_);
  and (_08851_, _08850_, _05253_);
  and (_08852_, _08325_, _05124_);
  and (_08854_, _08321_, _05122_);
  or (_08855_, _08854_, _08852_);
  and (_08856_, _08855_, _05293_);
  and (_08857_, _08337_, _05124_);
  and (_08858_, _08333_, _05122_);
  or (_08859_, _08858_, _08857_);
  and (_08860_, _08859_, _05299_);
  or (_08861_, _08860_, _08856_);
  or (_08862_, _08861_, _08851_);
  nor (_08863_, _08862_, _08847_);
  nor (_08864_, _08863_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _08864_, _08842_);
  and (_08866_, _05283_, word_in[25]);
  and (_08867_, _08352_, _05124_);
  and (_08868_, _08347_, _05122_);
  or (_08869_, _08868_, _08867_);
  and (_08870_, _08869_, _05251_);
  and (_08871_, _08383_, _05124_);
  and (_08872_, _08379_, _05122_);
  or (_08873_, _08872_, _08871_);
  and (_08874_, _08873_, _05253_);
  and (_08875_, _08373_, _05124_);
  and (_08876_, _08369_, _05122_);
  or (_08877_, _08876_, _08875_);
  and (_08878_, _08877_, _05293_);
  and (_08879_, _08363_, _05124_);
  and (_08880_, _08358_, _05122_);
  or (_08882_, _08880_, _08879_);
  and (_08883_, _08882_, _05299_);
  or (_08884_, _08883_, _08878_);
  or (_08885_, _08884_, _08874_);
  nor (_08887_, _08885_, _08870_);
  nor (_08888_, _08887_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _08888_, _08866_);
  and (_08890_, _05283_, word_in[26]);
  and (_08891_, _08399_, _05124_);
  and (_08892_, _08395_, _05122_);
  or (_08894_, _08892_, _08891_);
  and (_08895_, _08894_, _05251_);
  and (_08897_, _08410_, _05124_);
  and (_08899_, _08406_, _05122_);
  or (_08901_, _08899_, _08897_);
  and (_08902_, _08901_, _05253_);
  and (_08903_, _08421_, _05124_);
  and (_08905_, _08417_, _05122_);
  or (_08906_, _08905_, _08903_);
  and (_08907_, _08906_, _05293_);
  and (_08909_, _08432_, _05124_);
  and (_08911_, _08428_, _05122_);
  or (_08912_, _08911_, _08909_);
  and (_08913_, _08912_, _05299_);
  or (_08914_, _08913_, _08907_);
  or (_08915_, _08914_, _08902_);
  nor (_08916_, _08915_, _08895_);
  nor (_08917_, _08916_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _08917_, _08890_);
  and (_08918_, _05283_, word_in[27]);
  and (_08919_, _08446_, _05124_);
  and (_08921_, _08442_, _05122_);
  or (_08923_, _08921_, _08919_);
  and (_08924_, _08923_, _05251_);
  and (_08926_, _08456_, _05124_);
  and (_08927_, _08452_, _05122_);
  or (_08928_, _08927_, _08926_);
  and (_08930_, _08928_, _05253_);
  and (_08932_, _08467_, _05124_);
  and (_08934_, _08462_, _05122_);
  or (_08936_, _08934_, _08932_);
  and (_08937_, _08936_, _05293_);
  and (_08938_, _08479_, _05124_);
  and (_08939_, _08474_, _05122_);
  or (_08940_, _08939_, _08938_);
  and (_08942_, _08940_, _05299_);
  or (_08943_, _08942_, _08937_);
  or (_08944_, _08943_, _08930_);
  nor (_08945_, _08944_, _08924_);
  nor (_08946_, _08945_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _08946_, _08918_);
  and (_08947_, _05283_, word_in[28]);
  and (_08948_, _08494_, _05124_);
  and (_08949_, _08490_, _05122_);
  or (_08950_, _08949_, _08948_);
  and (_08951_, _08950_, _05251_);
  and (_08952_, _08504_, _05124_);
  and (_08953_, _08500_, _05122_);
  or (_08954_, _08953_, _08952_);
  and (_08955_, _08954_, _05253_);
  and (_08956_, _08517_, _05124_);
  and (_08957_, _08512_, _05122_);
  or (_08958_, _08957_, _08956_);
  and (_08959_, _08958_, _05293_);
  and (_08960_, _08530_, _05124_);
  and (_08961_, _08525_, _05122_);
  or (_08962_, _08961_, _08960_);
  and (_08963_, _08962_, _05299_);
  or (_08964_, _08963_, _08959_);
  or (_08965_, _08964_, _08955_);
  nor (_08966_, _08965_, _08951_);
  nor (_08967_, _08966_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _08967_, _08947_);
  and (_08968_, _05283_, word_in[29]);
  and (_08969_, _08545_, _05124_);
  and (_08970_, _08541_, _05122_);
  or (_08971_, _08970_, _08969_);
  and (_08972_, _08971_, _05251_);
  and (_08973_, _08555_, _05124_);
  and (_08974_, _08551_, _05122_);
  or (_08975_, _08974_, _08973_);
  and (_08976_, _08975_, _05253_);
  and (_08977_, _08566_, _05124_);
  and (_08978_, _08562_, _05122_);
  or (_08979_, _08978_, _08977_);
  and (_08980_, _08979_, _05293_);
  and (_08981_, _08578_, _05124_);
  and (_08982_, _08574_, _05122_);
  or (_08983_, _08982_, _08981_);
  and (_08985_, _08983_, _05299_);
  or (_08986_, _08985_, _08980_);
  or (_08988_, _08986_, _08976_);
  nor (_08989_, _08988_, _08972_);
  nor (_08991_, _08989_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _08991_, _08968_);
  and (_08993_, _05283_, word_in[30]);
  and (_08994_, _08630_, _05124_);
  and (_08995_, _08625_, _05122_);
  or (_08996_, _08995_, _08994_);
  and (_08998_, _08996_, _05253_);
  and (_08999_, _08595_, _05124_);
  and (_09001_, _08590_, _05122_);
  or (_09003_, _09001_, _08999_);
  and (_09004_, _09003_, _05251_);
  and (_09005_, _08618_, _05124_);
  and (_09006_, _08613_, _05122_);
  or (_09007_, _09006_, _09005_);
  and (_09008_, _09007_, _05293_);
  and (_09009_, _08605_, _05124_);
  and (_09011_, _08601_, _05122_);
  or (_09013_, _09011_, _09009_);
  and (_09014_, _09013_, _05299_);
  or (_09016_, _09014_, _09008_);
  or (_09017_, _09016_, _09004_);
  nor (_09018_, _09017_, _08998_);
  nor (_09019_, _09018_, _05283_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _09019_, _08993_);
  and (_02830_, t1_i, _23049_);
  and (_09021_, _01871_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_09022_, _24163_);
  or (_09023_, _03987_, _09022_);
  and (_09025_, _25071_, _22949_);
  and (_09026_, _23027_, _23017_);
  or (_09028_, _09026_, _09025_);
  or (_09029_, _09028_, _09023_);
  and (_09031_, _08650_, _22973_);
  and (_09032_, _23052_, _23009_);
  or (_09033_, _09032_, _24149_);
  or (_09034_, _09033_, _09031_);
  or (_09035_, _09034_, _09029_);
  and (_09037_, _09035_, _01913_);
  or (_26897_, _09037_, _09021_);
  and (_09040_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_09041_, _04300_, _26242_);
  or (_02889_, _09041_, _09040_);
  and (_09042_, _04915_, _23768_);
  and (_09043_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_02913_, _09043_, _09042_);
  and (_09044_, _08289_, _26242_);
  and (_09045_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_02924_, _09045_, _09044_);
  and (_09047_, _26260_, _26213_);
  not (_09049_, _09047_);
  and (_09050_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_09052_, _09047_, _26185_);
  or (_02981_, _09052_, _09050_);
  and (_09053_, _26421_, _23848_);
  and (_09054_, _09053_, _26242_);
  not (_09056_, _09053_);
  and (_09057_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_27267_, _09057_, _09054_);
  not (_09059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor (_09061_, _26096_, _09059_);
  nand (_09062_, _09061_, _26120_);
  not (_09064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_09066_, _26104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_09067_, _09066_, _09064_);
  or (_09068_, _09067_, _26122_);
  and (_09069_, _09068_, _26095_);
  nand (_09070_, _09069_, _09062_);
  not (_09072_, _05563_);
  and (_09074_, _26093_, _09059_);
  nor (_09076_, _09074_, _09072_);
  and (_09077_, _09076_, _09070_);
  and (_09078_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_09079_, _26133_, _25279_);
  or (_09080_, _09079_, _09078_);
  or (_09082_, _09080_, _09077_);
  and (_02990_, _09082_, _23049_);
  and (_09084_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_09085_, _09047_, _25927_);
  or (_27160_, _09085_, _09084_);
  and (_09087_, _26260_, _26190_);
  not (_09089_, _09087_);
  and (_09090_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_09092_, _09087_, _26242_);
  or (_03019_, _09092_, _09090_);
  and (_09094_, _04175_, _26242_);
  and (_09095_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_27115_, _09095_, _09094_);
  and (_09097_, _04175_, _26185_);
  and (_09098_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_03030_, _09098_, _09097_);
  and (_09100_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_09102_, _09087_, _26170_);
  or (_03061_, _09102_, _09100_);
  and (_09103_, _26260_, _25914_);
  not (_09104_, _09103_);
  and (_09106_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  and (_09107_, _09103_, _26185_);
  or (_03064_, _09107_, _09106_);
  and (_09110_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  and (_09111_, _09103_, _23830_);
  or (_03070_, _09111_, _09110_);
  and (_09112_, _04175_, _26085_);
  and (_09113_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_03072_, _09113_, _09112_);
  and (_09114_, _04175_, _23830_);
  and (_09115_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_03076_, _09115_, _09114_);
  and (_09116_, _02484_, _23830_);
  and (_09117_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_03081_, _09117_, _09116_);
  and (_09118_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  and (_09119_, _09103_, _23768_);
  or (_03083_, _09119_, _09118_);
  and (_09120_, _26351_, _25886_);
  and (_09121_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_27274_, _09121_, _09120_);
  and (_09122_, _04157_, _26202_);
  and (_09123_, _09122_, _23830_);
  not (_09124_, _09122_);
  and (_09125_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_03111_, _09125_, _09123_);
  and (_09126_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_09127_, _04300_, _26185_);
  or (_03112_, _09127_, _09126_);
  and (_09128_, _04157_, _23220_);
  and (_09129_, _09128_, _23830_);
  not (_09130_, _09128_);
  and (_09131_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or (_03128_, _09131_, _09129_);
  and (_09132_, _08289_, _23768_);
  and (_09133_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_03134_, _09133_, _09132_);
  and (_09134_, _08289_, _26170_);
  and (_09135_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or (_03141_, _09135_, _09134_);
  and (_09136_, _09128_, _23768_);
  and (_09137_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  or (_03143_, _09137_, _09136_);
  and (_09138_, _05551_, _25927_);
  and (_09139_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_03150_, _09139_, _09138_);
  and (_09140_, _04157_, _26072_);
  and (_09141_, _09140_, _26085_);
  not (_09142_, _09140_);
  and (_09143_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or (_03160_, _09143_, _09141_);
  and (_09144_, _09140_, _26170_);
  and (_09146_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or (_03171_, _09146_, _09144_);
  and (_09148_, _08289_, _25927_);
  and (_09149_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or (_03177_, _09149_, _09148_);
  and (_09150_, _05551_, _23768_);
  and (_09151_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_03179_, _09151_, _09150_);
  and (_09152_, _04157_, _25932_);
  and (_09153_, _09152_, _26242_);
  not (_09154_, _09152_);
  and (_09155_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_27155_, _09155_, _09153_);
  and (_09156_, _09152_, _25886_);
  and (_09158_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_03194_, _09158_, _09156_);
  nand (_09159_, _00190_, _25417_);
  and (_09160_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_09161_, _00216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_09162_, _00222_, _00196_);
  and (_09163_, _09162_, _09161_);
  and (_09164_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_09165_, _09164_, _09163_);
  nor (_09166_, _09165_, _00226_);
  or (_09167_, _09166_, _00190_);
  or (_09168_, _09167_, _09160_);
  and (_09169_, _09168_, _23049_);
  and (_03205_, _09169_, _09159_);
  and (_09170_, _04157_, _26150_);
  and (_09171_, _09170_, _26185_);
  not (_09172_, _09170_);
  and (_09173_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or (_03212_, _09173_, _09171_);
  and (_03215_, t0_i, _23049_);
  and (_09174_, _09170_, _25927_);
  and (_09175_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or (_03224_, _09175_, _09174_);
  and (_09176_, _04157_, _26224_);
  and (_09177_, _09176_, _26242_);
  not (_09178_, _09176_);
  and (_09179_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_03228_, _09179_, _09177_);
  and (_09180_, _09176_, _26170_);
  and (_09181_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_03236_, _09181_, _09180_);
  and (_09182_, _04157_, _26283_);
  and (_09184_, _09182_, _26185_);
  not (_09186_, _09182_);
  and (_09187_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or (_03244_, _09187_, _09184_);
  and (_09188_, _09182_, _23830_);
  and (_09189_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or (_03254_, _09189_, _09188_);
  and (_09190_, _09182_, _23768_);
  and (_09191_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  or (_27146_, _09191_, _09190_);
  and (_09192_, _05826_, _26242_);
  and (_09193_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_03271_, _09193_, _09192_);
  and (_09194_, _05826_, _26085_);
  and (_09195_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_03274_, _09195_, _09194_);
  and (_09196_, _04175_, _25886_);
  and (_09197_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_03276_, _09197_, _09196_);
  and (_09198_, _07645_, _25886_);
  and (_09199_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_03280_, _09199_, _09198_);
  and (_09200_, _04175_, _26170_);
  and (_09201_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_03285_, _09201_, _09200_);
  and (_09202_, _05771_, _25927_);
  and (_09203_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  or (_03295_, _09203_, _09202_);
  and (_09204_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_09205_, _26413_, _26185_);
  or (_03298_, _09205_, _09204_);
  and (_09206_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_09207_, _09047_, _25886_);
  or (_03303_, _09207_, _09206_);
  and (_09208_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_09209_, _09087_, _23830_);
  or (_03321_, _09209_, _09208_);
  and (_09211_, _09122_, _26185_);
  and (_09212_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_27158_, _09212_, _09211_);
  and (_09213_, _02484_, _25886_);
  and (_09214_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_03344_, _09214_, _09213_);
  and (_09215_, _09122_, _25927_);
  and (_09216_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_27157_, _09216_, _09215_);
  and (_09217_, _09128_, _26185_);
  and (_09218_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  or (_03348_, _09218_, _09217_);
  and (_09220_, _09128_, _26170_);
  and (_09221_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  or (_03350_, _09221_, _09220_);
  and (_09222_, _09140_, _26242_);
  and (_09223_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  or (_03352_, _09223_, _09222_);
  and (_09224_, _26273_, _26224_);
  and (_09225_, _09224_, _23830_);
  not (_09226_, _09224_);
  and (_09227_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_03362_, _09227_, _09225_);
  and (_09228_, _26374_, _26193_);
  and (_09229_, _09228_, _25886_);
  not (_09230_, _09228_);
  and (_09231_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_03366_, _09231_, _09229_);
  and (_09232_, _09152_, _23768_);
  and (_09233_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_03369_, _09233_, _09232_);
  and (_09234_, _09228_, _26170_);
  and (_09235_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_03373_, _09235_, _09234_);
  and (_09236_, _09170_, _25886_);
  and (_09237_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or (_27149_, _09237_, _09236_);
  and (_09239_, _09176_, _23830_);
  and (_09240_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_03399_, _09240_, _09239_);
  and (_09241_, _09228_, _25927_);
  and (_09242_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_03412_, _09242_, _09241_);
  and (_09244_, _07645_, _23768_);
  and (_09245_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_03417_, _09245_, _09244_);
  and (_09246_, _05771_, _25886_);
  and (_09247_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  or (_03420_, _09247_, _09246_);
  and (_09248_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_09249_, _09047_, _26242_);
  or (_03426_, _09249_, _09248_);
  and (_09250_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_09251_, _09087_, _23768_);
  or (_03435_, _09251_, _09250_);
  and (_09252_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  and (_09253_, _09103_, _25927_);
  or (_03445_, _09253_, _09252_);
  and (_09254_, _09140_, _25886_);
  and (_09255_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or (_03451_, _09255_, _09254_);
  and (_09256_, _09152_, _23830_);
  and (_09257_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_27154_, _09257_, _09256_);
  and (_09258_, _09170_, _26242_);
  and (_09259_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or (_03454_, _09259_, _09258_);
  and (_09260_, _09176_, _23768_);
  and (_09261_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_03460_, _09261_, _09260_);
  and (_09262_, _09182_, _25927_);
  and (_09263_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  or (_03466_, _09263_, _09262_);
  and (_09264_, _07645_, _23830_);
  and (_09265_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_03470_, _09265_, _09264_);
  and (_09266_, _05771_, _26085_);
  and (_09267_, _05773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or (_03473_, _09267_, _09266_);
  and (_09268_, _09122_, _26170_);
  and (_09269_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_03482_, _09269_, _09268_);
  and (_09270_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  and (_09271_, _26214_, _26170_);
  or (_03503_, _09271_, _09270_);
  and (_09272_, _07645_, _26085_);
  and (_09273_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_03506_, _09273_, _09272_);
  and (_09274_, _04812_, _26185_);
  and (_09275_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_03508_, _09275_, _09274_);
  and (_09276_, _09228_, _26185_);
  and (_09277_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_03510_, _09277_, _09276_);
  and (_09278_, _04812_, _23768_);
  and (_09279_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_03512_, _09279_, _09278_);
  and (_09280_, _02484_, _26085_);
  and (_09281_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_03516_, _09281_, _09280_);
  and (_09282_, _09228_, _26085_);
  and (_09283_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_03525_, _09283_, _09282_);
  and (_09284_, _03124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_09285_, _09284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_09286_, _09285_, _00221_);
  and (_09287_, _02638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or (_09288_, _09287_, _09286_);
  and (_09289_, _09288_, _00195_);
  or (_09290_, _09287_, _09285_);
  and (_09291_, _09290_, _02356_);
  nand (_09292_, _00209_, _00192_);
  and (_09293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_09294_, _09293_, _09292_);
  or (_09295_, _09294_, _00223_);
  or (_09296_, _09295_, _09291_);
  or (_09297_, _09296_, _09289_);
  and (_09298_, _09297_, _23049_);
  and (_03529_, _09298_, _02363_);
  and (_09299_, _09228_, _23830_);
  and (_09300_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_03531_, _09300_, _09299_);
  and (_09301_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_09302_, _26422_, _26170_);
  or (_03553_, _09302_, _09301_);
  and (_09304_, _26150_, _23779_);
  not (_09305_, _09304_);
  and (_09306_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_09307_, _09304_, _23830_);
  or (_03556_, _09307_, _09306_);
  nand (_09308_, _00071_, _25417_);
  and (_09309_, _01654_, _01666_);
  and (_09310_, _01669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_09311_, _09310_, _01658_);
  and (_09312_, _09311_, _09309_);
  and (_09313_, _09312_, _00083_);
  and (_09314_, _09313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_09315_, _09314_);
  and (_09316_, _09315_, _01673_);
  and (_09317_, _00084_, _00072_);
  nor (_09318_, _09317_, _01674_);
  or (_09319_, _09318_, _09316_);
  and (_09320_, _09319_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_09321_, _02497_, _00084_);
  or (_09322_, _09321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_09323_, _02498_, _02503_);
  and (_09324_, _09323_, _09322_);
  and (_09325_, _09314_, _01673_);
  and (_09326_, _09317_, _00074_);
  nor (_09327_, _09326_, _09325_);
  nor (_09328_, _09327_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_09330_, _09328_, _09324_);
  or (_09331_, _09330_, _09320_);
  or (_09332_, _09331_, _00071_);
  and (_09333_, _09332_, _00070_);
  and (_09334_, _09333_, _09308_);
  and (_09335_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_09336_, _09335_, _09334_);
  and (_03559_, _09336_, _23049_);
  nand (_09337_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_09338_, _09337_, _25891_);
  or (_09339_, _09338_, _00244_);
  and (_09340_, _26090_, _05639_);
  or (_09341_, _09340_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_09342_, _09341_, _25891_);
  and (_09343_, _09342_, _09339_);
  or (_09344_, _09343_, _25903_);
  nand (_09345_, _25903_, _25332_);
  and (_09346_, _09345_, _23049_);
  and (_03566_, _09346_, _09344_);
  and (_09347_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_09348_, _26413_, _26170_);
  or (_27069_, _09348_, _09347_);
  nor (_09349_, _26133_, _25332_);
  not (_09350_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_09351_, _26096_, _09350_);
  nand (_09352_, _09351_, _26120_);
  and (_09353_, _26109_, _26104_);
  or (_09354_, _09353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_09355_, _09354_, _05574_);
  and (_09356_, _09355_, _26095_);
  nand (_09357_, _09356_, _09352_);
  and (_09358_, _26093_, _09350_);
  nor (_09360_, _09358_, _09072_);
  and (_09361_, _09360_, _09357_);
  and (_09362_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_09363_, _09362_, _09361_);
  or (_09364_, _09363_, _09349_);
  and (_03574_, _09364_, _23049_);
  and (_09365_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  and (_09366_, _26214_, _23830_);
  or (_03577_, _09366_, _09365_);
  and (_09367_, _05551_, _26085_);
  and (_09368_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_03585_, _09368_, _09367_);
  and (_09369_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  and (_09370_, _00418_, _26185_);
  or (_03587_, _09370_, _09369_);
  and (_09371_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_09372_, _09371_, _26120_);
  nand (_09373_, _26114_, _26104_);
  nor (_09374_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_09375_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_09376_, _09375_, _26093_);
  or (_09377_, _09376_, _09374_);
  or (_09378_, _09377_, _09372_);
  nor (_09379_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_09380_, _09379_, _09072_);
  and (_09381_, _09380_, _09378_);
  and (_09382_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_09383_, _26142_, _25160_);
  or (_09384_, _09383_, _09382_);
  or (_09385_, _09384_, _09381_);
  and (_03589_, _09385_, _23049_);
  and (_09386_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_09387_, _09386_, _26120_);
  and (_09388_, _26111_, _26104_);
  or (_09389_, _09388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_09390_, _09388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_09391_, _09390_, _09389_);
  or (_09392_, _09391_, _26093_);
  or (_09393_, _09392_, _09387_);
  nor (_09394_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_09395_, _09394_, _09072_);
  and (_09396_, _09395_, _09393_);
  and (_09397_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_09398_, _26138_, _25283_);
  or (_09399_, _09398_, _09397_);
  or (_09400_, _09399_, _09396_);
  and (_03595_, _09400_, _23049_);
  and (_09401_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_09402_, _26321_, _26085_);
  or (_03600_, _09402_, _09401_);
  and (_09403_, _26322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_09404_, _26321_, _23768_);
  or (_03602_, _09404_, _09403_);
  and (_09405_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_09406_, _26417_, _25886_);
  or (_03605_, _09406_, _09405_);
  and (_09407_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_09408_, _00059_, _23830_);
  or (_03610_, _09408_, _09407_);
  and (_09409_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_09410_, _00141_, _23768_);
  or (_03613_, _09410_, _09409_);
  and (_09411_, _25891_, _25224_);
  nand (_09412_, _09411_, _23729_);
  or (_09413_, _09411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_09414_, _09413_, _25910_);
  and (_09415_, _09414_, _09412_);
  nor (_09416_, _25910_, _25279_);
  or (_09417_, _09416_, _09415_);
  and (_03615_, _09417_, _23049_);
  and (_09418_, _26193_, _23775_);
  and (_09419_, _09418_, _26085_);
  not (_09420_, _09418_);
  and (_09421_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_03617_, _09421_, _09419_);
  and (_09422_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_09423_, _02296_, _25927_);
  or (_03626_, _09423_, _09422_);
  and (_09424_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_09425_, _02564_, _23830_);
  or (_03629_, _09425_, _09424_);
  and (_09427_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_09428_, _02564_, _23768_);
  or (_03632_, _09428_, _09427_);
  and (_09431_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_09432_, _02615_, _23768_);
  or (_03641_, _09432_, _09431_);
  and (_09434_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  and (_09435_, _02019_, _26185_);
  or (_03667_, _09435_, _09434_);
  and (_09437_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_09438_, _04004_, _26242_);
  or (_03670_, _09438_, _09437_);
  and (_09439_, _05551_, _23830_);
  and (_09440_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_03673_, _09440_, _09439_);
  and (_09441_, _04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_09442_, _04004_, _25886_);
  or (_03676_, _09442_, _09441_);
  and (_09444_, _05551_, _25886_);
  and (_09446_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_03680_, _09446_, _09444_);
  and (_09448_, _09418_, _23830_);
  and (_09449_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_03682_, _09449_, _09448_);
  and (_09450_, _26072_, _23779_);
  not (_09451_, _09450_);
  and (_09452_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_09453_, _09450_, _26185_);
  or (_03692_, _09453_, _09452_);
  and (_09454_, _09228_, _23768_);
  and (_09455_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_03720_, _09455_, _09454_);
  and (_09456_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_09457_, _26185_, _25915_);
  or (_03727_, _09457_, _09456_);
  and (_09459_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_09460_, _04016_, _23768_);
  or (_03738_, _09460_, _09459_);
  and (_09461_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_09462_, _02296_, _26185_);
  or (_03743_, _09462_, _09461_);
  and (_09463_, _09418_, _26242_);
  and (_09464_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_03745_, _09464_, _09463_);
  and (_09465_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_09466_, _02615_, _26085_);
  or (_03749_, _09466_, _09465_);
  and (_09467_, _02826_, _25886_);
  and (_09468_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_03763_, _09468_, _09467_);
  and (_09469_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_09470_, _26602_, _25927_);
  or (_03765_, _09470_, _09469_);
  and (_09471_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_09472_, _02879_, _25886_);
  or (_27053_, _09472_, _09471_);
  and (_09473_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_09474_, _04820_, _26170_);
  or (_03782_, _09474_, _09473_);
  and (_09475_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_09476_, _26413_, _25886_);
  or (_03785_, _09476_, _09475_);
  and (_09477_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_09478_, _02564_, _26085_);
  or (_03794_, _09478_, _09477_);
  and (_09479_, _04223_, _25927_);
  and (_09480_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_03826_, _09480_, _09479_);
  and (_09481_, _04223_, _23768_);
  and (_09483_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_03844_, _09483_, _09481_);
  and (_09484_, _04157_, _23775_);
  and (_09485_, _09484_, _23830_);
  not (_09486_, _09484_);
  and (_09487_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or (_03850_, _09487_, _09485_);
  and (_09488_, _09484_, _25927_);
  and (_09489_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  or (_03857_, _09489_, _09488_);
  and (_09490_, _04157_, _26213_);
  and (_09491_, _09490_, _26085_);
  not (_09492_, _09490_);
  and (_09493_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_03866_, _09493_, _09491_);
  and (_09494_, _09490_, _23768_);
  and (_09495_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_27133_, _09495_, _09494_);
  and (_09496_, _04157_, _26190_);
  and (_09497_, _09496_, _26242_);
  not (_09498_, _09496_);
  and (_09499_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_03883_, _09499_, _09497_);
  and (_09500_, _09496_, _26085_);
  and (_09501_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_03886_, _09501_, _09500_);
  and (_09502_, _09496_, _23768_);
  and (_09503_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_03894_, _09503_, _09502_);
  and (_09504_, _26275_, _25886_);
  and (_09505_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_03901_, _09505_, _09504_);
  and (_09506_, _04157_, _25914_);
  and (_09507_, _09506_, _26170_);
  not (_09508_, _09506_);
  and (_09509_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or (_03903_, _09509_, _09507_);
  and (_09510_, _26202_, _26193_);
  and (_09511_, _09510_, _23830_);
  not (_09512_, _09510_);
  and (_09513_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or (_03921_, _09513_, _09511_);
  and (_09514_, _09510_, _26170_);
  and (_09515_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or (_03923_, _09515_, _09514_);
  and (_09516_, _04223_, _25886_);
  and (_09517_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_27112_, _09517_, _09516_);
  and (_09518_, _26193_, _23220_);
  and (_09519_, _09518_, _26242_);
  not (_09521_, _09518_);
  and (_09522_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_03937_, _09522_, _09519_);
  and (_09523_, _09518_, _23830_);
  and (_09524_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_03942_, _09524_, _09523_);
  and (_09525_, _04223_, _26170_);
  and (_09526_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_27111_, _09526_, _09525_);
  and (_09527_, _09518_, _25927_);
  and (_09528_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_27127_, _09528_, _09527_);
  and (_09529_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_09531_, _09304_, _26185_);
  or (_03953_, _09531_, _09529_);
  and (_09532_, _26193_, _25932_);
  and (_09533_, _09532_, _25927_);
  not (_09534_, _09532_);
  and (_09535_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_03959_, _09535_, _09533_);
  and (_09536_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  and (_09537_, _00418_, _25886_);
  or (_03971_, _09537_, _09536_);
  and (_09538_, _26340_, _26193_);
  and (_09539_, _09538_, _25886_);
  not (_09540_, _09538_);
  and (_09541_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_03972_, _09541_, _09539_);
  and (_09542_, _09538_, _25927_);
  and (_09543_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or (_03973_, _09543_, _09542_);
  and (_09544_, _26421_, _26193_);
  and (_09545_, _09544_, _26185_);
  not (_09546_, _09544_);
  and (_09547_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_27124_, _09547_, _09545_);
  and (_09548_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  and (_09549_, _26214_, _23768_);
  or (_03978_, _09549_, _09548_);
  and (_09550_, _07645_, _26170_);
  and (_09551_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_03979_, _09551_, _09550_);
  and (_09552_, _09544_, _25927_);
  and (_09553_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_03980_, _09553_, _09552_);
  and (_09554_, _04915_, _26085_);
  and (_09555_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_27122_, _09555_, _09554_);
  and (_09556_, _09224_, _26185_);
  and (_09557_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_03992_, _09557_, _09556_);
  and (_09558_, _26193_, _26072_);
  and (_09559_, _09558_, _26170_);
  not (_09560_, _09558_);
  and (_09561_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_03996_, _09561_, _09559_);
  and (_09562_, _09558_, _23768_);
  and (_09563_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_03998_, _09563_, _09562_);
  and (_09564_, _09532_, _26242_);
  and (_09565_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_04006_, _09565_, _09564_);
  and (_09566_, _02825_, _26190_);
  and (_09567_, _09566_, _26185_);
  not (_09568_, _09566_);
  and (_09569_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_04009_, _09569_, _09567_);
  and (_09570_, _09532_, _23830_);
  and (_09571_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_04011_, _09571_, _09570_);
  and (_09572_, _26301_, _26085_);
  and (_09573_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_04013_, _09573_, _09572_);
  and (_09574_, _09566_, _26085_);
  and (_09575_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_04021_, _09575_, _09574_);
  and (_09576_, _09490_, _26242_);
  and (_09577_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_04023_, _09577_, _09576_);
  and (_09578_, _09224_, _26085_);
  and (_09579_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_04028_, _09579_, _09578_);
  and (_09580_, _09496_, _26170_);
  and (_09581_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_04034_, _09581_, _09580_);
  and (_09583_, _09506_, _26242_);
  and (_09584_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  or (_04036_, _09584_, _09583_);
  and (_09586_, _09506_, _23830_);
  and (_09587_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or (_04039_, _09587_, _09586_);
  and (_09588_, _09510_, _26185_);
  and (_09589_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_04043_, _09589_, _09588_);
  and (_09592_, _05826_, _25886_);
  and (_09593_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_04046_, _09593_, _09592_);
  and (_09594_, _09544_, _25886_);
  and (_09595_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_27123_, _09595_, _09594_);
  and (_09596_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_09597_, _26085_, _23780_);
  or (_04073_, _09597_, _09596_);
  and (_09598_, _26615_, _26085_);
  and (_09599_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_04082_, _09599_, _09598_);
  and (_09600_, _02825_, _26283_);
  and (_09601_, _09600_, _26170_);
  not (_09603_, _09600_);
  and (_09605_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or (_04088_, _09605_, _09601_);
  and (_09606_, _09490_, _25927_);
  and (_09608_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_04099_, _09608_, _09606_);
  and (_09610_, _02825_, _23847_);
  and (_09611_, _09610_, _25886_);
  not (_09612_, _09610_);
  and (_09614_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_04102_, _09614_, _09611_);
  and (_09616_, _09610_, _26085_);
  and (_09618_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_04104_, _09618_, _09616_);
  and (_09619_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_09620_, _04300_, _23830_);
  or (_04109_, _09620_, _09619_);
  and (_09621_, _09610_, _26242_);
  and (_09622_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_04110_, _09622_, _09621_);
  and (_09623_, _26275_, _23830_);
  and (_09624_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_04115_, _09624_, _09623_);
  and (_09625_, _23961_, _23935_);
  or (_09627_, _24065_, _09625_);
  and (_09628_, _23947_, _24049_);
  and (_09629_, _23977_, _09628_);
  and (_09631_, _23928_, _22909_);
  and (_09632_, _09631_, _22934_);
  and (_09633_, _24004_, _09632_);
  or (_09634_, _09633_, _09629_);
  nor (_09635_, _09634_, _09627_);
  nand (_09637_, _09635_, _23985_);
  or (_09639_, _24030_, _24012_);
  or (_09641_, _09639_, _09637_);
  and (_09642_, _24005_, _23998_);
  and (_09643_, _24043_, _23943_);
  or (_09644_, _09643_, _09642_);
  and (_09645_, _23966_, _23946_);
  and (_09646_, _24005_, _09645_);
  and (_09647_, _09632_, _23923_);
  or (_09648_, _09647_, _09646_);
  or (_09649_, _09648_, _09644_);
  or (_09650_, _24042_, _24018_);
  not (_09651_, _23931_);
  nand (_09652_, _24080_, _09651_);
  or (_09654_, _09652_, _09650_);
  or (_09656_, _09654_, _09649_);
  or (_09657_, _09656_, _09641_);
  and (_09658_, _09657_, _22740_);
  and (_09659_, _22737_, _22734_);
  and (_09661_, _09659_, _22942_);
  nor (_09663_, _09661_, _08646_);
  or (_09664_, _09663_, rst);
  or (_26895_[1], _09664_, _09658_);
  and (_09665_, _09558_, _23830_);
  and (_09666_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_04124_, _09666_, _09665_);
  and (_09667_, _02825_, _26213_);
  and (_09668_, _09667_, _26242_);
  not (_09669_, _09667_);
  and (_09670_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_27030_, _09670_, _09668_);
  and (_09672_, _02825_, _23775_);
  and (_09673_, _09672_, _23768_);
  not (_09675_, _09672_);
  and (_09676_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or (_04133_, _09676_, _09673_);
  and (_09679_, _00068_, _25900_);
  nand (_09680_, _09679_, _25362_);
  and (_09682_, _00189_, _25900_);
  not (_09684_, _09682_);
  not (_09685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_09686_, _26096_, _26090_);
  nor (_09687_, _09686_, _09685_);
  and (_09688_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_09689_, _09688_, _09687_);
  or (_09690_, _09679_, _09689_);
  and (_09691_, _09690_, _09684_);
  and (_09692_, _09691_, _09680_);
  and (_09693_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_09694_, _09693_, _09692_);
  and (_04144_, _09694_, _23049_);
  and (_09696_, _09672_, _26170_);
  and (_09697_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or (_27031_, _09697_, _09696_);
  and (_09698_, _09672_, _25886_);
  and (_09700_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or (_04154_, _09700_, _09698_);
  and (_09702_, _09672_, _26185_);
  and (_09704_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or (_04158_, _09704_, _09702_);
  and (_09705_, _09532_, _26085_);
  and (_09706_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_04168_, _09706_, _09705_);
  and (_09707_, _09672_, _26242_);
  and (_09709_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or (_04171_, _09709_, _09707_);
  not (_09711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_09712_, _09686_, _09711_);
  and (_09713_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_09714_, _09713_, _09712_);
  or (_09715_, _09714_, _09679_);
  nand (_09716_, _09679_, _23761_);
  and (_09718_, _09716_, _09715_);
  or (_09719_, _09718_, _09682_);
  nand (_09720_, _09682_, _09711_);
  and (_09721_, _09720_, _23049_);
  and (_04173_, _09721_, _09719_);
  nand (_09722_, _09682_, _25160_);
  not (_09723_, _09686_);
  nor (_09724_, _09679_, _09723_);
  not (_09725_, _09724_);
  and (_09726_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_09728_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_09729_, _09728_, _09726_);
  or (_09730_, _09729_, _09682_);
  and (_09731_, _09730_, _23049_);
  and (_04174_, _09731_, _09722_);
  and (_09732_, _02825_, _26374_);
  and (_09733_, _09732_, _25927_);
  not (_09734_, _09732_);
  and (_09735_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or (_04178_, _09735_, _09733_);
  or (_09736_, _26104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_09737_, _26096_, _09711_);
  and (_09739_, _09737_, _26119_);
  or (_09741_, _09739_, _09066_);
  and (_09742_, _09741_, _09736_);
  or (_09743_, _09742_, _26093_);
  nand (_09744_, _26093_, _09711_);
  and (_09746_, _09744_, _05563_);
  and (_09748_, _09746_, _09743_);
  and (_09750_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_09752_, _26132_, _25283_);
  or (_09754_, _09752_, _09750_);
  or (_09755_, _09754_, _09748_);
  and (_04180_, _09755_, _23049_);
  and (_09756_, _25914_, _23230_);
  and (_09757_, _09756_, _26085_);
  not (_09758_, _09756_);
  and (_09759_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_04183_, _09759_, _09757_);
  and (_09760_, _09532_, _26170_);
  and (_09761_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or (_27126_, _09761_, _09760_);
  and (_09762_, _09732_, _26170_);
  and (_09763_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or (_04186_, _09763_, _09762_);
  and (_09765_, _09732_, _26085_);
  and (_09766_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or (_04188_, _09766_, _09765_);
  and (_09769_, _04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_09770_, _04016_, _26185_);
  or (_04191_, _09770_, _09769_);
  and (_09771_, _09532_, _25886_);
  and (_09772_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or (_04193_, _09772_, _09771_);
  and (_09773_, _09532_, _26185_);
  and (_09775_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_04213_, _09775_, _09773_);
  and (_09776_, _09732_, _26185_);
  and (_09777_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or (_04216_, _09777_, _09776_);
  and (_09780_, _02825_, _26258_);
  and (_09781_, _09780_, _23768_);
  not (_09782_, _09780_);
  and (_09784_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_04220_, _09784_, _09781_);
  and (_09786_, _00095_, _23220_);
  and (_09787_, _09786_, _25927_);
  not (_09788_, _09786_);
  and (_09789_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_04225_, _09789_, _09787_);
  and (_09791_, _00095_, _26072_);
  and (_09792_, _09791_, _25886_);
  not (_09793_, _09791_);
  and (_09794_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_04229_, _09794_, _09792_);
  and (_09795_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_09796_, _02879_, _26170_);
  or (_04238_, _09796_, _09795_);
  and (_09797_, _09780_, _25927_);
  and (_09798_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_04239_, _09798_, _09797_);
  and (_09799_, _09780_, _23830_);
  and (_09800_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_04242_, _09800_, _09799_);
  and (_09801_, _07104_, _26170_);
  and (_09803_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_04244_, _09803_, _09801_);
  and (_09804_, _02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_09805_, _02879_, _26085_);
  or (_27054_, _09805_, _09804_);
  and (_09806_, _09558_, _25927_);
  and (_09807_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_04253_, _09807_, _09806_);
  and (_09808_, _09558_, _25886_);
  and (_09809_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_04258_, _09809_, _09808_);
  and (_09810_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_09811_, _26602_, _23768_);
  or (_04260_, _09811_, _09810_);
  and (_09813_, _04915_, _25886_);
  and (_09814_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_04264_, _09814_, _09813_);
  and (_09815_, _09780_, _26085_);
  and (_09816_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_04266_, _09816_, _09815_);
  and (_09817_, _09780_, _26242_);
  and (_09818_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_04268_, _09818_, _09817_);
  and (_09819_, _02849_, _26242_);
  and (_09820_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or (_04270_, _09820_, _09819_);
  and (_09821_, _07104_, _23830_);
  and (_09822_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_27215_, _09822_, _09821_);
  and (_09823_, _09610_, _23768_);
  and (_09824_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_04276_, _09824_, _09823_);
  and (_09825_, _09600_, _23830_);
  and (_09826_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or (_04279_, _09826_, _09825_);
  and (_09827_, _02849_, _26085_);
  and (_09829_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or (_04285_, _09829_, _09827_);
  and (_09831_, _02826_, _26170_);
  and (_09832_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_04289_, _09832_, _09831_);
  and (_09835_, _04915_, _23830_);
  and (_09836_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_27121_, _09836_, _09835_);
  and (_09837_, _09224_, _25927_);
  and (_09838_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_04293_, _09838_, _09837_);
  and (_09839_, _04915_, _26185_);
  and (_09840_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_04310_, _09840_, _09839_);
  and (_09841_, _02826_, _26085_);
  and (_09842_, _02828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_04312_, _09842_, _09841_);
  and (_09844_, _09600_, _26085_);
  and (_09845_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or (_04315_, _09845_, _09844_);
  and (_09846_, _09600_, _26242_);
  and (_09847_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or (_04317_, _09847_, _09846_);
  and (_09849_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and (_09851_, _02792_, _26170_);
  or (_04320_, _09851_, _09849_);
  and (_09852_, _02825_, _26224_);
  and (_09854_, _09852_, _23768_);
  not (_09855_, _09852_);
  and (_09856_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_04324_, _09856_, _09854_);
  and (_09857_, _09852_, _25886_);
  and (_09858_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_04326_, _09858_, _09857_);
  and (_09859_, _07104_, _25886_);
  and (_09860_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_04328_, _09860_, _09859_);
  and (_09861_, _04915_, _26242_);
  and (_09862_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_04331_, _09862_, _09861_);
  and (_09863_, _02793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_09864_, _02792_, _23768_);
  or (_04336_, _09864_, _09863_);
  and (_09865_, _09852_, _23830_);
  and (_09866_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_04346_, _09866_, _09865_);
  and (_09867_, _09544_, _23768_);
  and (_09868_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_04354_, _09868_, _09867_);
  and (_09869_, _09852_, _26185_);
  and (_09870_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_04358_, _09870_, _09869_);
  and (_09871_, _09544_, _26170_);
  and (_09872_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_04361_, _09872_, _09871_);
  and (_09873_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_09874_, _02615_, _23830_);
  or (_04365_, _09874_, _09873_);
  and (_09876_, _09544_, _23830_);
  and (_09877_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_04371_, _09877_, _09876_);
  and (_09879_, _02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_09881_, _02615_, _26242_);
  or (_04380_, _09881_, _09879_);
  and (_09882_, _09544_, _26085_);
  and (_09883_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_04386_, _09883_, _09882_);
  and (_09884_, _02565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_09885_, _02564_, _26170_);
  or (_27047_, _09885_, _09884_);
  and (_09886_, _02825_, _26150_);
  and (_09887_, _09886_, _25927_);
  not (_09888_, _09886_);
  and (_09889_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or (_04393_, _09889_, _09887_);
  and (_09890_, _09886_, _25886_);
  and (_09891_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or (_04396_, _09891_, _09890_);
  and (_09892_, _09544_, _26242_);
  and (_09893_, _09546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_04419_, _09893_, _09892_);
  and (_09894_, _09886_, _23830_);
  and (_09895_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or (_04423_, _09895_, _09894_);
  and (_09896_, _09886_, _26185_);
  and (_09897_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or (_04426_, _09897_, _09896_);
  and (_09898_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_09899_, _02296_, _26085_);
  or (_04429_, _09899_, _09898_);
  and (_09900_, _09538_, _23768_);
  and (_09901_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_04435_, _09901_, _09900_);
  and (_09903_, _02825_, _26421_);
  and (_09904_, _09903_, _23768_);
  not (_09905_, _09903_);
  and (_09906_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or (_04439_, _09906_, _09904_);
  and (_09908_, _02297_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_09909_, _02296_, _25886_);
  or (_04442_, _09909_, _09908_);
  and (_09911_, _09224_, _25886_);
  and (_09913_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_04447_, _09913_, _09911_);
  and (_09914_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and (_09915_, _01962_, _25927_);
  or (_04450_, _09915_, _09914_);
  and (_09916_, _09538_, _26170_);
  and (_09917_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_04452_, _09917_, _09916_);
  and (_09918_, _09903_, _25927_);
  and (_09919_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or (_04456_, _09919_, _09918_);
  and (_09921_, _09538_, _23830_);
  and (_09922_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or (_04461_, _09922_, _09921_);
  and (_09923_, _01963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and (_09924_, _01962_, _26085_);
  or (_04466_, _09924_, _09923_);
  and (_09926_, _09903_, _25886_);
  and (_09928_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or (_04469_, _09928_, _09926_);
  and (_09931_, _00142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_09932_, _00141_, _26185_);
  or (_04473_, _09932_, _09931_);
  and (_09933_, _09538_, _26085_);
  and (_09935_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_04478_, _09935_, _09933_);
  and (_09936_, _09903_, _26085_);
  and (_09937_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or (_04486_, _09937_, _09936_);
  and (_09939_, _09538_, _26185_);
  and (_09940_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_27125_, _09940_, _09939_);
  and (_09942_, _00060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_09943_, _00059_, _25927_);
  or (_04493_, _09943_, _09942_);
  and (_09945_, _09791_, _26185_);
  and (_09946_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_04501_, _09946_, _09945_);
  and (_09948_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and (_09950_, _00022_, _25927_);
  or (_04504_, _09950_, _09948_);
  and (_09952_, _09538_, _26242_);
  and (_09954_, _09540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_04518_, _09954_, _09952_);
  and (_09956_, _02825_, _26340_);
  and (_09958_, _09956_, _25927_);
  not (_09960_, _09956_);
  and (_09961_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_04521_, _09961_, _09958_);
  and (_09962_, _09956_, _25886_);
  and (_09963_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_04528_, _09963_, _09962_);
  and (_09964_, _09532_, _23768_);
  and (_09965_, _09534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_04530_, _09965_, _09964_);
  and (_09966_, _07104_, _26242_);
  and (_09967_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_04535_, _09967_, _09966_);
  and (_09968_, _00023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_09970_, _00022_, _23830_);
  or (_04542_, _09970_, _09968_);
  and (_09972_, _09558_, _26085_);
  and (_09973_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_04544_, _09973_, _09972_);
  and (_09975_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_09977_, _26602_, _26185_);
  or (_04549_, _09977_, _09975_);
  and (_09978_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  and (_09979_, _06369_, _26242_);
  or (_04553_, _09979_, _09978_);
  and (_09980_, _09956_, _23830_);
  and (_09981_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_27036_, _09981_, _09980_);
  and (_09982_, _26603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_09983_, _26602_, _23830_);
  or (_04557_, _09983_, _09982_);
  and (_09986_, _09558_, _26185_);
  and (_09987_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_04559_, _09987_, _09986_);
  and (_09988_, _09786_, _26170_);
  and (_09989_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_04563_, _09989_, _09988_);
  and (_09991_, _09956_, _26242_);
  and (_09992_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_04565_, _09992_, _09991_);
  and (_09994_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_09996_, _26417_, _23768_);
  or (_04570_, _09996_, _09994_);
  and (_09998_, _02825_, _25932_);
  and (_09999_, _09998_, _23768_);
  not (_10000_, _09998_);
  and (_10001_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_04574_, _10001_, _09999_);
  and (_10002_, _09558_, _26242_);
  and (_10003_, _09560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_04578_, _10003_, _10002_);
  and (_10004_, _09998_, _26170_);
  and (_10005_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_04583_, _10005_, _10004_);
  and (_10006_, _26418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_10007_, _26417_, _26085_);
  or (_04586_, _10007_, _10006_);
  and (_10010_, _07104_, _26185_);
  and (_10011_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_04589_, _10011_, _10010_);
  and (_10012_, _09518_, _23768_);
  and (_10013_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_04593_, _10013_, _10012_);
  and (_10014_, _09998_, _25886_);
  and (_10015_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_04596_, _10015_, _10014_);
  and (_10016_, _09998_, _26185_);
  and (_10018_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_04599_, _10018_, _10016_);
  and (_10020_, _26255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_10021_, _26254_, _25886_);
  or (_04623_, _10021_, _10020_);
  and (_10024_, _09518_, _26170_);
  and (_10025_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_04625_, _10025_, _10024_);
  and (_10026_, _07104_, _26085_);
  and (_10028_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_04629_, _10028_, _10026_);
  and (_10029_, _02825_, _26072_);
  and (_10030_, _10029_, _25927_);
  not (_10031_, _10029_);
  and (_10032_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or (_27039_, _10032_, _10030_);
  and (_10033_, _10029_, _25886_);
  and (_10034_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or (_04634_, _10034_, _10033_);
  and (_10036_, _26206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_10037_, _26205_, _25927_);
  or (_04636_, _10037_, _10036_);
  and (_10038_, _09518_, _25886_);
  and (_10039_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_04639_, _10039_, _10038_);
  and (_10041_, _09518_, _26085_);
  and (_10042_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_04646_, _10042_, _10041_);
  and (_10043_, _10029_, _26085_);
  and (_10044_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or (_04650_, _10044_, _10043_);
  and (_10046_, _00016_, _26170_);
  and (_10047_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_04656_, _10047_, _10046_);
  and (_10049_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_10050_, _26085_, _25915_);
  or (_27061_, _10050_, _10049_);
  and (_10052_, _09518_, _26185_);
  and (_10053_, _09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_04665_, _10053_, _10052_);
  and (_10055_, _09510_, _23768_);
  and (_10056_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_04671_, _10056_, _10055_);
  and (_10057_, _10029_, _26242_);
  and (_10059_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or (_27041_, _10059_, _10057_);
  and (_10060_, _02849_, _23768_);
  and (_10061_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or (_04685_, _10061_, _10060_);
  and (_10063_, _09510_, _25927_);
  and (_10064_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_04689_, _10064_, _10063_);
  and (_10065_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_10066_, _25886_, _23780_);
  or (_04702_, _10066_, _10065_);
  and (_10067_, _09510_, _25886_);
  and (_10069_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or (_27128_, _10069_, _10067_);
  and (_10070_, _09510_, _26085_);
  and (_10072_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_04711_, _10072_, _10070_);
  and (_10073_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_10075_, _26242_, _23780_);
  or (_27066_, _10075_, _10073_);
  and (_10077_, _02849_, _25927_);
  and (_10079_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or (_04729_, _10079_, _10077_);
  and (_10080_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  and (_10082_, _02019_, _26170_);
  or (_04736_, _10082_, _10080_);
  and (_10084_, _09510_, _26242_);
  and (_10085_, _09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_04753_, _10085_, _10084_);
  and (_10086_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_10088_, _26413_, _26242_);
  or (_04756_, _10088_, _10086_);
  and (_10089_, _09506_, _23768_);
  and (_10090_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  or (_04759_, _10090_, _10089_);
  and (_10091_, _09667_, _23768_);
  and (_10092_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_27028_, _10092_, _10091_);
  and (_10093_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  and (_10094_, _02019_, _26242_);
  or (_27072_, _10094_, _10093_);
  and (_10096_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  and (_10097_, _02019_, _26085_);
  or (_04779_, _10097_, _10096_);
  and (_10098_, _04181_, _26185_);
  and (_10100_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or (_04781_, _10100_, _10098_);
  and (_10102_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  and (_10103_, _02010_, _23830_);
  or (_04785_, _10103_, _10102_);
  and (_10104_, _09506_, _25927_);
  and (_10106_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  or (_04788_, _10106_, _10104_);
  and (_10108_, _09566_, _26242_);
  and (_10109_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_04794_, _10109_, _10108_);
  and (_10111_, _09506_, _25886_);
  and (_10112_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or (_04797_, _10112_, _10111_);
  and (_10113_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_10115_, _04820_, _25927_);
  or (_27074_, _10115_, _10113_);
  and (_10118_, _09506_, _26085_);
  and (_10119_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or (_27129_, _10119_, _10118_);
  and (_10120_, _04181_, _26085_);
  and (_10121_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or (_04813_, _10121_, _10120_);
  and (_10122_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  and (_10123_, _02576_, _23768_);
  or (_04816_, _10123_, _10122_);
  and (_10124_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  and (_10126_, _02576_, _26185_);
  or (_04824_, _10126_, _10124_);
  and (_10127_, _09506_, _26185_);
  and (_10128_, _09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or (_04829_, _10128_, _10127_);
  and (_10130_, _09496_, _25927_);
  and (_10132_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_04839_, _10132_, _10130_);
  and (_10134_, _09566_, _25927_);
  and (_10135_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_04842_, _10135_, _10134_);
  and (_10137_, _09224_, _26170_);
  and (_10138_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_04844_, _10138_, _10137_);
  and (_10139_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_10140_, _09304_, _26242_);
  or (_04846_, _10140_, _10139_);
  and (_10143_, _05826_, _23830_);
  and (_10145_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_04864_, _10145_, _10143_);
  and (_10147_, _09496_, _25886_);
  and (_10148_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_04867_, _10148_, _10147_);
  and (_10150_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  and (_10152_, _01996_, _25927_);
  or (_04869_, _10152_, _10150_);
  or (_10155_, _01617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  not (_10156_, _01618_);
  and (_10157_, _10156_, _02554_);
  and (_10158_, _10157_, _10155_);
  and (_10159_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_10160_, _10159_, _10158_);
  and (_10162_, _10160_, _02363_);
  and (_10164_, _01612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_10166_, _10164_, _01627_);
  or (_10167_, _10166_, _10162_);
  nor (_10169_, _01612_, _25160_);
  or (_10170_, _10169_, _10167_);
  and (_04871_, _10170_, _23049_);
  and (_10172_, _09566_, _23768_);
  and (_10173_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_04874_, _10173_, _10172_);
  and (_10175_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_10176_, _26422_, _26185_);
  or (_04877_, _10176_, _10175_);
  and (_10178_, _01625_, _00209_);
  or (_10180_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_10183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand (_10184_, _10183_, _02531_);
  and (_10185_, _10184_, _01614_);
  nand (_10187_, _10185_, _01625_);
  and (_10189_, _10187_, _10180_);
  or (_10190_, _10189_, _00190_);
  nand (_10191_, _00190_, _23761_);
  and (_10192_, _10191_, _23049_);
  and (_04883_, _10192_, _10190_);
  and (_10193_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  and (_10194_, _01996_, _26242_);
  or (_27086_, _10194_, _10193_);
  and (_10196_, _09496_, _23830_);
  and (_10198_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_27130_, _10198_, _10196_);
  and (_10200_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  and (_10201_, _01996_, _23830_);
  or (_27084_, _10201_, _10200_);
  or (_10202_, _00222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_10203_, _02539_, _00221_);
  and (_10204_, _10203_, _00195_);
  and (_10205_, _10204_, _10202_);
  or (_10206_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_10207_, _02539_, _02656_);
  and (_10208_, _10207_, _10206_);
  or (_10209_, _10208_, _10183_);
  nor (_10210_, _10209_, _10205_);
  nand (_10212_, _10210_, _02363_);
  nand (_10213_, _00226_, _23761_);
  or (_10214_, _01612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_10215_, _10214_, _23049_);
  and (_10216_, _10215_, _10213_);
  and (_04891_, _10216_, _10212_);
  and (_10218_, _25932_, _23779_);
  not (_10220_, _10218_);
  and (_10221_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  and (_10222_, _10218_, _26185_);
  or (_27087_, _10222_, _10221_);
  and (_10225_, _07104_, _23768_);
  and (_10226_, _07106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_27214_, _10226_, _10225_);
  and (_10229_, _09496_, _26185_);
  and (_10231_, _09498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_27131_, _10231_, _10229_);
  nor (_10233_, _25858_, _24307_);
  nor (_10235_, _01361_, _01358_);
  nor (_10236_, _10235_, _24307_);
  and (_10237_, _10236_, _22748_);
  nor (_10238_, _10236_, _22748_);
  nor (_10240_, _10238_, _10237_);
  nor (_10242_, _10240_, _10233_);
  and (_10243_, _22750_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_10244_, _10243_, _10233_);
  nor (_10245_, _10244_, _24087_);
  or (_10246_, _10245_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_10248_, _10246_, _10242_);
  and (_26927_[2], _10248_, _23049_);
  and (_10250_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_10251_, _09450_, _26085_);
  or (_27088_, _10251_, _10250_);
  and (_10252_, _04181_, _26242_);
  and (_10254_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or (_27213_, _10254_, _10252_);
  and (_10255_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  and (_10256_, _00089_, _26242_);
  or (_27168_, _10256_, _10255_);
  and (_10257_, _09490_, _26170_);
  and (_10258_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_27134_, _10258_, _10257_);
  and (_10259_, _23779_, _23220_);
  not (_10260_, _10259_);
  and (_10262_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_10264_, _10259_, _23830_);
  or (_27094_, _10264_, _10262_);
  and (_10265_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_10266_, _10259_, _25927_);
  or (_27092_, _10266_, _10265_);
  nand (_10267_, _00069_, _25160_);
  and (_10268_, _05692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_10270_, _05696_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not (_10271_, _00071_);
  nand (_10272_, _05697_, _10271_);
  and (_10273_, _10272_, _10270_);
  or (_10274_, _10273_, _10268_);
  or (_10275_, _10271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_10276_, _10275_, _10274_);
  or (_10278_, _10276_, _00069_);
  and (_10279_, _10278_, _23049_);
  and (_04919_, _10279_, _10267_);
  and (_10281_, _05826_, _26185_);
  and (_10282_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_27145_, _10282_, _10281_);
  and (_10283_, _26202_, _23779_);
  not (_10284_, _10283_);
  and (_10285_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  and (_10286_, _10283_, _26170_);
  or (_27096_, _10286_, _10285_);
  and (_10287_, _09566_, _25886_);
  and (_10288_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_27027_, _10288_, _10287_);
  and (_10289_, _09490_, _25886_);
  and (_10290_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_27135_, _10290_, _10289_);
  or (_10291_, _10271_, _25258_);
  and (_10293_, _02497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_10295_, _10293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_10296_, _10295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_10297_, _10295_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_10298_, _10297_, _02503_);
  and (_10299_, _10297_, _09310_);
  or (_10301_, _09310_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_10303_, _10301_, _01672_);
  nor (_10304_, _10303_, _10299_);
  or (_10305_, _10304_, _10298_);
  and (_10306_, _10305_, _10296_);
  and (_10307_, _00079_, _00072_);
  and (_10308_, _10307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_10309_, _10308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_10311_, _10308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_10312_, _10311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_10313_, _10312_, _10309_);
  or (_10314_, _10313_, _10306_);
  or (_10315_, _10314_, _00071_);
  and (_10316_, _10315_, _00070_);
  and (_10318_, _10316_, _10291_);
  and (_10320_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_10321_, _10320_, _10318_);
  and (_04926_, _10321_, _23049_);
  and (_10324_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  and (_10325_, _10283_, _26242_);
  or (_27099_, _10325_, _10324_);
  and (_10326_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_10327_, _09304_, _26085_);
  or (_27081_, _10327_, _10326_);
  and (_10328_, _09490_, _23830_);
  and (_10329_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_27136_, _10329_, _10328_);
  and (_10330_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  and (_10331_, _10283_, _23830_);
  or (_27098_, _10331_, _10330_);
  and (_10333_, _09490_, _26185_);
  and (_10335_, _09492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_27137_, _10335_, _10333_);
  and (_10336_, _09566_, _26170_);
  and (_10337_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_27026_, _10337_, _10336_);
  not (_10338_, _02406_);
  or (_10340_, _10338_, _25258_);
  or (_10342_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_10344_, _10342_, _23049_);
  and (_04947_, _10344_, _10340_);
  and (_10347_, _02484_, _26170_);
  and (_10348_, _02486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_27101_, _10348_, _10347_);
  and (_10351_, _26194_, _23768_);
  and (_10352_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_27102_, _10352_, _10351_);
  and (_10354_, _09484_, _23768_);
  and (_10355_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  or (_27138_, _10355_, _10354_);
  and (_10357_, _26194_, _26085_);
  and (_10358_, _26196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_27105_, _10358_, _10357_);
  and (_10360_, _09484_, _26170_);
  and (_10361_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or (_27139_, _10361_, _10360_);
  and (_10363_, _04812_, _25886_);
  and (_10365_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_27106_, _10365_, _10363_);
  and (_10366_, _09418_, _25886_);
  and (_10368_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_27110_, _10368_, _10366_);
  and (_10369_, _09484_, _25886_);
  and (_10370_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or (_27140_, _10370_, _10369_);
  and (_10371_, _09418_, _23768_);
  and (_10372_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_27108_, _10372_, _10371_);
  and (_10375_, _02825_, _25914_);
  and (_10377_, _10375_, _25886_);
  not (_10378_, _10375_);
  and (_10380_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or (_27025_, _10380_, _10377_);
  and (_10382_, _04181_, _23768_);
  and (_10383_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or (_27212_, _10383_, _10382_);
  and (_10384_, _10375_, _26170_);
  and (_10385_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or (_27024_, _10385_, _10384_);
  and (_10386_, _10375_, _25927_);
  and (_10387_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or (_27023_, _10387_, _10386_);
  and (_10388_, _05557_, _26242_);
  and (_10389_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_26974_, _10389_, _10388_);
  and (_10390_, _04027_, _26242_);
  and (_10391_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or (_05013_, _10391_, _10390_);
  and (_10392_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  and (_10393_, _10283_, _25886_);
  or (_27097_, _10393_, _10392_);
  and (_10394_, _05755_, _25886_);
  and (_10395_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_05043_, _10395_, _10394_);
  and (_10396_, _09182_, _26170_);
  and (_10397_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or (_05050_, _10397_, _10396_);
  and (_10398_, _05755_, _26170_);
  and (_10399_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_05054_, _10399_, _10398_);
  and (_10400_, _10375_, _26185_);
  and (_10401_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or (_05062_, _10401_, _10400_);
  and (_10402_, _10375_, _26085_);
  and (_10403_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or (_05074_, _10403_, _10402_);
  and (_10404_, _26213_, _23848_);
  and (_10405_, _10404_, _26170_);
  not (_10406_, _10404_);
  and (_10408_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_05101_, _10408_, _10405_);
  and (_10409_, _04181_, _26170_);
  and (_10410_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or (_05114_, _10410_, _10409_);
  and (_10411_, _04181_, _25927_);
  and (_10412_, _04184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or (_05123_, _10412_, _10411_);
  and (_10414_, _10404_, _25927_);
  and (_10415_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_27254_, _10415_, _10414_);
  and (_10416_, _00115_, _25927_);
  and (_10417_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_27067_, _10417_, _10416_);
  and (_10418_, _23227_, _23183_);
  and (_10419_, _26191_, _10418_);
  and (_10420_, _10419_, _26202_);
  and (_10422_, _10420_, _26085_);
  not (_10423_, _10420_);
  and (_10424_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or (_05172_, _10424_, _10422_);
  and (_10425_, _09791_, _26085_);
  and (_10426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_27015_, _10426_, _10425_);
  and (_10427_, _04027_, _26170_);
  and (_10428_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or (_05204_, _10428_, _10427_);
  and (_10429_, _09791_, _23830_);
  and (_10430_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_05207_, _10430_, _10429_);
  and (_10431_, _05755_, _25927_);
  and (_10432_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_05211_, _10432_, _10431_);
  and (_10433_, _04027_, _25927_);
  and (_10434_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or (_05213_, _10434_, _10433_);
  and (_10435_, _10420_, _26242_);
  and (_10436_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_05231_, _10436_, _10435_);
  and (_10437_, _04027_, _23768_);
  and (_10438_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or (_05233_, _10438_, _10437_);
  and (_10439_, _09756_, _23830_);
  and (_10440_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_05244_, _10440_, _10439_);
  and (_10441_, _09756_, _26185_);
  and (_10442_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_05250_, _10442_, _10441_);
  and (_10443_, _09182_, _25886_);
  and (_10445_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or (_27147_, _10445_, _10443_);
  and (_10446_, _10404_, _23768_);
  and (_10447_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_05262_, _10447_, _10446_);
  and (_10448_, _09786_, _23768_);
  and (_10450_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_05273_, _10450_, _10448_);
  and (_10451_, _09182_, _26085_);
  and (_10452_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  or (_27148_, _10452_, _10451_);
  and (_10453_, _09791_, _26242_);
  and (_10454_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_05291_, _10454_, _10453_);
  and (_10455_, _26202_, _26175_);
  and (_10456_, _10455_, _26185_);
  not (_10457_, _10455_);
  and (_10458_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_05298_, _10458_, _10456_);
  and (_10459_, _09182_, _26242_);
  and (_10460_, _09186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or (_05308_, _10460_, _10459_);
  and (_10461_, _04027_, _26085_);
  and (_10462_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or (_05311_, _10462_, _10461_);
  and (_10463_, _00095_, _25932_);
  and (_10464_, _10463_, _26185_);
  not (_10465_, _10463_);
  and (_10466_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_05335_, _10466_, _10464_);
  and (_10468_, _10463_, _26242_);
  and (_10469_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_05339_, _10469_, _10468_);
  and (_10471_, _10420_, _23768_);
  and (_10472_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or (_05343_, _10472_, _10471_);
  and (_10473_, _04027_, _23830_);
  and (_10474_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or (_05345_, _10474_, _10473_);
  and (_10475_, _26421_, _25938_);
  and (_10476_, _10475_, _26085_);
  not (_10477_, _10475_);
  and (_10478_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_05347_, _10478_, _10476_);
  and (_10479_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_10480_, _04120_, _26185_);
  or (_05349_, _10480_, _10479_);
  and (_10481_, _10475_, _23830_);
  and (_10482_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_05353_, _10482_, _10481_);
  and (_10483_, _10419_, _23220_);
  and (_10485_, _10483_, _26242_);
  not (_10486_, _10483_);
  and (_10487_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_27020_, _10487_, _10485_);
  and (_10488_, _10483_, _26185_);
  and (_10489_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_05364_, _10489_, _10488_);
  and (_10492_, _09791_, _23768_);
  and (_10493_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_05371_, _10493_, _10492_);
  and (_10494_, _09791_, _26170_);
  and (_10495_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_05378_, _10495_, _10494_);
  and (_10497_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  and (_10499_, _26541_, _26085_);
  or (_05381_, _10499_, _10497_);
  and (_10501_, _04027_, _25886_);
  and (_10502_, _04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or (_05386_, _10502_, _10501_);
  and (_10503_, _09791_, _25927_);
  and (_10504_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_05391_, _10504_, _10503_);
  and (_10506_, _04125_, _25886_);
  and (_10507_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or (_05413_, _10507_, _10506_);
  and (_10508_, _09053_, _23768_);
  and (_10509_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_05415_, _10509_, _10508_);
  and (_10510_, _10420_, _26170_);
  and (_10511_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_27022_, _10511_, _10510_);
  and (_10513_, _04163_, _23768_);
  and (_10514_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or (_05426_, _10514_, _10513_);
  and (_10515_, _10420_, _25927_);
  and (_10516_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_27021_, _10516_, _10515_);
  and (_10517_, _00115_, _26170_);
  and (_10518_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_05433_, _10518_, _10517_);
  and (_10521_, _04035_, _26170_);
  and (_10522_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_05436_, _10522_, _10521_);
  and (_10524_, _04175_, _25927_);
  and (_10525_, _04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_05440_, _10525_, _10524_);
  and (_10528_, _04163_, _25927_);
  and (_10529_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or (_05443_, _10529_, _10528_);
  and (_10530_, _04125_, _26185_);
  and (_10531_, _04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_05446_, _10531_, _10530_);
  and (_10532_, _09756_, _26242_);
  and (_10533_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_05448_, _10533_, _10532_);
  and (_10534_, _00115_, _23768_);
  and (_10535_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_05450_, _10535_, _10534_);
  and (_10538_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_10539_, _01608_, _23768_);
  or (_05454_, _10539_, _10538_);
  and (_10540_, _04035_, _25927_);
  and (_10541_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_05459_, _10541_, _10540_);
  and (_10542_, _04159_, _26085_);
  and (_10543_, _04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_05464_, _10543_, _10542_);
  and (_10544_, _00115_, _26185_);
  and (_10545_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_05468_, _10545_, _10544_);
  and (_10547_, _00115_, _25886_);
  and (_10548_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_05473_, _10548_, _10547_);
  and (_10549_, _08289_, _25886_);
  and (_10550_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or (_05480_, _10550_, _10549_);
  and (_10551_, _10483_, _23768_);
  and (_10552_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_05484_, _10552_, _10551_);
  and (_10553_, _00115_, _23830_);
  and (_10554_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_05486_, _10554_, _10553_);
  and (_10556_, _05557_, _26185_);
  and (_10558_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_05504_, _10558_, _10556_);
  and (_10559_, _04163_, _23830_);
  and (_10561_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  or (_05509_, _10561_, _10559_);
  and (_10562_, _00095_, _26202_);
  and (_10564_, _10562_, _26185_);
  not (_10565_, _10562_);
  and (_10566_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_05521_, _10566_, _10564_);
  and (_10567_, _04163_, _25886_);
  and (_10568_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  or (_05523_, _10568_, _10567_);
  and (_10569_, _10562_, _26085_);
  and (_10570_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_27043_, _10570_, _10569_);
  and (_10571_, _10483_, _25927_);
  and (_10573_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_05527_, _10573_, _10571_);
  and (_10575_, _04163_, _26085_);
  and (_10577_, _04165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or (_27141_, _10577_, _10575_);
  and (_10578_, _10562_, _23830_);
  and (_10579_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_05534_, _10579_, _10578_);
  and (_10581_, _04915_, _25927_);
  and (_10582_, _04917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_05537_, _10582_, _10581_);
  and (_10583_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_10584_, _26422_, _25927_);
  or (_05539_, _10584_, _10583_);
  and (_10585_, _08289_, _26185_);
  and (_10586_, _08291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_05544_, _10586_, _10585_);
  and (_10588_, _05826_, _25927_);
  and (_10589_, _05829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_05577_, _10589_, _10588_);
  and (_10591_, _04035_, _23830_);
  and (_10592_, _04038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_05579_, _10592_, _10591_);
  and (_10594_, _10562_, _26242_);
  and (_10595_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_05582_, _10595_, _10594_);
  and (_10596_, _10483_, _25886_);
  and (_10597_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_27019_, _10597_, _10596_);
  and (_10598_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_10599_, _10598_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_10600_, _10598_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_10602_, _10600_, _10599_);
  and (_05603_, _10602_, _23049_);
  and (_05606_, _24792_, _23049_);
  and (_05609_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _23049_);
  and (_10603_, _10483_, _23830_);
  and (_10605_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_05614_, _10605_, _10603_);
  and (_10607_, _04223_, _23830_);
  and (_10608_, _04226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or (_05617_, _10608_, _10607_);
  and (_10609_, _09484_, _26242_);
  and (_10610_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or (_05620_, _10610_, _10609_);
  and (_10612_, _09786_, _26242_);
  and (_10613_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_05622_, _10613_, _10612_);
  and (_10614_, _26733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_10615_, _26660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_10616_, _26660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_10617_, _10616_, _10615_);
  nor (_10618_, _10617_, _26732_);
  or (_10619_, _10618_, _26657_);
  or (_10621_, _10619_, _10614_);
  or (_10622_, _10617_, _26736_);
  and (_10623_, _10622_, _23049_);
  and (_05629_, _10623_, _10621_);
  and (_10624_, _09786_, _26185_);
  and (_10625_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_05631_, _10625_, _10624_);
  nand (_10627_, _26733_, _26659_);
  nand (_10629_, _10615_, _26657_);
  and (_10630_, _10629_, _23049_);
  and (_05635_, _10630_, _10627_);
  and (_10632_, _09484_, _26085_);
  and (_10633_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  or (_05638_, _10633_, _10632_);
  and (_10634_, _09786_, _26085_);
  and (_10635_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_27032_, _10635_, _10634_);
  and (_10637_, _26687_, _26675_);
  nand (_10638_, _26690_, _10637_);
  or (_10640_, _26703_, _26690_);
  and (_10641_, _10640_, _26660_);
  and (_10643_, _10641_, _10638_);
  or (_10644_, _10643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_10645_, _26712_, _26732_);
  or (_10646_, _26684_, _26665_);
  and (_10647_, _10646_, _10645_);
  or (_10649_, _10647_, _26692_);
  and (_10650_, _26692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_10651_, _10650_, _26736_);
  and (_10652_, _10651_, _23049_);
  and (_10653_, _10652_, _10649_);
  and (_05643_, _10653_, _10644_);
  and (_10655_, _09418_, _26185_);
  and (_10657_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_05645_, _10657_, _10655_);
  and (_10660_, _09228_, _26242_);
  and (_10661_, _09230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_05647_, _10661_, _10660_);
  and (_10662_, _09484_, _26185_);
  and (_10663_, _09486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or (_05649_, _10663_, _10662_);
  and (_10664_, _04041_, _26185_);
  and (_10666_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_05678_, _10666_, _10664_);
  and (_10667_, _10562_, _26170_);
  and (_10668_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_05681_, _10668_, _10667_);
  and (_10670_, _10419_, _26072_);
  and (_10672_, _10670_, _26170_);
  not (_10673_, _10670_);
  and (_10675_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_05685_, _10675_, _10672_);
  and (_10676_, _10562_, _25927_);
  and (_10677_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_05689_, _10677_, _10676_);
  and (_10680_, _10562_, _23768_);
  and (_10681_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_05707_, _10681_, _10680_);
  and (_10682_, _10670_, _25927_);
  and (_10683_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_05710_, _10683_, _10682_);
  and (_10685_, _04041_, _26085_);
  and (_10686_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_05713_, _10686_, _10685_);
  and (_10688_, _10670_, _23768_);
  and (_10689_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_05716_, _10689_, _10688_);
  and (_10690_, _04041_, _23830_);
  and (_10691_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_05725_, _10691_, _10690_);
  and (_10693_, _09786_, _23830_);
  and (_10695_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_05730_, _10695_, _10693_);
  and (_10697_, _09786_, _25886_);
  and (_10698_, _09788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_05737_, _10698_, _10697_);
  and (_10699_, _02849_, _26170_);
  and (_10700_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or (_05749_, _10700_, _10699_);
  and (_10702_, _10670_, _26185_);
  and (_10703_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_05754_, _10703_, _10702_);
  and (_10704_, _10029_, _26185_);
  and (_10705_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or (_05756_, _10705_, _10704_);
  and (_10706_, _10670_, _26085_);
  and (_10707_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_05760_, _10707_, _10706_);
  and (_10710_, _10029_, _26170_);
  and (_10711_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or (_27040_, _10711_, _10710_);
  and (_10714_, _10029_, _23768_);
  and (_10715_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or (_05763_, _10715_, _10714_);
  and (_10717_, _09998_, _26242_);
  and (_10719_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_05767_, _10719_, _10717_);
  and (_10721_, _01604_, _23768_);
  and (_10722_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_27235_, _10722_, _10721_);
  and (_10724_, _00095_, _26340_);
  and (_10725_, _10724_, _25927_);
  not (_10726_, _10724_);
  and (_10728_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_05769_, _10728_, _10725_);
  and (_10731_, _09998_, _23830_);
  and (_10732_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_05775_, _10732_, _10731_);
  and (_10734_, _10670_, _23830_);
  and (_10736_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_05778_, _10736_, _10734_);
  and (_10738_, _10724_, _23768_);
  and (_10739_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_05782_, _10739_, _10738_);
  and (_10740_, _09956_, _26085_);
  and (_10742_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_05789_, _10742_, _10740_);
  and (_10745_, _04041_, _26242_);
  and (_10746_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_05803_, _10746_, _10745_);
  and (_10748_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  and (_10750_, _10283_, _26085_);
  or (_05805_, _10750_, _10748_);
  and (_10751_, _09956_, _23768_);
  and (_10752_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_05807_, _10752_, _10751_);
  and (_10754_, _10404_, _25886_);
  and (_10756_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_05810_, _10756_, _10754_);
  and (_10759_, _09903_, _23830_);
  and (_10760_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or (_27035_, _10760_, _10759_);
  and (_10761_, _10404_, _26085_);
  and (_10762_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_27255_, _10762_, _10761_);
  and (_10763_, _09903_, _26170_);
  and (_10765_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or (_05817_, _10765_, _10763_);
  and (_10766_, _10724_, _26085_);
  and (_10767_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_05821_, _10767_, _10766_);
  and (_10768_, _10419_, _25932_);
  and (_10769_, _10768_, _25886_);
  not (_10770_, _10768_);
  and (_10772_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_05825_, _10772_, _10769_);
  and (_10775_, _10404_, _23830_);
  and (_10776_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_05828_, _10776_, _10775_);
  not (_10777_, _04851_);
  not (_10779_, _04870_);
  and (_10780_, _04887_, _04886_);
  and (_10782_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_10783_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_10784_, _10783_, _10782_);
  and (_10785_, _10784_, _04847_);
  not (_10786_, _04847_);
  and (_10788_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_10789_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_10790_, _10789_, _10788_);
  and (_10791_, _10790_, _10786_);
  or (_10793_, _10791_, _10785_);
  or (_10794_, _10793_, _10779_);
  not (_10795_, _04880_);
  and (_10797_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_10798_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_10800_, _10798_, _10797_);
  and (_10802_, _10800_, _04847_);
  and (_10804_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_10806_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_10807_, _10806_, _10804_);
  and (_10808_, _10807_, _10786_);
  or (_10810_, _10808_, _10802_);
  or (_10812_, _10810_, _04870_);
  and (_10814_, _10812_, _10795_);
  and (_10815_, _10814_, _10794_);
  or (_10816_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_10818_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_10820_, _10818_, _10816_);
  and (_10822_, _10820_, _04847_);
  or (_10823_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_10825_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_10826_, _10825_, _10823_);
  and (_10827_, _10826_, _10786_);
  or (_10828_, _10827_, _10822_);
  or (_10830_, _10828_, _10779_);
  or (_10832_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_10833_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_10834_, _10833_, _10832_);
  and (_10835_, _10834_, _04847_);
  or (_10836_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_10837_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_10838_, _10837_, _10836_);
  and (_10839_, _10838_, _10786_);
  or (_10840_, _10839_, _10835_);
  or (_10841_, _10840_, _04870_);
  and (_10842_, _10841_, _04880_);
  and (_10844_, _10842_, _10830_);
  or (_10846_, _10844_, _10815_);
  or (_10848_, _10846_, _10777_);
  not (_10849_, _04853_);
  and (_10850_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_10851_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_10852_, _10851_, _10850_);
  and (_10853_, _10852_, _04847_);
  and (_10855_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_10856_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_10857_, _10856_, _10855_);
  and (_10858_, _10857_, _10786_);
  or (_10859_, _10858_, _10853_);
  or (_10860_, _10859_, _10779_);
  and (_10861_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_10862_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_10863_, _10862_, _10861_);
  and (_10864_, _10863_, _04847_);
  and (_10865_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_10867_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_10868_, _10867_, _10865_);
  and (_10869_, _10868_, _10786_);
  or (_10870_, _10869_, _10864_);
  or (_10872_, _10870_, _04870_);
  and (_10873_, _10872_, _10795_);
  and (_10875_, _10873_, _10860_);
  or (_10876_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_10877_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_10878_, _10877_, _10786_);
  and (_10879_, _10878_, _10876_);
  or (_10881_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_10882_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_10883_, _10882_, _04847_);
  and (_10884_, _10883_, _10881_);
  or (_10885_, _10884_, _10879_);
  or (_10886_, _10885_, _10779_);
  or (_10887_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_10888_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_10890_, _10888_, _10786_);
  and (_10891_, _10890_, _10887_);
  or (_10893_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_10895_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_10896_, _10895_, _04847_);
  and (_10897_, _10896_, _10893_);
  or (_10898_, _10897_, _10891_);
  or (_10899_, _10898_, _04870_);
  and (_10901_, _10899_, _04880_);
  and (_10902_, _10901_, _10886_);
  or (_10904_, _10902_, _10875_);
  or (_10905_, _10904_, _04851_);
  and (_10906_, _10905_, _10849_);
  and (_10907_, _10906_, _10848_);
  and (_10909_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_10910_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_10911_, _10910_, _10909_);
  and (_10912_, _10911_, _04847_);
  and (_10913_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_10914_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_10916_, _10914_, _10913_);
  and (_10918_, _10916_, _10786_);
  or (_10921_, _10918_, _10912_);
  and (_10923_, _10921_, _04870_);
  and (_10924_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_10925_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_10926_, _10925_, _10924_);
  and (_10927_, _10926_, _04847_);
  and (_10929_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_10930_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_10932_, _10930_, _10929_);
  and (_10933_, _10932_, _10786_);
  or (_10935_, _10933_, _10927_);
  and (_10936_, _10935_, _10779_);
  or (_10937_, _10936_, _04880_);
  or (_10938_, _10937_, _10923_);
  or (_10939_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_10940_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_10942_, _10940_, _10786_);
  and (_10943_, _10942_, _10939_);
  or (_10944_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_10946_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_10947_, _10946_, _04847_);
  and (_10948_, _10947_, _10944_);
  or (_10949_, _10948_, _10943_);
  and (_10950_, _10949_, _04870_);
  or (_10951_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_10952_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_10953_, _10952_, _10786_);
  and (_10954_, _10953_, _10951_);
  or (_10956_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_10958_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_10959_, _10958_, _04847_);
  and (_10960_, _10959_, _10956_);
  or (_10961_, _10960_, _10954_);
  and (_10962_, _10961_, _10779_);
  or (_10963_, _10962_, _10795_);
  or (_10964_, _10963_, _10950_);
  and (_10965_, _10964_, _10938_);
  or (_10966_, _10965_, _04851_);
  and (_10967_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_10968_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_10969_, _10968_, _10967_);
  and (_10970_, _10969_, _04847_);
  and (_10971_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_10972_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_10974_, _10972_, _10971_);
  and (_10975_, _10974_, _10786_);
  or (_10977_, _10975_, _10970_);
  and (_10978_, _10977_, _04870_);
  and (_10980_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_10981_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_10983_, _10981_, _10980_);
  and (_10985_, _10983_, _04847_);
  and (_10986_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_10987_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_10988_, _10987_, _10986_);
  and (_10990_, _10988_, _10786_);
  or (_10991_, _10990_, _10985_);
  and (_10993_, _10991_, _10779_);
  or (_10994_, _10993_, _04880_);
  or (_10995_, _10994_, _10978_);
  or (_10996_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_10998_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_10999_, _10998_, _10996_);
  and (_11000_, _10999_, _04847_);
  or (_11001_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_11003_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_11005_, _11003_, _11001_);
  and (_11007_, _11005_, _10786_);
  or (_11008_, _11007_, _11000_);
  and (_11010_, _11008_, _04870_);
  or (_11012_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_11014_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_11016_, _11014_, _11012_);
  and (_11017_, _11016_, _04847_);
  or (_11018_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_11019_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_11020_, _11019_, _11018_);
  and (_11021_, _11020_, _10786_);
  or (_11022_, _11021_, _11017_);
  and (_11023_, _11022_, _10779_);
  or (_11025_, _11023_, _10795_);
  or (_11026_, _11025_, _11010_);
  and (_11028_, _11026_, _10995_);
  or (_11030_, _11028_, _10777_);
  and (_11031_, _11030_, _04853_);
  and (_11032_, _11031_, _10966_);
  or (_11034_, _11032_, _10907_);
  or (_11036_, _11034_, _04858_);
  not (_11038_, _04858_);
  and (_11040_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and (_11042_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_11043_, _11042_, _11040_);
  and (_11044_, _11043_, _04847_);
  and (_11045_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and (_11047_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_11049_, _11047_, _11045_);
  and (_11050_, _11049_, _10786_);
  or (_11051_, _11050_, _11044_);
  and (_11053_, _11051_, _04870_);
  and (_11054_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and (_11056_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_11058_, _11056_, _11054_);
  and (_11059_, _11058_, _04847_);
  and (_11060_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and (_11062_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_11064_, _11062_, _11060_);
  and (_11065_, _11064_, _10786_);
  or (_11067_, _11065_, _11059_);
  and (_11069_, _11067_, _10779_);
  or (_11070_, _11069_, _04880_);
  or (_11071_, _11070_, _11053_);
  or (_11072_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_11074_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and (_11075_, _11074_, _11072_);
  and (_11076_, _11075_, _04847_);
  or (_11077_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_11079_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  and (_11080_, _11079_, _11077_);
  and (_11082_, _11080_, _10786_);
  or (_11084_, _11082_, _11076_);
  and (_11085_, _11084_, _04870_);
  or (_11087_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_11088_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and (_11089_, _11088_, _11087_);
  and (_11091_, _11089_, _04847_);
  or (_11093_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_11095_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  and (_11097_, _11095_, _11093_);
  and (_11099_, _11097_, _10786_);
  or (_11101_, _11099_, _11091_);
  and (_11102_, _11101_, _10779_);
  or (_11103_, _11102_, _10795_);
  or (_11105_, _11103_, _11085_);
  and (_11106_, _11105_, _11071_);
  or (_11107_, _11106_, _04851_);
  and (_11109_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_11110_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_11111_, _11110_, _11109_);
  and (_11112_, _11111_, _04847_);
  and (_11113_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_11114_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_11116_, _11114_, _11113_);
  and (_11117_, _11116_, _10786_);
  or (_11118_, _11117_, _11112_);
  and (_11119_, _11118_, _04870_);
  and (_11120_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_11122_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_11123_, _11122_, _11120_);
  and (_11125_, _11123_, _04847_);
  and (_11127_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_11129_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_11130_, _11129_, _11127_);
  and (_11131_, _11130_, _10786_);
  or (_11132_, _11131_, _11125_);
  and (_11133_, _11132_, _10779_);
  or (_11135_, _11133_, _04880_);
  or (_11136_, _11135_, _11119_);
  or (_11138_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_11140_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_11142_, _11140_, _11138_);
  and (_11143_, _11142_, _04847_);
  or (_11144_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_11146_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_11147_, _11146_, _11144_);
  and (_11148_, _11147_, _10786_);
  or (_11149_, _11148_, _11143_);
  and (_11150_, _11149_, _04870_);
  or (_11151_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_11153_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_11154_, _11153_, _11151_);
  and (_11155_, _11154_, _04847_);
  or (_11156_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_11158_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_11160_, _11158_, _11156_);
  and (_11162_, _11160_, _10786_);
  or (_11164_, _11162_, _11155_);
  and (_11166_, _11164_, _10779_);
  or (_11168_, _11166_, _10795_);
  or (_11169_, _11168_, _11150_);
  and (_11170_, _11169_, _11136_);
  or (_11171_, _11170_, _10777_);
  and (_11172_, _11171_, _04853_);
  and (_11173_, _11172_, _11107_);
  and (_11175_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_11176_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_11177_, _11176_, _11175_);
  and (_11178_, _11177_, _10786_);
  and (_11179_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_11180_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_11181_, _11180_, _11179_);
  and (_11182_, _11181_, _04847_);
  or (_11184_, _11182_, _11178_);
  or (_11185_, _11184_, _10779_);
  and (_11187_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_11188_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_11189_, _11188_, _11187_);
  and (_11191_, _11189_, _10786_);
  and (_11192_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_11193_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_11194_, _11193_, _11192_);
  and (_11195_, _11194_, _04847_);
  or (_11196_, _11195_, _11191_);
  or (_11197_, _11196_, _04870_);
  and (_11199_, _11197_, _10795_);
  and (_11200_, _11199_, _11185_);
  or (_11201_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_11202_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_11204_, _11202_, _04847_);
  and (_11205_, _11204_, _11201_);
  or (_11206_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_11207_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_11208_, _11207_, _10786_);
  and (_11210_, _11208_, _11206_);
  or (_11212_, _11210_, _11205_);
  or (_11213_, _11212_, _10779_);
  or (_11214_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_11216_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_11217_, _11216_, _04847_);
  and (_11218_, _11217_, _11214_);
  or (_11219_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_11220_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_11221_, _11220_, _10786_);
  and (_11222_, _11221_, _11219_);
  or (_11224_, _11222_, _11218_);
  or (_11226_, _11224_, _04870_);
  and (_11227_, _11226_, _04880_);
  and (_11228_, _11227_, _11213_);
  or (_11230_, _11228_, _11200_);
  and (_11231_, _11230_, _10777_);
  and (_11233_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_11235_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_11237_, _11235_, _04847_);
  or (_11239_, _11237_, _11233_);
  and (_11241_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_11242_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_11243_, _11242_, _10786_);
  or (_11245_, _11243_, _11241_);
  and (_11247_, _11245_, _11239_);
  or (_11249_, _11247_, _10779_);
  and (_11250_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_11252_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_11253_, _11252_, _04847_);
  or (_11254_, _11253_, _11250_);
  and (_11255_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_11257_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_11259_, _11257_, _10786_);
  or (_11261_, _11259_, _11255_);
  and (_11262_, _11261_, _11254_);
  or (_11263_, _11262_, _04870_);
  and (_11264_, _11263_, _10795_);
  and (_11266_, _11264_, _11249_);
  or (_11267_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_11268_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_11270_, _11268_, _11267_);
  or (_11272_, _11270_, _10786_);
  or (_11273_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_11275_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_11277_, _11275_, _11273_);
  or (_11279_, _11277_, _04847_);
  and (_11281_, _11279_, _11272_);
  or (_11283_, _11281_, _10779_);
  or (_11285_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_11286_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_11287_, _11286_, _11285_);
  or (_11288_, _11287_, _10786_);
  or (_11290_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_11292_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_11294_, _11292_, _11290_);
  or (_11296_, _11294_, _04847_);
  and (_11298_, _11296_, _11288_);
  or (_11300_, _11298_, _04870_);
  and (_11302_, _11300_, _04880_);
  and (_11304_, _11302_, _11283_);
  or (_11305_, _11304_, _11266_);
  and (_11306_, _11305_, _04851_);
  or (_11307_, _11306_, _11231_);
  and (_11308_, _11307_, _10849_);
  or (_11310_, _11308_, _11173_);
  or (_11311_, _11310_, _11038_);
  and (_11312_, _11311_, _11036_);
  or (_11314_, _11312_, _25445_);
  and (_11315_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_11317_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_11319_, _11317_, _11315_);
  and (_11320_, _11319_, _04847_);
  and (_11321_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_11322_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_11324_, _11322_, _11321_);
  and (_11325_, _11324_, _10786_);
  or (_11327_, _11325_, _11320_);
  or (_11329_, _11327_, _10779_);
  and (_11331_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_11332_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_11333_, _11332_, _11331_);
  and (_11334_, _11333_, _04847_);
  and (_11335_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_11336_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_11338_, _11336_, _11335_);
  and (_11340_, _11338_, _10786_);
  or (_11341_, _11340_, _11334_);
  or (_11343_, _11341_, _04870_);
  and (_11345_, _11343_, _10795_);
  and (_11347_, _11345_, _11329_);
  or (_11348_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_11350_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_11352_, _11350_, _11348_);
  and (_11354_, _11352_, _04847_);
  or (_11355_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_11357_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_11358_, _11357_, _11355_);
  and (_11361_, _11358_, _10786_);
  or (_11363_, _11361_, _11354_);
  or (_11364_, _11363_, _10779_);
  or (_11366_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_11367_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_11368_, _11367_, _11366_);
  and (_11369_, _11368_, _04847_);
  or (_11370_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_11371_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_11372_, _11371_, _11370_);
  and (_11373_, _11372_, _10786_);
  or (_11374_, _11373_, _11369_);
  or (_11375_, _11374_, _04870_);
  and (_11376_, _11375_, _04880_);
  and (_11377_, _11376_, _11364_);
  or (_11378_, _11377_, _11347_);
  and (_11379_, _11378_, _04851_);
  and (_11380_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_11381_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_11382_, _11381_, _11380_);
  and (_11383_, _11382_, _04847_);
  and (_11384_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_11385_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_11386_, _11385_, _11384_);
  and (_11387_, _11386_, _10786_);
  or (_11388_, _11387_, _11383_);
  or (_11389_, _11388_, _10779_);
  and (_11390_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_11391_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_11392_, _11391_, _11390_);
  and (_11393_, _11392_, _04847_);
  and (_11394_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_11395_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_11396_, _11395_, _11394_);
  and (_11397_, _11396_, _10786_);
  or (_11399_, _11397_, _11393_);
  or (_11400_, _11399_, _04870_);
  and (_11401_, _11400_, _10795_);
  and (_11402_, _11401_, _11389_);
  or (_11404_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_11405_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_11406_, _11405_, _10786_);
  and (_11407_, _11406_, _11404_);
  or (_11408_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_11409_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_11410_, _11409_, _04847_);
  and (_11411_, _11410_, _11408_);
  or (_11412_, _11411_, _11407_);
  or (_11413_, _11412_, _10779_);
  or (_11414_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_11415_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_11416_, _11415_, _10786_);
  and (_11417_, _11416_, _11414_);
  or (_11419_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_11420_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_11421_, _11420_, _04847_);
  and (_11422_, _11421_, _11419_);
  or (_11424_, _11422_, _11417_);
  or (_11425_, _11424_, _04870_);
  and (_11426_, _11425_, _04880_);
  and (_11427_, _11426_, _11413_);
  or (_11428_, _11427_, _11402_);
  and (_11430_, _11428_, _10777_);
  or (_11431_, _11430_, _11379_);
  and (_11433_, _11431_, _10849_);
  and (_11434_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_11435_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_11436_, _11435_, _11434_);
  and (_11437_, _11436_, _04847_);
  and (_11438_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_11439_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_11440_, _11439_, _11438_);
  and (_11441_, _11440_, _10786_);
  or (_11442_, _11441_, _11437_);
  and (_11443_, _11442_, _04870_);
  and (_11444_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_11445_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_11447_, _11445_, _11444_);
  and (_11449_, _11447_, _04847_);
  and (_11450_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_11452_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_11453_, _11452_, _11450_);
  and (_11454_, _11453_, _10786_);
  or (_11456_, _11454_, _11449_);
  and (_11457_, _11456_, _10779_);
  or (_11458_, _11457_, _11443_);
  and (_11460_, _11458_, _10795_);
  or (_11461_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_11462_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_11463_, _11462_, _10786_);
  and (_11464_, _11463_, _11461_);
  or (_11465_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_11467_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_11468_, _11467_, _04847_);
  and (_11469_, _11468_, _11465_);
  or (_11470_, _11469_, _11464_);
  and (_11471_, _11470_, _04870_);
  or (_11472_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_11473_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_11474_, _11473_, _10786_);
  and (_11475_, _11474_, _11472_);
  or (_11476_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_11477_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_11478_, _11477_, _04847_);
  and (_11480_, _11478_, _11476_);
  or (_11482_, _11480_, _11475_);
  and (_11483_, _11482_, _10779_);
  or (_11484_, _11483_, _11471_);
  and (_11485_, _11484_, _04880_);
  or (_11486_, _11485_, _11460_);
  and (_11488_, _11486_, _10777_);
  and (_11489_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_11490_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_11492_, _11490_, _11489_);
  and (_11493_, _11492_, _04847_);
  and (_11494_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_11495_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_11496_, _11495_, _11494_);
  and (_11497_, _11496_, _10786_);
  or (_11498_, _11497_, _11493_);
  and (_11499_, _11498_, _04870_);
  and (_11500_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_11501_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_11502_, _11501_, _11500_);
  and (_11504_, _11502_, _04847_);
  and (_11505_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_11506_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_11507_, _11506_, _11505_);
  and (_11508_, _11507_, _10786_);
  or (_11509_, _11508_, _11504_);
  and (_11510_, _11509_, _10779_);
  or (_11511_, _11510_, _11499_);
  and (_11512_, _11511_, _10795_);
  or (_11513_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_11514_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_11515_, _11514_, _11513_);
  and (_11516_, _11515_, _04847_);
  or (_11517_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_11518_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_11519_, _11518_, _11517_);
  and (_11521_, _11519_, _10786_);
  or (_11522_, _11521_, _11516_);
  and (_11524_, _11522_, _04870_);
  or (_11525_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_11526_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_11527_, _11526_, _11525_);
  and (_11528_, _11527_, _04847_);
  or (_11529_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_11530_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_11531_, _11530_, _11529_);
  and (_11533_, _11531_, _10786_);
  or (_11535_, _11533_, _11528_);
  and (_11537_, _11535_, _10779_);
  or (_11538_, _11537_, _11524_);
  and (_11539_, _11538_, _04880_);
  or (_11540_, _11539_, _11512_);
  and (_11541_, _11540_, _04851_);
  or (_11542_, _11541_, _11488_);
  and (_11543_, _11542_, _04853_);
  or (_11544_, _11543_, _11433_);
  or (_11545_, _11544_, _04858_);
  and (_11546_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_11547_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_11548_, _11547_, _11546_);
  and (_11549_, _11548_, _04847_);
  and (_11551_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_11553_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_11555_, _11553_, _11551_);
  and (_11557_, _11555_, _10786_);
  or (_11559_, _11557_, _11549_);
  or (_11562_, _11559_, _10779_);
  and (_11564_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_11566_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_11568_, _11566_, _11564_);
  and (_11569_, _11568_, _04847_);
  and (_11570_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_11571_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_11573_, _11571_, _11570_);
  and (_11575_, _11573_, _10786_);
  or (_11577_, _11575_, _11569_);
  or (_11579_, _11577_, _04870_);
  and (_11580_, _11579_, _10795_);
  and (_11582_, _11580_, _11562_);
  or (_11583_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_11584_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_11586_, _11584_, _10786_);
  and (_11587_, _11586_, _11583_);
  or (_11588_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_11589_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_11590_, _11589_, _04847_);
  and (_11592_, _11590_, _11588_);
  or (_11593_, _11592_, _11587_);
  or (_11594_, _11593_, _10779_);
  or (_11595_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_11596_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_11597_, _11596_, _10786_);
  and (_11598_, _11597_, _11595_);
  or (_11599_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_11600_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_11601_, _11600_, _04847_);
  and (_11602_, _11601_, _11599_);
  or (_11603_, _11602_, _11598_);
  or (_11604_, _11603_, _04870_);
  and (_11605_, _11604_, _04880_);
  and (_11606_, _11605_, _11594_);
  or (_11607_, _11606_, _11582_);
  and (_11608_, _11607_, _10777_);
  and (_11609_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_11610_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_11611_, _11610_, _11609_);
  and (_11612_, _11611_, _04847_);
  and (_11613_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_11614_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_11615_, _11614_, _11613_);
  and (_11616_, _11615_, _10786_);
  or (_11617_, _11616_, _11612_);
  or (_11618_, _11617_, _10779_);
  and (_11619_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_11620_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_11621_, _11620_, _11619_);
  and (_11622_, _11621_, _04847_);
  and (_11623_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_11624_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_11625_, _11624_, _11623_);
  and (_11626_, _11625_, _10786_);
  or (_11627_, _11626_, _11622_);
  or (_11629_, _11627_, _04870_);
  and (_11630_, _11629_, _10795_);
  and (_11631_, _11630_, _11618_);
  or (_11632_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_11633_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_11634_, _11633_, _11632_);
  and (_11635_, _11634_, _04847_);
  or (_11636_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_11637_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_11638_, _11637_, _11636_);
  and (_11639_, _11638_, _10786_);
  or (_11640_, _11639_, _11635_);
  or (_11641_, _11640_, _10779_);
  or (_11642_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_11643_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_11644_, _11643_, _11642_);
  and (_11645_, _11644_, _04847_);
  or (_11646_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_11647_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_11648_, _11647_, _11646_);
  and (_11649_, _11648_, _10786_);
  or (_11650_, _11649_, _11645_);
  or (_11651_, _11650_, _04870_);
  and (_11652_, _11651_, _04880_);
  and (_11653_, _11652_, _11641_);
  or (_11654_, _11653_, _11631_);
  and (_11655_, _11654_, _04851_);
  or (_11656_, _11655_, _11608_);
  and (_11657_, _11656_, _10849_);
  or (_11658_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_11659_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_11660_, _11659_, _11658_);
  and (_11661_, _11660_, _04847_);
  or (_11662_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_11663_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_11664_, _11663_, _11662_);
  and (_11665_, _11664_, _10786_);
  or (_11666_, _11665_, _11661_);
  and (_11667_, _11666_, _10779_);
  or (_11668_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_11669_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _04847_);
  or (_11672_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_11673_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_11674_, _11673_, _11672_);
  and (_11675_, _11674_, _10786_);
  or (_11676_, _11675_, _11671_);
  and (_11677_, _11676_, _04870_);
  or (_11678_, _11677_, _11667_);
  and (_11679_, _11678_, _04880_);
  and (_11680_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_11681_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_11682_, _11681_, _11680_);
  and (_11684_, _11682_, _04847_);
  and (_11685_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_11686_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_11687_, _11686_, _11685_);
  and (_11688_, _11687_, _10786_);
  or (_11689_, _11688_, _11684_);
  and (_11690_, _11689_, _10779_);
  and (_11691_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_11692_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_11693_, _11692_, _11691_);
  and (_11694_, _11693_, _04847_);
  and (_11695_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_11696_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_11697_, _11696_, _11695_);
  and (_11698_, _11697_, _10786_);
  or (_11699_, _11698_, _11694_);
  and (_11700_, _11699_, _04870_);
  or (_11701_, _11700_, _11690_);
  and (_11702_, _11701_, _10795_);
  or (_11703_, _11702_, _11679_);
  and (_11704_, _11703_, _04851_);
  or (_11705_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_11706_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_11707_, _11706_, _10786_);
  and (_11708_, _11707_, _11705_);
  or (_11709_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_11710_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_11711_, _11710_, _04847_);
  and (_11712_, _11711_, _11709_);
  or (_11713_, _11712_, _11708_);
  and (_11714_, _11713_, _10779_);
  or (_11715_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_11716_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_11717_, _11716_, _10786_);
  and (_11718_, _11717_, _11715_);
  or (_11719_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_11720_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_11721_, _11720_, _04847_);
  and (_11722_, _11721_, _11719_);
  or (_11723_, _11722_, _11718_);
  and (_11724_, _11723_, _04870_);
  or (_11725_, _11724_, _11714_);
  and (_11726_, _11725_, _04880_);
  and (_11727_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_11728_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_11729_, _11728_, _11727_);
  and (_11730_, _11729_, _04847_);
  and (_11731_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_11732_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_11733_, _11732_, _11731_);
  and (_11734_, _11733_, _10786_);
  or (_11735_, _11734_, _11730_);
  and (_11736_, _11735_, _10779_);
  and (_11737_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_11738_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_11739_, _11738_, _11737_);
  and (_11740_, _11739_, _04847_);
  and (_11741_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_11742_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_11743_, _11742_, _11741_);
  and (_11744_, _11743_, _10786_);
  or (_11745_, _11744_, _11740_);
  and (_11746_, _11745_, _04870_);
  or (_11747_, _11746_, _11736_);
  and (_11748_, _11747_, _10795_);
  or (_11749_, _11748_, _11726_);
  and (_11750_, _11749_, _10777_);
  or (_11751_, _11750_, _11704_);
  and (_11752_, _11751_, _04853_);
  or (_11753_, _11752_, _11657_);
  or (_11755_, _11753_, _11038_);
  and (_11756_, _11755_, _11545_);
  or (_11757_, _11756_, _03372_);
  and (_11758_, _11757_, _11314_);
  or (_11759_, _11758_, _04902_);
  not (_11760_, _04902_);
  or (_11761_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_11762_, _11761_, _23049_);
  and (_05830_, _11762_, _11759_);
  and (_11763_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_11764_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_11765_, _11764_, _11763_);
  and (_11766_, _11765_, _04847_);
  and (_11767_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_11768_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_11769_, _11768_, _11767_);
  and (_11770_, _11769_, _10786_);
  or (_11771_, _11770_, _11766_);
  or (_11772_, _11771_, _10779_);
  and (_11773_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_11775_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_11776_, _11775_, _11773_);
  and (_11777_, _11776_, _04847_);
  and (_11778_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_11779_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_11780_, _11779_, _11778_);
  and (_11781_, _11780_, _10786_);
  or (_11782_, _11781_, _11777_);
  or (_11783_, _11782_, _04870_);
  and (_11784_, _11783_, _10795_);
  and (_11785_, _11784_, _11772_);
  or (_11786_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_11787_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_11788_, _11787_, _11786_);
  and (_11789_, _11788_, _04847_);
  or (_11790_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_11791_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_11792_, _11791_, _11790_);
  and (_11793_, _11792_, _10786_);
  or (_11794_, _11793_, _11789_);
  or (_11796_, _11794_, _10779_);
  or (_11797_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_11798_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_11799_, _11798_, _11797_);
  and (_11800_, _11799_, _04847_);
  or (_11801_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_11802_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_11803_, _11802_, _11801_);
  and (_11804_, _11803_, _10786_);
  or (_11805_, _11804_, _11800_);
  or (_11806_, _11805_, _04870_);
  and (_11807_, _11806_, _04880_);
  and (_11808_, _11807_, _11796_);
  or (_11809_, _11808_, _11785_);
  and (_11810_, _11809_, _04851_);
  and (_11811_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_11812_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_11813_, _11812_, _11811_);
  and (_11814_, _11813_, _04847_);
  and (_11815_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_11816_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_11817_, _11816_, _11815_);
  and (_11818_, _11817_, _10786_);
  or (_11819_, _11818_, _11814_);
  or (_11820_, _11819_, _10779_);
  and (_11821_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_11822_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_11823_, _11822_, _11821_);
  and (_11824_, _11823_, _04847_);
  and (_11825_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_11826_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_11827_, _11826_, _11825_);
  and (_11828_, _11827_, _10786_);
  or (_11829_, _11828_, _11824_);
  or (_11830_, _11829_, _04870_);
  and (_11831_, _11830_, _10795_);
  and (_11832_, _11831_, _11820_);
  or (_11833_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_11834_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_11835_, _11834_, _10786_);
  and (_11836_, _11835_, _11833_);
  or (_11837_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_11838_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_11839_, _11838_, _04847_);
  and (_11840_, _11839_, _11837_);
  or (_11841_, _11840_, _11836_);
  or (_11842_, _11841_, _10779_);
  or (_11843_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_11844_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_11845_, _11844_, _10786_);
  and (_11847_, _11845_, _11843_);
  or (_11848_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_11849_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_11850_, _11849_, _04847_);
  and (_11851_, _11850_, _11848_);
  or (_11852_, _11851_, _11847_);
  or (_11853_, _11852_, _04870_);
  and (_11854_, _11853_, _04880_);
  and (_11855_, _11854_, _11842_);
  or (_11856_, _11855_, _11832_);
  and (_11857_, _11856_, _10777_);
  or (_11858_, _11857_, _11810_);
  and (_11859_, _11858_, _10849_);
  and (_11860_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_11861_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_11862_, _11861_, _11860_);
  and (_11863_, _11862_, _04847_);
  and (_11864_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_11865_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_11866_, _11865_, _11864_);
  and (_11867_, _11866_, _10786_);
  or (_11868_, _11867_, _11863_);
  and (_11869_, _11868_, _04870_);
  and (_11870_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_11871_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_11872_, _11871_, _11870_);
  and (_11873_, _11872_, _04847_);
  and (_11874_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_11875_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_11876_, _11875_, _11874_);
  and (_11877_, _11876_, _10786_);
  or (_11878_, _11877_, _11873_);
  and (_11879_, _11878_, _10779_);
  or (_11880_, _11879_, _11869_);
  and (_11881_, _11880_, _10795_);
  or (_11882_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_11883_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_11884_, _11883_, _10786_);
  and (_11885_, _11884_, _11882_);
  or (_11886_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_11887_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_11888_, _11887_, _04847_);
  and (_11889_, _11888_, _11886_);
  or (_11890_, _11889_, _11885_);
  and (_11891_, _11890_, _04870_);
  or (_11892_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_11893_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_11894_, _11893_, _10786_);
  and (_11895_, _11894_, _11892_);
  or (_11896_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_11897_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_11898_, _11897_, _04847_);
  and (_11899_, _11898_, _11896_);
  or (_11900_, _11899_, _11895_);
  and (_11901_, _11900_, _10779_);
  or (_11902_, _11901_, _11891_);
  and (_11903_, _11902_, _04880_);
  or (_11904_, _11903_, _11881_);
  and (_11905_, _11904_, _10777_);
  and (_11906_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_11907_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_11908_, _11907_, _11906_);
  and (_11909_, _11908_, _04847_);
  and (_11910_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_11911_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_11912_, _11911_, _11910_);
  and (_11913_, _11912_, _10786_);
  or (_11914_, _11913_, _11909_);
  and (_11915_, _11914_, _04870_);
  and (_11916_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_11917_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_11918_, _11917_, _11916_);
  and (_11919_, _11918_, _04847_);
  and (_11920_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_11921_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_11922_, _11921_, _11920_);
  and (_11923_, _11922_, _10786_);
  or (_11924_, _11923_, _11919_);
  and (_11925_, _11924_, _10779_);
  or (_11926_, _11925_, _11915_);
  and (_11928_, _11926_, _10795_);
  or (_11929_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_11930_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_11931_, _11930_, _11929_);
  and (_11932_, _11931_, _04847_);
  or (_11933_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_11934_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_11935_, _11934_, _11933_);
  and (_11936_, _11935_, _10786_);
  or (_11937_, _11936_, _11932_);
  and (_11938_, _11937_, _04870_);
  or (_11939_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_11940_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_11941_, _11940_, _11939_);
  and (_11942_, _11941_, _04847_);
  or (_11943_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_11944_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_11945_, _11944_, _11943_);
  and (_11946_, _11945_, _10786_);
  or (_11947_, _11946_, _11942_);
  and (_11948_, _11947_, _10779_);
  or (_11949_, _11948_, _11938_);
  and (_11950_, _11949_, _04880_);
  or (_11951_, _11950_, _11928_);
  and (_11952_, _11951_, _04851_);
  or (_11953_, _11952_, _11905_);
  and (_11954_, _11953_, _04853_);
  or (_11955_, _11954_, _11859_);
  or (_11956_, _11955_, _04858_);
  and (_11957_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_11959_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_11960_, _11959_, _11957_);
  and (_11961_, _11960_, _04847_);
  and (_11962_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_11963_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_11964_, _11963_, _11962_);
  and (_11965_, _11964_, _10786_);
  or (_11966_, _11965_, _11961_);
  or (_11967_, _11966_, _10779_);
  and (_11968_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_11969_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_11970_, _11969_, _11968_);
  and (_11971_, _11970_, _04847_);
  and (_11972_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_11973_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_11974_, _11973_, _11972_);
  and (_11975_, _11974_, _10786_);
  or (_11976_, _11975_, _11971_);
  or (_11977_, _11976_, _04870_);
  and (_11978_, _11977_, _10795_);
  and (_11979_, _11978_, _11967_);
  or (_11980_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_11981_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_11982_, _11981_, _10786_);
  and (_11983_, _11982_, _11980_);
  or (_11984_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_11985_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_11986_, _11985_, _04847_);
  and (_11987_, _11986_, _11984_);
  or (_11988_, _11987_, _11983_);
  or (_11989_, _11988_, _10779_);
  or (_11990_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_11991_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_11992_, _11991_, _10786_);
  and (_11993_, _11992_, _11990_);
  or (_11994_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_11995_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_11996_, _11995_, _04847_);
  and (_11997_, _11996_, _11994_);
  or (_11998_, _11997_, _11993_);
  or (_12000_, _11998_, _04870_);
  and (_12001_, _12000_, _04880_);
  and (_12002_, _12001_, _11989_);
  or (_12003_, _12002_, _11979_);
  and (_12004_, _12003_, _10777_);
  and (_12005_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_12006_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_12007_, _12006_, _12005_);
  and (_12008_, _12007_, _04847_);
  and (_12009_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_12010_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_12011_, _12010_, _12009_);
  and (_12012_, _12011_, _10786_);
  or (_12013_, _12012_, _12008_);
  or (_12014_, _12013_, _10779_);
  and (_12015_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_12016_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_12017_, _12016_, _12015_);
  and (_12018_, _12017_, _04847_);
  and (_12019_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_12020_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_12021_, _12020_, _12019_);
  and (_12022_, _12021_, _10786_);
  or (_12023_, _12022_, _12018_);
  or (_12024_, _12023_, _04870_);
  and (_12025_, _12024_, _10795_);
  and (_12026_, _12025_, _12014_);
  or (_12027_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_12028_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_12029_, _12028_, _12027_);
  and (_12032_, _12029_, _04847_);
  or (_12033_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_12034_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_12035_, _12034_, _12033_);
  and (_12036_, _12035_, _10786_);
  or (_12037_, _12036_, _12032_);
  or (_12038_, _12037_, _10779_);
  or (_12039_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_12040_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_12041_, _12040_, _12039_);
  and (_12042_, _12041_, _04847_);
  or (_12043_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_12044_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_12045_, _12044_, _12043_);
  and (_12046_, _12045_, _10786_);
  or (_12047_, _12046_, _12042_);
  or (_12048_, _12047_, _04870_);
  and (_12049_, _12048_, _04880_);
  and (_12050_, _12049_, _12038_);
  or (_12051_, _12050_, _12026_);
  and (_12052_, _12051_, _04851_);
  or (_12053_, _12052_, _12004_);
  and (_12055_, _12053_, _10849_);
  or (_12056_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_12057_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_12058_, _12057_, _12056_);
  and (_12059_, _12058_, _04847_);
  or (_12060_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_12061_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_12062_, _12061_, _12060_);
  and (_12063_, _12062_, _10786_);
  or (_12064_, _12063_, _12059_);
  and (_12065_, _12064_, _10779_);
  or (_12066_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_12067_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_12068_, _12067_, _12066_);
  and (_12069_, _12068_, _04847_);
  or (_12070_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_12071_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_12073_, _12071_, _12070_);
  and (_12074_, _12073_, _10786_);
  or (_12075_, _12074_, _12069_);
  and (_12076_, _12075_, _04870_);
  or (_12077_, _12076_, _12065_);
  and (_12078_, _12077_, _04880_);
  and (_12079_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_12080_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_12081_, _12080_, _12079_);
  and (_12082_, _12081_, _04847_);
  and (_12083_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_12085_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_12086_, _12085_, _12083_);
  and (_12087_, _12086_, _10786_);
  or (_12088_, _12087_, _12082_);
  and (_12089_, _12088_, _10779_);
  and (_12090_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_12091_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_12092_, _12091_, _12090_);
  and (_12093_, _12092_, _04847_);
  and (_12094_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_12095_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_12096_, _12095_, _12094_);
  and (_12097_, _12096_, _10786_);
  or (_12099_, _12097_, _12093_);
  and (_12100_, _12099_, _04870_);
  or (_12101_, _12100_, _12089_);
  and (_12102_, _12101_, _10795_);
  or (_12103_, _12102_, _12078_);
  and (_12105_, _12103_, _04851_);
  or (_12106_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_12108_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_12109_, _12108_, _10786_);
  and (_12110_, _12109_, _12106_);
  or (_12111_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_12112_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_12113_, _12112_, _04847_);
  and (_12114_, _12113_, _12111_);
  or (_12115_, _12114_, _12110_);
  and (_12116_, _12115_, _10779_);
  or (_12117_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_12118_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and (_12119_, _12118_, _10786_);
  and (_12120_, _12119_, _12117_);
  or (_12121_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_12122_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and (_12123_, _12122_, _04847_);
  and (_12124_, _12123_, _12121_);
  or (_12125_, _12124_, _12120_);
  and (_12126_, _12125_, _04870_);
  or (_12127_, _12126_, _12116_);
  and (_12129_, _12127_, _04880_);
  and (_12130_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_12131_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_12132_, _12131_, _12130_);
  and (_12134_, _12132_, _04847_);
  and (_12136_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_12137_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_12138_, _12137_, _12136_);
  and (_12139_, _12138_, _10786_);
  or (_12140_, _12139_, _12134_);
  and (_12142_, _12140_, _10779_);
  and (_12143_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_12144_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_12145_, _12144_, _12143_);
  and (_12146_, _12145_, _04847_);
  and (_12147_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and (_12148_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_12149_, _12148_, _12147_);
  and (_12150_, _12149_, _10786_);
  or (_12152_, _12150_, _12146_);
  and (_12153_, _12152_, _04870_);
  or (_12154_, _12153_, _12142_);
  and (_12155_, _12154_, _10795_);
  or (_12156_, _12155_, _12129_);
  and (_12157_, _12156_, _10777_);
  or (_12158_, _12157_, _12105_);
  and (_12160_, _12158_, _04853_);
  or (_12161_, _12160_, _12055_);
  or (_12162_, _12161_, _11038_);
  and (_12163_, _12162_, _11956_);
  or (_12165_, _12163_, _25445_);
  and (_12167_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_12168_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_12169_, _12168_, _12167_);
  and (_12170_, _12169_, _04847_);
  and (_12171_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_12173_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_12175_, _12173_, _12171_);
  and (_12177_, _12175_, _10786_);
  or (_12178_, _12177_, _12170_);
  or (_12179_, _12178_, _10779_);
  and (_12180_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_12181_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_12182_, _12181_, _12180_);
  and (_12183_, _12182_, _04847_);
  and (_12184_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_12185_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_12186_, _12185_, _12184_);
  and (_12187_, _12186_, _10786_);
  or (_12188_, _12187_, _12183_);
  or (_12190_, _12188_, _04870_);
  and (_12191_, _12190_, _10795_);
  and (_12192_, _12191_, _12179_);
  or (_12193_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_12194_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_12195_, _12194_, _12193_);
  and (_12196_, _12195_, _04847_);
  or (_12198_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_12200_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_12201_, _12200_, _12198_);
  and (_12202_, _12201_, _10786_);
  or (_12203_, _12202_, _12196_);
  or (_12204_, _12203_, _10779_);
  or (_12206_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_12207_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_12209_, _12207_, _12206_);
  and (_12210_, _12209_, _04847_);
  or (_12211_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_12212_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_12213_, _12212_, _12211_);
  and (_12214_, _12213_, _10786_);
  or (_12216_, _12214_, _12210_);
  or (_12217_, _12216_, _04870_);
  and (_12218_, _12217_, _04880_);
  and (_12219_, _12218_, _12204_);
  or (_12220_, _12219_, _12192_);
  and (_12222_, _12220_, _04851_);
  and (_12223_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_12224_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_12225_, _12224_, _12223_);
  and (_12226_, _12225_, _04847_);
  and (_12227_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_12229_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_12231_, _12229_, _12227_);
  and (_12233_, _12231_, _10786_);
  or (_12234_, _12233_, _12226_);
  or (_12235_, _12234_, _10779_);
  and (_12236_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_12237_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_12238_, _12237_, _12236_);
  and (_12239_, _12238_, _04847_);
  and (_12240_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_12241_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_12243_, _12241_, _12240_);
  and (_12244_, _12243_, _10786_);
  or (_12245_, _12244_, _12239_);
  or (_12247_, _12245_, _04870_);
  and (_12249_, _12247_, _10795_);
  and (_12250_, _12249_, _12235_);
  or (_12251_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_12253_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_12254_, _12253_, _10786_);
  and (_12256_, _12254_, _12251_);
  or (_12257_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_12258_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_12259_, _12258_, _04847_);
  and (_12260_, _12259_, _12257_);
  or (_12262_, _12260_, _12256_);
  or (_12263_, _12262_, _10779_);
  or (_12264_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_12265_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_12266_, _12265_, _10786_);
  and (_12267_, _12266_, _12264_);
  or (_12268_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_12269_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_12270_, _12269_, _04847_);
  and (_12271_, _12270_, _12268_);
  or (_12272_, _12271_, _12267_);
  or (_12273_, _12272_, _04870_);
  and (_12274_, _12273_, _04880_);
  and (_12275_, _12274_, _12263_);
  or (_12276_, _12275_, _12250_);
  and (_12277_, _12276_, _10777_);
  or (_12278_, _12277_, _12222_);
  and (_12279_, _12278_, _10849_);
  and (_12280_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_12281_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_12282_, _12281_, _12280_);
  and (_12283_, _12282_, _04847_);
  and (_12284_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_12285_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_12286_, _12285_, _12284_);
  and (_12287_, _12286_, _10786_);
  or (_12288_, _12287_, _12283_);
  and (_12289_, _12288_, _04870_);
  and (_12290_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_12291_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_12292_, _12291_, _12290_);
  and (_12293_, _12292_, _04847_);
  and (_12294_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_12295_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_12296_, _12295_, _12294_);
  and (_12297_, _12296_, _10786_);
  or (_12298_, _12297_, _12293_);
  and (_12299_, _12298_, _10779_);
  or (_12300_, _12299_, _12289_);
  and (_12301_, _12300_, _10795_);
  or (_12302_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_12303_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_12304_, _12303_, _10786_);
  and (_12306_, _12304_, _12302_);
  or (_12307_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_12308_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_12309_, _12308_, _04847_);
  and (_12310_, _12309_, _12307_);
  or (_12311_, _12310_, _12306_);
  and (_12312_, _12311_, _04870_);
  or (_12313_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_12314_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_12315_, _12314_, _10786_);
  and (_12316_, _12315_, _12313_);
  or (_12317_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_12318_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_12319_, _12318_, _04847_);
  and (_12320_, _12319_, _12317_);
  or (_12321_, _12320_, _12316_);
  and (_12322_, _12321_, _10779_);
  or (_12323_, _12322_, _12312_);
  and (_12324_, _12323_, _04880_);
  or (_12325_, _12324_, _12301_);
  and (_12326_, _12325_, _10777_);
  and (_12327_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_12328_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_12329_, _12328_, _12327_);
  and (_12330_, _12329_, _04847_);
  and (_12331_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_12332_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_12333_, _12332_, _12331_);
  and (_12334_, _12333_, _10786_);
  or (_12335_, _12334_, _12330_);
  and (_12336_, _12335_, _04870_);
  and (_12337_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_12338_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_12339_, _12338_, _12337_);
  and (_12340_, _12339_, _04847_);
  and (_12341_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_12342_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_12343_, _12342_, _12341_);
  and (_12344_, _12343_, _10786_);
  or (_12345_, _12344_, _12340_);
  and (_12347_, _12345_, _10779_);
  or (_12348_, _12347_, _12336_);
  and (_12349_, _12348_, _10795_);
  or (_12350_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_12351_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_12352_, _12351_, _12350_);
  and (_12353_, _12352_, _04847_);
  or (_12354_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_12355_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_12356_, _12355_, _12354_);
  and (_12357_, _12356_, _10786_);
  or (_12358_, _12357_, _12353_);
  and (_12359_, _12358_, _04870_);
  or (_12360_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_12361_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_12362_, _12361_, _12360_);
  and (_12363_, _12362_, _04847_);
  or (_12364_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_12365_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_12366_, _12365_, _12364_);
  and (_12367_, _12366_, _10786_);
  or (_12368_, _12367_, _12363_);
  and (_12369_, _12368_, _10779_);
  or (_12370_, _12369_, _12359_);
  and (_12371_, _12370_, _04880_);
  or (_12372_, _12371_, _12349_);
  and (_12373_, _12372_, _04851_);
  or (_12374_, _12373_, _12326_);
  and (_12375_, _12374_, _04853_);
  or (_12376_, _12375_, _12279_);
  or (_12377_, _12376_, _04858_);
  and (_12378_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_12379_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_12380_, _12379_, _12378_);
  and (_12381_, _12380_, _04847_);
  and (_12382_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_12383_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_12384_, _12383_, _12382_);
  and (_12385_, _12384_, _10786_);
  or (_12386_, _12385_, _12381_);
  or (_12387_, _12386_, _10779_);
  and (_12388_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_12389_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_12390_, _12389_, _12388_);
  and (_12391_, _12390_, _04847_);
  and (_12392_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_12393_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_12394_, _12393_, _12392_);
  and (_12395_, _12394_, _10786_);
  or (_12396_, _12395_, _12391_);
  or (_12398_, _12396_, _04870_);
  and (_12399_, _12398_, _10795_);
  and (_12400_, _12399_, _12387_);
  or (_12401_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_12402_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_12403_, _12402_, _10786_);
  and (_12404_, _12403_, _12401_);
  or (_12405_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_12406_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_12407_, _12406_, _04847_);
  and (_12408_, _12407_, _12405_);
  or (_12409_, _12408_, _12404_);
  or (_12410_, _12409_, _10779_);
  or (_12411_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_12412_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_12413_, _12412_, _10786_);
  and (_12414_, _12413_, _12411_);
  or (_12415_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_12416_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_12417_, _12416_, _04847_);
  and (_12418_, _12417_, _12415_);
  or (_12419_, _12418_, _12414_);
  or (_12420_, _12419_, _04870_);
  and (_12421_, _12420_, _04880_);
  and (_12422_, _12421_, _12410_);
  or (_12423_, _12422_, _12400_);
  and (_12424_, _12423_, _10777_);
  and (_12425_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_12426_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_12427_, _12426_, _12425_);
  and (_12428_, _12427_, _04847_);
  and (_12429_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_12430_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_12431_, _12430_, _12429_);
  and (_12432_, _12431_, _10786_);
  or (_12433_, _12432_, _12428_);
  or (_12434_, _12433_, _10779_);
  and (_12435_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_12436_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_12437_, _12436_, _12435_);
  and (_12438_, _12437_, _04847_);
  and (_12439_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_12440_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_12441_, _12440_, _12439_);
  and (_12442_, _12441_, _10786_);
  or (_12443_, _12442_, _12438_);
  or (_12444_, _12443_, _04870_);
  and (_12445_, _12444_, _10795_);
  and (_12446_, _12445_, _12434_);
  or (_12447_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_12448_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_12449_, _12448_, _12447_);
  and (_12450_, _12449_, _04847_);
  or (_12451_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_12452_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_12453_, _12452_, _12451_);
  and (_12454_, _12453_, _10786_);
  or (_12455_, _12454_, _12450_);
  or (_12456_, _12455_, _10779_);
  or (_12457_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_12458_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_12459_, _12458_, _12457_);
  and (_12460_, _12459_, _04847_);
  or (_12461_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_12462_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_12463_, _12462_, _12461_);
  and (_12464_, _12463_, _10786_);
  or (_12465_, _12464_, _12460_);
  or (_12466_, _12465_, _04870_);
  and (_12467_, _12466_, _04880_);
  and (_12468_, _12467_, _12456_);
  or (_12469_, _12468_, _12446_);
  and (_12470_, _12469_, _04851_);
  or (_12471_, _12470_, _12424_);
  and (_12472_, _12471_, _10849_);
  or (_12473_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_12474_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_12475_, _12474_, _12473_);
  and (_12476_, _12475_, _04847_);
  or (_12477_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_12478_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_12479_, _12478_, _12477_);
  and (_12480_, _12479_, _10786_);
  or (_12481_, _12480_, _12476_);
  and (_12482_, _12481_, _10779_);
  or (_12483_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_12484_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_12485_, _12484_, _12483_);
  and (_12486_, _12485_, _04847_);
  or (_12487_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_12488_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_12489_, _12488_, _12487_);
  and (_12490_, _12489_, _10786_);
  or (_12491_, _12490_, _12486_);
  and (_12492_, _12491_, _04870_);
  or (_12493_, _12492_, _12482_);
  and (_12494_, _12493_, _04880_);
  and (_12495_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_12496_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_12497_, _12496_, _12495_);
  and (_12498_, _12497_, _04847_);
  and (_12499_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_12500_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_12501_, _12500_, _12499_);
  and (_12502_, _12501_, _10786_);
  or (_12503_, _12502_, _12498_);
  and (_12504_, _12503_, _10779_);
  and (_12505_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_12506_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_12507_, _12506_, _12505_);
  and (_12509_, _12507_, _04847_);
  and (_12510_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_12511_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_12512_, _12511_, _12510_);
  and (_12513_, _12512_, _10786_);
  or (_12514_, _12513_, _12509_);
  and (_12515_, _12514_, _04870_);
  or (_12516_, _12515_, _12504_);
  and (_12517_, _12516_, _10795_);
  or (_12518_, _12517_, _12494_);
  and (_12519_, _12518_, _04851_);
  or (_12520_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_12521_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_12522_, _12521_, _10786_);
  and (_12523_, _12522_, _12520_);
  or (_12524_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_12525_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_12526_, _12525_, _04847_);
  and (_12527_, _12526_, _12524_);
  or (_12528_, _12527_, _12523_);
  and (_12529_, _12528_, _10779_);
  or (_12530_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_12531_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_12532_, _12531_, _10786_);
  and (_12533_, _12532_, _12530_);
  or (_12534_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_12535_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_12536_, _12535_, _04847_);
  and (_12537_, _12536_, _12534_);
  or (_12538_, _12537_, _12533_);
  and (_12539_, _12538_, _04870_);
  or (_12540_, _12539_, _12529_);
  and (_12541_, _12540_, _04880_);
  and (_12542_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_12543_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_12544_, _12543_, _12542_);
  and (_12545_, _12544_, _04847_);
  and (_12546_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_12547_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_12548_, _12547_, _12546_);
  and (_12549_, _12548_, _10786_);
  or (_12550_, _12549_, _12545_);
  and (_12551_, _12550_, _10779_);
  and (_12552_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_12553_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_12554_, _12553_, _12552_);
  and (_12555_, _12554_, _04847_);
  and (_12556_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_12557_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_12558_, _12557_, _12556_);
  and (_12559_, _12558_, _10786_);
  or (_12560_, _12559_, _12555_);
  and (_12561_, _12560_, _04870_);
  or (_12562_, _12561_, _12551_);
  and (_12563_, _12562_, _10795_);
  or (_12564_, _12563_, _12541_);
  and (_12565_, _12564_, _10777_);
  or (_12566_, _12565_, _12519_);
  and (_12567_, _12566_, _04853_);
  or (_12568_, _12567_, _12472_);
  or (_12569_, _12568_, _11038_);
  and (_12570_, _12569_, _12377_);
  or (_12571_, _12570_, _03372_);
  and (_12572_, _12571_, _12165_);
  or (_12573_, _12572_, _04902_);
  or (_12574_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_12575_, _12574_, _23049_);
  and (_05832_, _12575_, _12573_);
  and (_12576_, _09886_, _26085_);
  and (_12577_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or (_05834_, _12577_, _12576_);
  and (_12578_, _10724_, _23830_);
  and (_12579_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_05836_, _12579_, _12578_);
  and (_12580_, _09886_, _26170_);
  and (_12581_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or (_27034_, _12581_, _12580_);
  and (_12582_, _10724_, _25886_);
  and (_12583_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_05845_, _12583_, _12582_);
  and (_12584_, _10768_, _26170_);
  and (_12585_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_05848_, _12585_, _12584_);
  and (_12586_, _09886_, _23768_);
  and (_12587_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or (_05851_, _12587_, _12586_);
  and (_12588_, _09852_, _26242_);
  and (_12589_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_05853_, _12589_, _12588_);
  and (_12590_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  and (_12591_, _10283_, _26185_);
  or (_05858_, _12591_, _12590_);
  and (_12592_, _09852_, _26085_);
  and (_12593_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_05865_, _12593_, _12592_);
  and (_12594_, _26548_, _25536_);
  nand (_12595_, _12594_, _23729_);
  or (_12596_, _12594_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_12597_, _12596_, _26547_);
  and (_12598_, _12597_, _12595_);
  nor (_12599_, _26547_, _25417_);
  or (_12600_, _12599_, _12598_);
  and (_05868_, _12600_, _23049_);
  nand (_12601_, _23167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_12602_, _12601_, _26523_);
  or (_12603_, _12602_, _00244_);
  and (_12604_, _12603_, _26621_);
  nand (_12605_, _26621_, _23167_);
  and (_12606_, _12605_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_12607_, _12606_, _26624_);
  or (_12609_, _12607_, _12604_);
  nand (_12610_, _26624_, _25332_);
  and (_12611_, _12610_, _23049_);
  and (_05873_, _12611_, _12609_);
  and (_12612_, _09852_, _25927_);
  and (_12613_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_05877_, _12613_, _12612_);
  and (_12614_, _09600_, _26185_);
  and (_12615_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or (_05881_, _12615_, _12614_);
  and (_12616_, _06946_, _26242_);
  and (_12617_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_05884_, _12617_, _12616_);
  and (_12618_, _04041_, _23768_);
  and (_12619_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_27207_, _12619_, _12618_);
  and (_12620_, _01564_, _23830_);
  and (_12621_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_05888_, _12621_, _12620_);
  and (_12622_, _09610_, _25927_);
  and (_12624_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_05890_, _12624_, _12622_);
  and (_12625_, _01564_, _25886_);
  and (_12626_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_05894_, _12626_, _12625_);
  and (_12627_, _09780_, _26185_);
  and (_12628_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_05914_, _12628_, _12627_);
  and (_12629_, _10768_, _26242_);
  and (_12630_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_05916_, _12630_, _12629_);
  and (_12631_, _09780_, _26170_);
  and (_12632_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_05921_, _12632_, _12631_);
  and (_12633_, _10768_, _26185_);
  and (_12634_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or (_27016_, _12634_, _12633_);
  and (_12635_, _10768_, _26085_);
  and (_12636_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or (_05924_, _12636_, _12635_);
  and (_12638_, _25916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_12639_, _26242_, _25915_);
  or (_27062_, _12639_, _12638_);
  and (_12640_, _01564_, _26242_);
  and (_12641_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_05931_, _12641_, _12640_);
  and (_12642_, _09732_, _26242_);
  and (_12643_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or (_05933_, _12643_, _12642_);
  and (_12644_, _09732_, _25886_);
  and (_12645_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or (_05941_, _12645_, _12644_);
  and (_12646_, _01564_, _26185_);
  and (_12647_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_05952_, _12647_, _12646_);
  and (_12648_, _09672_, _23830_);
  and (_12649_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or (_05956_, _12649_, _12648_);
  and (_12650_, _26283_, _26273_);
  and (_12651_, _12650_, _26185_);
  not (_12652_, _12650_);
  and (_12653_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or (_05959_, _12653_, _12651_);
  and (_12654_, _01564_, _26085_);
  and (_12655_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_05962_, _12655_, _12654_);
  and (_12656_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_12657_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_12658_, _12657_, _12656_);
  and (_12659_, _12658_, _04847_);
  and (_12660_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_12661_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_12662_, _12661_, _12660_);
  and (_12663_, _12662_, _10786_);
  or (_12664_, _12663_, _12659_);
  or (_12665_, _12664_, _10779_);
  and (_12666_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_12667_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_12668_, _12667_, _12666_);
  and (_12669_, _12668_, _04847_);
  and (_12670_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_12671_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_12672_, _12671_, _12670_);
  and (_12673_, _12672_, _10786_);
  or (_12674_, _12673_, _12669_);
  or (_12675_, _12674_, _04870_);
  and (_12676_, _12675_, _10795_);
  and (_12677_, _12676_, _12665_);
  or (_12678_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_12679_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_12680_, _12679_, _12678_);
  and (_12681_, _12680_, _04847_);
  or (_12682_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_12683_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_12684_, _12683_, _12682_);
  and (_12685_, _12684_, _10786_);
  or (_12686_, _12685_, _12681_);
  or (_12687_, _12686_, _10779_);
  or (_12688_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_12689_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_12690_, _12689_, _12688_);
  and (_12691_, _12690_, _04847_);
  or (_12692_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_12693_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_12694_, _12693_, _12692_);
  and (_12695_, _12694_, _10786_);
  or (_12696_, _12695_, _12691_);
  or (_12697_, _12696_, _04870_);
  and (_12698_, _12697_, _04880_);
  and (_12699_, _12698_, _12687_);
  or (_12700_, _12699_, _12677_);
  and (_12701_, _12700_, _04851_);
  and (_12702_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_12703_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_12704_, _12703_, _12702_);
  and (_12705_, _12704_, _04847_);
  and (_12706_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_12707_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_12708_, _12707_, _12706_);
  and (_12709_, _12708_, _10786_);
  or (_12710_, _12709_, _12705_);
  or (_12711_, _12710_, _10779_);
  and (_12712_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_12713_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_12714_, _12713_, _12712_);
  and (_12715_, _12714_, _04847_);
  and (_12716_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_12717_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_12718_, _12717_, _12716_);
  and (_12719_, _12718_, _10786_);
  or (_12720_, _12719_, _12715_);
  or (_12721_, _12720_, _04870_);
  and (_12722_, _12721_, _10795_);
  and (_12723_, _12722_, _12711_);
  or (_12724_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_12725_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_12726_, _12725_, _10786_);
  and (_12727_, _12726_, _12724_);
  or (_12728_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_12729_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_12730_, _12729_, _04847_);
  and (_12731_, _12730_, _12728_);
  or (_12732_, _12731_, _12727_);
  or (_12733_, _12732_, _10779_);
  or (_12734_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_12735_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_12736_, _12735_, _10786_);
  and (_12737_, _12736_, _12734_);
  or (_12738_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_12739_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_12740_, _12739_, _04847_);
  and (_12741_, _12740_, _12738_);
  or (_12742_, _12741_, _12737_);
  or (_12743_, _12742_, _04870_);
  and (_12744_, _12743_, _04880_);
  and (_12745_, _12744_, _12733_);
  or (_12746_, _12745_, _12723_);
  and (_12747_, _12746_, _10777_);
  or (_12748_, _12747_, _12701_);
  and (_12749_, _12748_, _10849_);
  and (_12751_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_12752_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_12753_, _12752_, _12751_);
  and (_12754_, _12753_, _04847_);
  and (_12755_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_12756_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_12757_, _12756_, _12755_);
  and (_12758_, _12757_, _10786_);
  or (_12759_, _12758_, _12754_);
  and (_12760_, _12759_, _04870_);
  and (_12761_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_12762_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_12763_, _12762_, _12761_);
  and (_12764_, _12763_, _04847_);
  and (_12765_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_12766_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_12767_, _12766_, _12765_);
  and (_12768_, _12767_, _10786_);
  or (_12769_, _12768_, _12764_);
  and (_12770_, _12769_, _10779_);
  or (_12771_, _12770_, _12760_);
  and (_12772_, _12771_, _10795_);
  or (_12773_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_12774_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_12775_, _12774_, _10786_);
  and (_12776_, _12775_, _12773_);
  or (_12777_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_12778_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_12779_, _12778_, _04847_);
  and (_12780_, _12779_, _12777_);
  or (_12781_, _12780_, _12776_);
  and (_12782_, _12781_, _04870_);
  or (_12783_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_12784_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_12785_, _12784_, _10786_);
  and (_12786_, _12785_, _12783_);
  or (_12787_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_12788_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_12789_, _12788_, _04847_);
  and (_12790_, _12789_, _12787_);
  or (_12792_, _12790_, _12786_);
  and (_12793_, _12792_, _10779_);
  or (_12794_, _12793_, _12782_);
  and (_12795_, _12794_, _04880_);
  or (_12796_, _12795_, _12772_);
  and (_12797_, _12796_, _10777_);
  and (_12798_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_12799_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_12800_, _12799_, _12798_);
  and (_12801_, _12800_, _04847_);
  and (_12802_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_12803_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_12804_, _12803_, _12802_);
  and (_12805_, _12804_, _10786_);
  or (_12806_, _12805_, _12801_);
  and (_12807_, _12806_, _04870_);
  and (_12808_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_12809_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_12810_, _12809_, _12808_);
  and (_12811_, _12810_, _04847_);
  and (_12813_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_12814_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_12815_, _12814_, _12813_);
  and (_12816_, _12815_, _10786_);
  or (_12817_, _12816_, _12811_);
  and (_12818_, _12817_, _10779_);
  or (_12819_, _12818_, _12807_);
  and (_12820_, _12819_, _10795_);
  or (_12821_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_12822_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_12823_, _12822_, _12821_);
  and (_12824_, _12823_, _04847_);
  or (_12825_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_12826_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_12827_, _12826_, _12825_);
  and (_12828_, _12827_, _10786_);
  or (_12829_, _12828_, _12824_);
  and (_12830_, _12829_, _04870_);
  or (_12831_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_12832_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_12833_, _12832_, _12831_);
  and (_12834_, _12833_, _04847_);
  or (_12835_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_12836_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, _10786_);
  or (_12839_, _12838_, _12834_);
  and (_12840_, _12839_, _10779_);
  or (_12841_, _12840_, _12830_);
  and (_12842_, _12841_, _04880_);
  or (_12843_, _12842_, _12820_);
  and (_12844_, _12843_, _04851_);
  or (_12845_, _12844_, _12797_);
  and (_12846_, _12845_, _04853_);
  or (_12847_, _12846_, _12749_);
  or (_12848_, _12847_, _04858_);
  and (_12849_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_12850_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_12851_, _12850_, _12849_);
  and (_12852_, _12851_, _04847_);
  and (_12853_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_12854_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_12855_, _12854_, _12853_);
  and (_12856_, _12855_, _10786_);
  or (_12857_, _12856_, _12852_);
  or (_12858_, _12857_, _10779_);
  and (_12859_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_12860_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_12861_, _12860_, _12859_);
  and (_12862_, _12861_, _04847_);
  and (_12863_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_12864_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_12865_, _12864_, _12863_);
  and (_12866_, _12865_, _10786_);
  or (_12867_, _12866_, _12862_);
  or (_12868_, _12867_, _04870_);
  and (_12869_, _12868_, _10795_);
  and (_12870_, _12869_, _12858_);
  or (_12871_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_12872_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_12873_, _12872_, _10786_);
  and (_12874_, _12873_, _12871_);
  or (_12875_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_12876_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_12877_, _12876_, _04847_);
  and (_12878_, _12877_, _12875_);
  or (_12879_, _12878_, _12874_);
  or (_12880_, _12879_, _10779_);
  or (_12881_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_12882_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_12883_, _12882_, _10786_);
  and (_12884_, _12883_, _12881_);
  or (_12885_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_12886_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_12887_, _12886_, _04847_);
  and (_12888_, _12887_, _12885_);
  or (_12889_, _12888_, _12884_);
  or (_12890_, _12889_, _04870_);
  and (_12891_, _12890_, _04880_);
  and (_12892_, _12891_, _12880_);
  or (_12893_, _12892_, _12870_);
  and (_12894_, _12893_, _10777_);
  and (_12895_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_12896_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_12897_, _12896_, _12895_);
  and (_12898_, _12897_, _04847_);
  and (_12899_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_12900_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _10786_);
  or (_12903_, _12902_, _12898_);
  or (_12904_, _12903_, _10779_);
  and (_12905_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_12906_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_12907_, _12906_, _12905_);
  and (_12908_, _12907_, _04847_);
  and (_12909_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_12910_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_12911_, _12910_, _12909_);
  and (_12912_, _12911_, _10786_);
  or (_12913_, _12912_, _12908_);
  or (_12914_, _12913_, _04870_);
  and (_12915_, _12914_, _10795_);
  and (_12916_, _12915_, _12904_);
  or (_12917_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_12918_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_12919_, _12918_, _12917_);
  and (_12920_, _12919_, _04847_);
  or (_12921_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_12922_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_12924_, _12922_, _12921_);
  and (_12925_, _12924_, _10786_);
  or (_12926_, _12925_, _12920_);
  or (_12927_, _12926_, _10779_);
  or (_12928_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_12929_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_12930_, _12929_, _12928_);
  and (_12931_, _12930_, _04847_);
  or (_12932_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_12933_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_12934_, _12933_, _12932_);
  and (_12935_, _12934_, _10786_);
  or (_12936_, _12935_, _12931_);
  or (_12937_, _12936_, _04870_);
  and (_12938_, _12937_, _04880_);
  and (_12939_, _12938_, _12927_);
  or (_12940_, _12939_, _12916_);
  and (_12941_, _12940_, _04851_);
  or (_12942_, _12941_, _12894_);
  and (_12943_, _12942_, _10849_);
  or (_12945_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_12946_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_12947_, _12946_, _12945_);
  and (_12948_, _12947_, _04847_);
  or (_12949_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_12950_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _10786_);
  or (_12953_, _12952_, _12948_);
  and (_12954_, _12953_, _10779_);
  or (_12955_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_12956_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_12957_, _12956_, _12955_);
  and (_12958_, _12957_, _04847_);
  or (_12959_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_12960_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_12961_, _12960_, _12959_);
  and (_12962_, _12961_, _10786_);
  or (_12963_, _12962_, _12958_);
  and (_12964_, _12963_, _04870_);
  or (_12965_, _12964_, _12954_);
  and (_12966_, _12965_, _04880_);
  and (_12967_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_12968_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_12969_, _12968_, _12967_);
  and (_12970_, _12969_, _04847_);
  and (_12971_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_12972_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_12973_, _12972_, _12971_);
  and (_12974_, _12973_, _10786_);
  or (_12975_, _12974_, _12970_);
  and (_12976_, _12975_, _10779_);
  and (_12977_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_12978_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_12979_, _12978_, _12977_);
  and (_12980_, _12979_, _04847_);
  and (_12981_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_12982_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_12983_, _12982_, _12981_);
  and (_12984_, _12983_, _10786_);
  or (_12985_, _12984_, _12980_);
  and (_12986_, _12985_, _04870_);
  or (_12987_, _12986_, _12976_);
  and (_12988_, _12987_, _10795_);
  or (_12989_, _12988_, _12966_);
  and (_12990_, _12989_, _04851_);
  or (_12991_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_12992_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_12993_, _12992_, _10786_);
  and (_12994_, _12993_, _12991_);
  or (_12995_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_12996_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_12997_, _12996_, _04847_);
  and (_12998_, _12997_, _12995_);
  or (_12999_, _12998_, _12994_);
  and (_13000_, _12999_, _10779_);
  or (_13001_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_13002_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_13003_, _13002_, _10786_);
  and (_13004_, _13003_, _13001_);
  or (_13005_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_13006_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_13007_, _13006_, _04847_);
  and (_13008_, _13007_, _13005_);
  or (_13009_, _13008_, _13004_);
  and (_13010_, _13009_, _04870_);
  or (_13011_, _13010_, _13000_);
  and (_13012_, _13011_, _04880_);
  and (_13013_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_13014_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_13015_, _13014_, _13013_);
  and (_13016_, _13015_, _04847_);
  and (_13017_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_13018_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_13019_, _13018_, _13017_);
  and (_13020_, _13019_, _10786_);
  or (_13021_, _13020_, _13016_);
  and (_13022_, _13021_, _10779_);
  and (_13023_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_13024_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_13025_, _13024_, _13023_);
  and (_13026_, _13025_, _04847_);
  and (_13027_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_13028_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_13029_, _13028_, _13027_);
  and (_13030_, _13029_, _10786_);
  or (_13031_, _13030_, _13026_);
  and (_13032_, _13031_, _04870_);
  or (_13033_, _13032_, _13022_);
  and (_13034_, _13033_, _10795_);
  or (_13035_, _13034_, _13012_);
  and (_13036_, _13035_, _10777_);
  or (_13037_, _13036_, _12990_);
  and (_13038_, _13037_, _04853_);
  or (_13039_, _13038_, _12943_);
  or (_13040_, _13039_, _11038_);
  and (_13041_, _13040_, _12848_);
  or (_13042_, _13041_, _25445_);
  and (_13043_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_13044_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_13045_, _13044_, _13043_);
  and (_13046_, _13045_, _04847_);
  and (_13047_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_13048_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_13049_, _13048_, _13047_);
  and (_13050_, _13049_, _10786_);
  or (_13051_, _13050_, _13046_);
  or (_13052_, _13051_, _10779_);
  and (_13053_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_13054_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_13055_, _13054_, _13053_);
  and (_13056_, _13055_, _04847_);
  and (_13057_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_13058_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_13059_, _13058_, _13057_);
  and (_13060_, _13059_, _10786_);
  or (_13061_, _13060_, _13056_);
  or (_13062_, _13061_, _04870_);
  and (_13063_, _13062_, _10795_);
  and (_13064_, _13063_, _13052_);
  or (_13065_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_13066_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_13067_, _13066_, _13065_);
  and (_13068_, _13067_, _04847_);
  or (_13069_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_13070_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_13071_, _13070_, _13069_);
  and (_13072_, _13071_, _10786_);
  or (_13073_, _13072_, _13068_);
  or (_13074_, _13073_, _10779_);
  or (_13075_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_13076_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_13077_, _13076_, _13075_);
  and (_13078_, _13077_, _04847_);
  or (_13079_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_13080_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_13081_, _13080_, _13079_);
  and (_13082_, _13081_, _10786_);
  or (_13083_, _13082_, _13078_);
  or (_13084_, _13083_, _04870_);
  and (_13085_, _13084_, _04880_);
  and (_13086_, _13085_, _13074_);
  or (_13087_, _13086_, _13064_);
  and (_13088_, _13087_, _04851_);
  and (_13089_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_13090_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_13091_, _13090_, _13089_);
  and (_13092_, _13091_, _04847_);
  and (_13093_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_13094_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_13096_, _13094_, _13093_);
  and (_13097_, _13096_, _10786_);
  or (_13098_, _13097_, _13092_);
  or (_13099_, _13098_, _10779_);
  and (_13100_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_13101_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_13102_, _13101_, _13100_);
  and (_13103_, _13102_, _04847_);
  and (_13104_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_13105_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _10786_);
  or (_13108_, _13107_, _13103_);
  or (_13109_, _13108_, _04870_);
  and (_13110_, _13109_, _10795_);
  and (_13111_, _13110_, _13099_);
  or (_13112_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_13113_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_13114_, _13113_, _10786_);
  and (_13115_, _13114_, _13112_);
  or (_13116_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_13117_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_13118_, _13117_, _04847_);
  and (_13119_, _13118_, _13116_);
  or (_13120_, _13119_, _13115_);
  or (_13121_, _13120_, _10779_);
  or (_13122_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_13123_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_13124_, _13123_, _10786_);
  and (_13125_, _13124_, _13122_);
  or (_13126_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_13127_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_13128_, _13127_, _04847_);
  and (_13129_, _13128_, _13126_);
  or (_13130_, _13129_, _13125_);
  or (_13131_, _13130_, _04870_);
  and (_13132_, _13131_, _04880_);
  and (_13133_, _13132_, _13121_);
  or (_13134_, _13133_, _13111_);
  and (_13135_, _13134_, _10777_);
  or (_13136_, _13135_, _13088_);
  and (_13137_, _13136_, _10849_);
  and (_13138_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_13139_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_13140_, _13139_, _13138_);
  and (_13141_, _13140_, _04847_);
  and (_13142_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_13143_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _10786_);
  or (_13146_, _13145_, _13141_);
  and (_13147_, _13146_, _04870_);
  and (_13148_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_13149_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_13150_, _13149_, _13148_);
  and (_13151_, _13150_, _04847_);
  and (_13152_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_13153_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_13154_, _13153_, _13152_);
  and (_13155_, _13154_, _10786_);
  or (_13156_, _13155_, _13151_);
  and (_13157_, _13156_, _10779_);
  or (_13158_, _13157_, _13147_);
  and (_13159_, _13158_, _10795_);
  or (_13160_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_13161_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_13162_, _13161_, _10786_);
  and (_13163_, _13162_, _13160_);
  or (_13164_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_13165_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_13166_, _13165_, _04847_);
  and (_13167_, _13166_, _13164_);
  or (_13168_, _13167_, _13163_);
  and (_13169_, _13168_, _04870_);
  or (_13170_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_13171_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_13172_, _13171_, _10786_);
  and (_13173_, _13172_, _13170_);
  or (_13174_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_13175_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_13176_, _13175_, _04847_);
  and (_13177_, _13176_, _13174_);
  or (_13178_, _13177_, _13173_);
  and (_13179_, _13178_, _10779_);
  or (_13180_, _13179_, _13169_);
  and (_13181_, _13180_, _04880_);
  or (_13182_, _13181_, _13159_);
  and (_13183_, _13182_, _10777_);
  and (_13184_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_13185_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_13186_, _13185_, _13184_);
  and (_13187_, _13186_, _04847_);
  and (_13188_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_13189_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_13190_, _13189_, _13188_);
  and (_13191_, _13190_, _10786_);
  or (_13192_, _13191_, _13187_);
  and (_13193_, _13192_, _04870_);
  and (_13194_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_13195_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_13196_, _13195_, _13194_);
  and (_13197_, _13196_, _04847_);
  and (_13198_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_13199_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_13200_, _13199_, _13198_);
  and (_13201_, _13200_, _10786_);
  or (_13202_, _13201_, _13197_);
  and (_13203_, _13202_, _10779_);
  or (_13204_, _13203_, _13193_);
  and (_13205_, _13204_, _10795_);
  or (_13206_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_13207_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_13208_, _13207_, _13206_);
  and (_13209_, _13208_, _04847_);
  or (_13210_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_13211_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_13212_, _13211_, _13210_);
  and (_13213_, _13212_, _10786_);
  or (_13214_, _13213_, _13209_);
  and (_13215_, _13214_, _04870_);
  or (_13217_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_13218_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_13219_, _13218_, _13217_);
  and (_13220_, _13219_, _04847_);
  or (_13221_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_13222_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_13223_, _13222_, _13221_);
  and (_13224_, _13223_, _10786_);
  or (_13225_, _13224_, _13220_);
  and (_13226_, _13225_, _10779_);
  or (_13227_, _13226_, _13215_);
  and (_13228_, _13227_, _04880_);
  or (_13229_, _13228_, _13205_);
  and (_13230_, _13229_, _04851_);
  or (_13231_, _13230_, _13183_);
  and (_13232_, _13231_, _04853_);
  or (_13233_, _13232_, _13137_);
  or (_13234_, _13233_, _04858_);
  and (_13235_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_13236_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_13237_, _13236_, _13235_);
  and (_13238_, _13237_, _04847_);
  and (_13239_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_13240_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_13241_, _13240_, _13239_);
  and (_13242_, _13241_, _10786_);
  or (_13243_, _13242_, _13238_);
  or (_13244_, _13243_, _10779_);
  and (_13245_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_13246_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_13247_, _13246_, _13245_);
  and (_13248_, _13247_, _04847_);
  and (_13249_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_13250_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_13251_, _13250_, _13249_);
  and (_13252_, _13251_, _10786_);
  or (_13253_, _13252_, _13248_);
  or (_13254_, _13253_, _04870_);
  and (_13255_, _13254_, _10795_);
  and (_13256_, _13255_, _13244_);
  or (_13257_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_13258_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_13259_, _13258_, _10786_);
  and (_13260_, _13259_, _13257_);
  or (_13261_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_13262_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_13263_, _13262_, _04847_);
  and (_13264_, _13263_, _13261_);
  or (_13265_, _13264_, _13260_);
  or (_13266_, _13265_, _10779_);
  or (_13267_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_13268_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_13269_, _13268_, _10786_);
  and (_13270_, _13269_, _13267_);
  or (_13271_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_13272_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_13273_, _13272_, _04847_);
  and (_13274_, _13273_, _13271_);
  or (_13275_, _13274_, _13270_);
  or (_13276_, _13275_, _04870_);
  and (_13277_, _13276_, _04880_);
  and (_13278_, _13277_, _13266_);
  or (_13279_, _13278_, _13256_);
  and (_13280_, _13279_, _10777_);
  and (_13281_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_13282_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_13283_, _13282_, _13281_);
  and (_13284_, _13283_, _04847_);
  and (_13285_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_13286_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_13287_, _13286_, _13285_);
  and (_13288_, _13287_, _10786_);
  or (_13289_, _13288_, _13284_);
  or (_13290_, _13289_, _10779_);
  and (_13291_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_13292_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_13293_, _13292_, _13291_);
  and (_13294_, _13293_, _04847_);
  and (_13295_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_13296_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_13297_, _13296_, _13295_);
  and (_13298_, _13297_, _10786_);
  or (_13299_, _13298_, _13294_);
  or (_13300_, _13299_, _04870_);
  and (_13301_, _13300_, _10795_);
  and (_13302_, _13301_, _13290_);
  or (_13303_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_13304_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_13305_, _13304_, _13303_);
  and (_13306_, _13305_, _04847_);
  or (_13307_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_13308_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_13309_, _13308_, _13307_);
  and (_13310_, _13309_, _10786_);
  or (_13311_, _13310_, _13306_);
  or (_13312_, _13311_, _10779_);
  or (_13313_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_13314_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_13315_, _13314_, _13313_);
  and (_13316_, _13315_, _04847_);
  or (_13317_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_13318_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_13319_, _13318_, _13317_);
  and (_13320_, _13319_, _10786_);
  or (_13321_, _13320_, _13316_);
  or (_13322_, _13321_, _04870_);
  and (_13323_, _13322_, _04880_);
  and (_13324_, _13323_, _13312_);
  or (_13325_, _13324_, _13302_);
  and (_13326_, _13325_, _04851_);
  or (_13328_, _13326_, _13280_);
  and (_13329_, _13328_, _10849_);
  or (_13330_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_13331_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_13332_, _13331_, _13330_);
  and (_13333_, _13332_, _04847_);
  or (_13334_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_13335_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_13336_, _13335_, _13334_);
  and (_13337_, _13336_, _10786_);
  or (_13338_, _13337_, _13333_);
  and (_13339_, _13338_, _10779_);
  or (_13340_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_13341_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_13342_, _13341_, _13340_);
  and (_13343_, _13342_, _04847_);
  or (_13344_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_13345_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_13346_, _13345_, _13344_);
  and (_13347_, _13346_, _10786_);
  or (_13349_, _13347_, _13343_);
  and (_13350_, _13349_, _04870_);
  or (_13351_, _13350_, _13339_);
  and (_13352_, _13351_, _04880_);
  and (_13353_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_13354_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _04847_);
  and (_13357_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_13358_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_13359_, _13358_, _13357_);
  and (_13360_, _13359_, _10786_);
  or (_13361_, _13360_, _13356_);
  and (_13362_, _13361_, _10779_);
  and (_13363_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_13364_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_13365_, _13364_, _13363_);
  and (_13366_, _13365_, _04847_);
  and (_13367_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_13368_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_13369_, _13368_, _13367_);
  and (_13370_, _13369_, _10786_);
  or (_13371_, _13370_, _13366_);
  and (_13372_, _13371_, _04870_);
  or (_13373_, _13372_, _13362_);
  and (_13374_, _13373_, _10795_);
  or (_13375_, _13374_, _13352_);
  and (_13376_, _13375_, _04851_);
  or (_13377_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_13378_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_13380_, _13378_, _10786_);
  and (_13381_, _13380_, _13377_);
  or (_13382_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_13383_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_13384_, _13383_, _04847_);
  and (_13385_, _13384_, _13382_);
  or (_13386_, _13385_, _13381_);
  and (_13387_, _13386_, _10779_);
  or (_13388_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_13389_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_13390_, _13389_, _10786_);
  and (_13391_, _13390_, _13388_);
  or (_13392_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_13393_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_13394_, _13393_, _04847_);
  and (_13395_, _13394_, _13392_);
  or (_13396_, _13395_, _13391_);
  and (_13397_, _13396_, _04870_);
  or (_13398_, _13397_, _13387_);
  and (_13399_, _13398_, _04880_);
  and (_13400_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_13401_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_13402_, _13401_, _13400_);
  and (_13403_, _13402_, _04847_);
  and (_13404_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_13405_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_13406_, _13405_, _13404_);
  and (_13407_, _13406_, _10786_);
  or (_13408_, _13407_, _13403_);
  and (_13409_, _13408_, _10779_);
  and (_13410_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_13411_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_13412_, _13411_, _13410_);
  and (_13413_, _13412_, _04847_);
  and (_13414_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_13415_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_13416_, _13415_, _13414_);
  and (_13417_, _13416_, _10786_);
  or (_13418_, _13417_, _13413_);
  and (_13419_, _13418_, _04870_);
  or (_13420_, _13419_, _13409_);
  and (_13421_, _13420_, _10795_);
  or (_13422_, _13421_, _13399_);
  and (_13423_, _13422_, _10777_);
  or (_13424_, _13423_, _13376_);
  and (_13425_, _13424_, _04853_);
  or (_13426_, _13425_, _13329_);
  or (_13427_, _13426_, _11038_);
  and (_13428_, _13427_, _13234_);
  or (_13429_, _13428_, _03372_);
  and (_13430_, _13429_, _13042_);
  or (_13431_, _13430_, _04902_);
  or (_13432_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_13433_, _13432_, _23049_);
  and (_05973_, _13433_, _13431_);
  and (_13434_, _09600_, _23768_);
  and (_13435_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or (_05979_, _13435_, _13434_);
  and (_13436_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_13437_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_13438_, _13437_, _13436_);
  and (_13439_, _13438_, _04847_);
  and (_13440_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_13441_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_13442_, _13441_, _13440_);
  and (_13443_, _13442_, _10786_);
  or (_13444_, _13443_, _13439_);
  or (_13445_, _13444_, _10779_);
  and (_13446_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_13447_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_13448_, _13447_, _13446_);
  and (_13449_, _13448_, _04847_);
  and (_13450_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_13451_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_13452_, _13451_, _13450_);
  and (_13453_, _13452_, _10786_);
  or (_13454_, _13453_, _13449_);
  or (_13455_, _13454_, _04870_);
  and (_13456_, _13455_, _10795_);
  and (_13457_, _13456_, _13445_);
  or (_13458_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_13459_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_13460_, _13459_, _13458_);
  and (_13461_, _13460_, _04847_);
  or (_13462_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_13463_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_13464_, _13463_, _13462_);
  and (_13465_, _13464_, _10786_);
  or (_13466_, _13465_, _13461_);
  or (_13467_, _13466_, _10779_);
  or (_13468_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_13469_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_13470_, _13469_, _13468_);
  and (_13471_, _13470_, _04847_);
  or (_13472_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_13473_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_13474_, _13473_, _13472_);
  and (_13475_, _13474_, _10786_);
  or (_13476_, _13475_, _13471_);
  or (_13477_, _13476_, _04870_);
  and (_13478_, _13477_, _04880_);
  and (_13479_, _13478_, _13467_);
  or (_13480_, _13479_, _13457_);
  and (_13481_, _13480_, _04851_);
  and (_13482_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_13483_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_13484_, _13483_, _13482_);
  and (_13485_, _13484_, _04847_);
  and (_13486_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_13487_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_13489_, _13487_, _13486_);
  and (_13490_, _13489_, _10786_);
  or (_13491_, _13490_, _13485_);
  or (_13492_, _13491_, _10779_);
  and (_13493_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_13494_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_13495_, _13494_, _13493_);
  and (_13496_, _13495_, _04847_);
  and (_13497_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_13498_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_13499_, _13498_, _13497_);
  and (_13500_, _13499_, _10786_);
  or (_13501_, _13500_, _13496_);
  or (_13502_, _13501_, _04870_);
  and (_13503_, _13502_, _10795_);
  and (_13504_, _13503_, _13492_);
  or (_13505_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_13506_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_13507_, _13506_, _10786_);
  and (_13508_, _13507_, _13505_);
  or (_13509_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_13510_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_13511_, _13510_, _04847_);
  and (_13512_, _13511_, _13509_);
  or (_13513_, _13512_, _13508_);
  or (_13514_, _13513_, _10779_);
  or (_13515_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_13516_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_13517_, _13516_, _10786_);
  and (_13518_, _13517_, _13515_);
  or (_13519_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_13520_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_13521_, _13520_, _04847_);
  and (_13522_, _13521_, _13519_);
  or (_13523_, _13522_, _13518_);
  or (_13524_, _13523_, _04870_);
  and (_13525_, _13524_, _04880_);
  and (_13526_, _13525_, _13514_);
  or (_13527_, _13526_, _13504_);
  and (_13528_, _13527_, _10777_);
  or (_13529_, _13528_, _13481_);
  and (_13530_, _13529_, _10849_);
  and (_13531_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_13532_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_13533_, _13532_, _13531_);
  and (_13534_, _13533_, _04847_);
  and (_13535_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_13536_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_13537_, _13536_, _13535_);
  and (_13538_, _13537_, _10786_);
  or (_13539_, _13538_, _13534_);
  and (_13540_, _13539_, _04870_);
  and (_13541_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_13542_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_13543_, _13542_, _13541_);
  and (_13544_, _13543_, _04847_);
  and (_13545_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_13546_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_13547_, _13546_, _13545_);
  and (_13548_, _13547_, _10786_);
  or (_13549_, _13548_, _13544_);
  and (_13550_, _13549_, _10779_);
  or (_13551_, _13550_, _13540_);
  and (_13552_, _13551_, _10795_);
  or (_13553_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_13554_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_13555_, _13554_, _10786_);
  and (_13556_, _13555_, _13553_);
  or (_13557_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_13558_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_13559_, _13558_, _04847_);
  and (_13560_, _13559_, _13557_);
  or (_13561_, _13560_, _13556_);
  and (_13562_, _13561_, _04870_);
  or (_13563_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_13564_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_13565_, _13564_, _10786_);
  and (_13566_, _13565_, _13563_);
  or (_13567_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_13568_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_13570_, _13568_, _04847_);
  and (_13571_, _13570_, _13567_);
  or (_13572_, _13571_, _13566_);
  and (_13573_, _13572_, _10779_);
  or (_13574_, _13573_, _13562_);
  and (_13575_, _13574_, _04880_);
  or (_13576_, _13575_, _13552_);
  and (_13577_, _13576_, _10777_);
  and (_13578_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_13579_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_13580_, _13579_, _13578_);
  and (_13581_, _13580_, _04847_);
  and (_13582_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_13583_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_13584_, _13583_, _13582_);
  and (_13585_, _13584_, _10786_);
  or (_13586_, _13585_, _13581_);
  and (_13587_, _13586_, _04870_);
  and (_13588_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_13589_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_13590_, _13589_, _13588_);
  and (_13591_, _13590_, _04847_);
  and (_13592_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_13593_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_13594_, _13593_, _13592_);
  and (_13595_, _13594_, _10786_);
  or (_13596_, _13595_, _13591_);
  and (_13597_, _13596_, _10779_);
  or (_13598_, _13597_, _13587_);
  and (_13599_, _13598_, _10795_);
  or (_13600_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_13601_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_13602_, _13601_, _13600_);
  and (_13603_, _13602_, _04847_);
  or (_13604_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_13605_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_13606_, _13605_, _13604_);
  and (_13607_, _13606_, _10786_);
  or (_13608_, _13607_, _13603_);
  and (_13609_, _13608_, _04870_);
  or (_13610_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_13611_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_13612_, _13611_, _13610_);
  and (_13613_, _13612_, _04847_);
  or (_13614_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_13615_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_13616_, _13615_, _13614_);
  and (_13617_, _13616_, _10786_);
  or (_13618_, _13617_, _13613_);
  and (_13619_, _13618_, _10779_);
  or (_13621_, _13619_, _13609_);
  and (_13622_, _13621_, _04880_);
  or (_13623_, _13622_, _13599_);
  and (_13624_, _13623_, _04851_);
  or (_13625_, _13624_, _13577_);
  and (_13626_, _13625_, _04853_);
  or (_13627_, _13626_, _13530_);
  or (_13628_, _13627_, _04858_);
  and (_13629_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_13630_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_13631_, _13630_, _13629_);
  and (_13632_, _13631_, _04847_);
  and (_13633_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_13634_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_13635_, _13634_, _13633_);
  and (_13636_, _13635_, _10786_);
  or (_13637_, _13636_, _13632_);
  or (_13638_, _13637_, _10779_);
  and (_13639_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_13640_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_13641_, _13640_, _13639_);
  and (_13642_, _13641_, _04847_);
  and (_13643_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_13644_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_13645_, _13644_, _13643_);
  and (_13646_, _13645_, _10786_);
  or (_13647_, _13646_, _13642_);
  or (_13648_, _13647_, _04870_);
  and (_13649_, _13648_, _10795_);
  and (_13650_, _13649_, _13638_);
  or (_13651_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_13652_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_13653_, _13652_, _10786_);
  and (_13654_, _13653_, _13651_);
  or (_13655_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_13656_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_13657_, _13656_, _04847_);
  and (_13658_, _13657_, _13655_);
  or (_13659_, _13658_, _13654_);
  or (_13660_, _13659_, _10779_);
  or (_13661_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_13662_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_13663_, _13662_, _10786_);
  and (_13664_, _13663_, _13661_);
  or (_13665_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_13666_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_13667_, _13666_, _04847_);
  and (_13668_, _13667_, _13665_);
  or (_13669_, _13668_, _13664_);
  or (_13670_, _13669_, _04870_);
  and (_13671_, _13670_, _04880_);
  and (_13672_, _13671_, _13660_);
  or (_13673_, _13672_, _13650_);
  and (_13674_, _13673_, _10777_);
  and (_13675_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_13676_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_13677_, _13676_, _13675_);
  and (_13678_, _13677_, _04847_);
  and (_13679_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_13680_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_13681_, _13680_, _13679_);
  and (_13682_, _13681_, _10786_);
  or (_13683_, _13682_, _13678_);
  or (_13684_, _13683_, _10779_);
  and (_13685_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_13686_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_13687_, _13686_, _13685_);
  and (_13688_, _13687_, _04847_);
  and (_13689_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_13690_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_13691_, _13690_, _13689_);
  and (_13692_, _13691_, _10786_);
  or (_13693_, _13692_, _13688_);
  or (_13694_, _13693_, _04870_);
  and (_13695_, _13694_, _10795_);
  and (_13696_, _13695_, _13684_);
  or (_13697_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_13698_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_13699_, _13698_, _13697_);
  and (_13700_, _13699_, _04847_);
  or (_13701_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_13702_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_13703_, _13702_, _13701_);
  and (_13704_, _13703_, _10786_);
  or (_13705_, _13704_, _13700_);
  or (_13706_, _13705_, _10779_);
  or (_13707_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_13708_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_13709_, _13708_, _13707_);
  and (_13710_, _13709_, _04847_);
  or (_13711_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_13712_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_13713_, _13712_, _13711_);
  and (_13714_, _13713_, _10786_);
  or (_13715_, _13714_, _13710_);
  or (_13716_, _13715_, _04870_);
  and (_13717_, _13716_, _04880_);
  and (_13718_, _13717_, _13706_);
  or (_13719_, _13718_, _13696_);
  and (_13720_, _13719_, _04851_);
  or (_13721_, _13720_, _13674_);
  and (_13722_, _13721_, _10849_);
  or (_13723_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_13724_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_13725_, _13724_, _13723_);
  and (_13726_, _13725_, _04847_);
  or (_13727_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_13728_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_13729_, _13728_, _13727_);
  and (_13730_, _13729_, _10786_);
  or (_13731_, _13730_, _13726_);
  and (_13732_, _13731_, _10779_);
  or (_13733_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_13734_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_13735_, _13734_, _13733_);
  and (_13736_, _13735_, _04847_);
  or (_13737_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_13738_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_13739_, _13738_, _13737_);
  and (_13740_, _13739_, _10786_);
  or (_13741_, _13740_, _13736_);
  and (_13742_, _13741_, _04870_);
  or (_13743_, _13742_, _13732_);
  and (_13744_, _13743_, _04880_);
  and (_13745_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_13746_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_13747_, _13746_, _13745_);
  and (_13748_, _13747_, _04847_);
  and (_13749_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_13750_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_13751_, _13750_, _13749_);
  and (_13752_, _13751_, _10786_);
  or (_13753_, _13752_, _13748_);
  and (_13754_, _13753_, _10779_);
  and (_13755_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_13756_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_13757_, _13756_, _13755_);
  and (_13758_, _13757_, _04847_);
  and (_13759_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_13760_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_13762_, _13760_, _13759_);
  and (_13763_, _13762_, _10786_);
  or (_13764_, _13763_, _13758_);
  and (_13765_, _13764_, _04870_);
  or (_13766_, _13765_, _13754_);
  and (_13767_, _13766_, _10795_);
  or (_13768_, _13767_, _13744_);
  and (_13769_, _13768_, _04851_);
  or (_13770_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_13771_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_13772_, _13771_, _10786_);
  and (_13773_, _13772_, _13770_);
  or (_13774_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_13775_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_13776_, _13775_, _04847_);
  and (_13777_, _13776_, _13774_);
  or (_13778_, _13777_, _13773_);
  and (_13779_, _13778_, _10779_);
  or (_13780_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_13781_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_13782_, _13781_, _10786_);
  and (_13783_, _13782_, _13780_);
  or (_13784_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_13785_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_13786_, _13785_, _04847_);
  and (_13787_, _13786_, _13784_);
  or (_13788_, _13787_, _13783_);
  and (_13789_, _13788_, _04870_);
  or (_13790_, _13789_, _13779_);
  and (_13791_, _13790_, _04880_);
  and (_13792_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_13793_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_13794_, _13793_, _13792_);
  and (_13795_, _13794_, _04847_);
  and (_13796_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_13797_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_13798_, _13797_, _13796_);
  and (_13799_, _13798_, _10786_);
  or (_13800_, _13799_, _13795_);
  and (_13801_, _13800_, _10779_);
  and (_13802_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_13803_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_13804_, _13803_, _13802_);
  and (_13805_, _13804_, _04847_);
  and (_13806_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_13807_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_13808_, _13807_, _13806_);
  and (_13809_, _13808_, _10786_);
  or (_13810_, _13809_, _13805_);
  and (_13811_, _13810_, _04870_);
  or (_13812_, _13811_, _13801_);
  and (_13813_, _13812_, _10795_);
  or (_13814_, _13813_, _13791_);
  and (_13815_, _13814_, _10777_);
  or (_13816_, _13815_, _13769_);
  and (_13817_, _13816_, _04853_);
  or (_13818_, _13817_, _13722_);
  or (_13819_, _13818_, _11038_);
  and (_13820_, _13819_, _13628_);
  or (_13821_, _13820_, _25445_);
  and (_13822_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_13823_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_13824_, _13823_, _13822_);
  and (_13825_, _13824_, _04847_);
  and (_13826_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_13827_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_13828_, _13827_, _13826_);
  and (_13829_, _13828_, _10786_);
  or (_13830_, _13829_, _13825_);
  or (_13831_, _13830_, _10779_);
  and (_13832_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_13833_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_13834_, _13833_, _13832_);
  and (_13835_, _13834_, _04847_);
  and (_13836_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_13837_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_13838_, _13837_, _13836_);
  and (_13839_, _13838_, _10786_);
  or (_13840_, _13839_, _13835_);
  or (_13841_, _13840_, _04870_);
  and (_13842_, _13841_, _10795_);
  and (_13843_, _13842_, _13831_);
  or (_13844_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_13845_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_13846_, _13845_, _13844_);
  and (_13847_, _13846_, _04847_);
  or (_13848_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_13849_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_13850_, _13849_, _13848_);
  and (_13851_, _13850_, _10786_);
  or (_13852_, _13851_, _13847_);
  or (_13853_, _13852_, _10779_);
  or (_13854_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_13855_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_13856_, _13855_, _13854_);
  and (_13857_, _13856_, _04847_);
  or (_13858_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_13859_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_13860_, _13859_, _13858_);
  and (_13861_, _13860_, _10786_);
  or (_13862_, _13861_, _13857_);
  or (_13863_, _13862_, _04870_);
  and (_13864_, _13863_, _04880_);
  and (_13865_, _13864_, _13853_);
  or (_13866_, _13865_, _13843_);
  and (_13867_, _13866_, _04851_);
  and (_13868_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_13869_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_13870_, _13869_, _13868_);
  and (_13871_, _13870_, _04847_);
  and (_13872_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_13873_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_13874_, _13873_, _13872_);
  and (_13875_, _13874_, _10786_);
  or (_13876_, _13875_, _13871_);
  or (_13877_, _13876_, _10779_);
  and (_13878_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_13879_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_13880_, _13879_, _13878_);
  and (_13881_, _13880_, _04847_);
  and (_13882_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_13883_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_13884_, _13883_, _13882_);
  and (_13885_, _13884_, _10786_);
  or (_13886_, _13885_, _13881_);
  or (_13887_, _13886_, _04870_);
  and (_13888_, _13887_, _10795_);
  and (_13889_, _13888_, _13877_);
  or (_13890_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_13891_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_13892_, _13891_, _10786_);
  and (_13893_, _13892_, _13890_);
  or (_13894_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_13895_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_13896_, _13895_, _04847_);
  and (_13897_, _13896_, _13894_);
  or (_13898_, _13897_, _13893_);
  or (_13899_, _13898_, _10779_);
  or (_13900_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_13901_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_13902_, _13901_, _10786_);
  and (_13903_, _13902_, _13900_);
  or (_13904_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_13905_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_13906_, _13905_, _04847_);
  and (_13907_, _13906_, _13904_);
  or (_13908_, _13907_, _13903_);
  or (_13909_, _13908_, _04870_);
  and (_13910_, _13909_, _04880_);
  and (_13911_, _13910_, _13899_);
  or (_13912_, _13911_, _13889_);
  and (_13913_, _13912_, _10777_);
  or (_13914_, _13913_, _13867_);
  and (_13915_, _13914_, _10849_);
  and (_13916_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_13917_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_13918_, _13917_, _13916_);
  and (_13919_, _13918_, _04847_);
  and (_13920_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_13921_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_13922_, _13921_, _13920_);
  and (_13923_, _13922_, _10786_);
  or (_13924_, _13923_, _13919_);
  and (_13925_, _13924_, _04870_);
  and (_13926_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_13927_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_13928_, _13927_, _13926_);
  and (_13929_, _13928_, _04847_);
  and (_13930_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_13931_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_13932_, _13931_, _13930_);
  and (_13933_, _13932_, _10786_);
  or (_13934_, _13933_, _13929_);
  and (_13935_, _13934_, _10779_);
  or (_13936_, _13935_, _13925_);
  and (_13937_, _13936_, _10795_);
  or (_13938_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_13939_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_13940_, _13939_, _10786_);
  and (_13941_, _13940_, _13938_);
  or (_13942_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_13943_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_13944_, _13943_, _04847_);
  and (_13945_, _13944_, _13942_);
  or (_13946_, _13945_, _13941_);
  and (_13947_, _13946_, _04870_);
  or (_13948_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_13949_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_13950_, _13949_, _10786_);
  and (_13951_, _13950_, _13948_);
  or (_13952_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_13953_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_13954_, _13953_, _04847_);
  and (_13955_, _13954_, _13952_);
  or (_13956_, _13955_, _13951_);
  and (_13957_, _13956_, _10779_);
  or (_13958_, _13957_, _13947_);
  and (_13959_, _13958_, _04880_);
  or (_13960_, _13959_, _13937_);
  and (_13961_, _13960_, _10777_);
  and (_13962_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_13963_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_13964_, _13963_, _13962_);
  and (_13965_, _13964_, _04847_);
  and (_13966_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_13967_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_13968_, _13967_, _13966_);
  and (_13969_, _13968_, _10786_);
  or (_13970_, _13969_, _13965_);
  and (_13971_, _13970_, _04870_);
  and (_13972_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_13973_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_13974_, _13973_, _13972_);
  and (_13975_, _13974_, _04847_);
  and (_13976_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_13977_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_13978_, _13977_, _13976_);
  and (_13979_, _13978_, _10786_);
  or (_13980_, _13979_, _13975_);
  and (_13981_, _13980_, _10779_);
  or (_13982_, _13981_, _13971_);
  and (_13983_, _13982_, _10795_);
  or (_13984_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_13985_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_13986_, _13985_, _13984_);
  and (_13987_, _13986_, _04847_);
  or (_13988_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_13989_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_13990_, _13989_, _13988_);
  and (_13991_, _13990_, _10786_);
  or (_13992_, _13991_, _13987_);
  and (_13993_, _13992_, _04870_);
  or (_13994_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_13995_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_13996_, _13995_, _13994_);
  and (_13997_, _13996_, _04847_);
  or (_13998_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_13999_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_14000_, _13999_, _13998_);
  and (_14001_, _14000_, _10786_);
  or (_14002_, _14001_, _13997_);
  and (_14003_, _14002_, _10779_);
  or (_14004_, _14003_, _13993_);
  and (_14005_, _14004_, _04880_);
  or (_14006_, _14005_, _13983_);
  and (_14007_, _14006_, _04851_);
  or (_14008_, _14007_, _13961_);
  and (_14009_, _14008_, _04853_);
  or (_14010_, _14009_, _13915_);
  or (_14011_, _14010_, _04858_);
  and (_14012_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_14013_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_14014_, _14013_, _14012_);
  and (_14015_, _14014_, _04847_);
  and (_14016_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_14017_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_14018_, _14017_, _14016_);
  and (_14019_, _14018_, _10786_);
  or (_14020_, _14019_, _14015_);
  or (_14021_, _14020_, _10779_);
  and (_14022_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_14023_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_14024_, _14023_, _14022_);
  and (_14025_, _14024_, _04847_);
  and (_14026_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_14027_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_14028_, _14027_, _14026_);
  and (_14029_, _14028_, _10786_);
  or (_14030_, _14029_, _14025_);
  or (_14031_, _14030_, _04870_);
  and (_14033_, _14031_, _10795_);
  and (_14034_, _14033_, _14021_);
  or (_14035_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_14036_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_14037_, _14036_, _10786_);
  and (_14038_, _14037_, _14035_);
  or (_14039_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_14040_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_14041_, _14040_, _04847_);
  and (_14042_, _14041_, _14039_);
  or (_14043_, _14042_, _14038_);
  or (_14044_, _14043_, _10779_);
  or (_14045_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_14046_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_14047_, _14046_, _10786_);
  and (_14048_, _14047_, _14045_);
  or (_14049_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_14050_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_14051_, _14050_, _04847_);
  and (_14052_, _14051_, _14049_);
  or (_14053_, _14052_, _14048_);
  or (_14054_, _14053_, _04870_);
  and (_14055_, _14054_, _04880_);
  and (_14056_, _14055_, _14044_);
  or (_14057_, _14056_, _14034_);
  and (_14058_, _14057_, _10777_);
  and (_14059_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_14060_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_14061_, _14060_, _14059_);
  and (_14062_, _14061_, _04847_);
  and (_14063_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_14064_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_14065_, _14064_, _14063_);
  and (_14066_, _14065_, _10786_);
  or (_14067_, _14066_, _14062_);
  or (_14068_, _14067_, _10779_);
  and (_14069_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_14070_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_14071_, _14070_, _14069_);
  and (_14072_, _14071_, _04847_);
  and (_14074_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_14075_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_14076_, _14075_, _14074_);
  and (_14077_, _14076_, _10786_);
  or (_14078_, _14077_, _14072_);
  or (_14079_, _14078_, _04870_);
  and (_14080_, _14079_, _10795_);
  and (_14081_, _14080_, _14068_);
  or (_14082_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_14083_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_14084_, _14083_, _14082_);
  and (_14085_, _14084_, _04847_);
  or (_14086_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_14087_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_14088_, _14087_, _14086_);
  and (_14089_, _14088_, _10786_);
  or (_14090_, _14089_, _14085_);
  or (_14091_, _14090_, _10779_);
  or (_14092_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_14093_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_14094_, _14093_, _14092_);
  and (_14095_, _14094_, _04847_);
  or (_14096_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_14097_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_14098_, _14097_, _14096_);
  and (_14099_, _14098_, _10786_);
  or (_14100_, _14099_, _14095_);
  or (_14101_, _14100_, _04870_);
  and (_14102_, _14101_, _04880_);
  and (_14103_, _14102_, _14091_);
  or (_14104_, _14103_, _14081_);
  and (_14105_, _14104_, _04851_);
  or (_14106_, _14105_, _14058_);
  and (_14107_, _14106_, _10849_);
  or (_14108_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_14109_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_14110_, _14109_, _14108_);
  and (_14111_, _14110_, _04847_);
  or (_14112_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_14113_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_14114_, _14113_, _14112_);
  and (_14115_, _14114_, _10786_);
  or (_14116_, _14115_, _14111_);
  and (_14117_, _14116_, _10779_);
  or (_14118_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_14119_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_14120_, _14119_, _14118_);
  and (_14121_, _14120_, _04847_);
  or (_14122_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_14123_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_14124_, _14123_, _14122_);
  and (_14125_, _14124_, _10786_);
  or (_14126_, _14125_, _14121_);
  and (_14127_, _14126_, _04870_);
  or (_14128_, _14127_, _14117_);
  and (_14129_, _14128_, _04880_);
  and (_14130_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_14131_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_14132_, _14131_, _14130_);
  and (_14133_, _14132_, _04847_);
  and (_14134_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_14135_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_14136_, _14135_, _14134_);
  and (_14137_, _14136_, _10786_);
  or (_14138_, _14137_, _14133_);
  and (_14139_, _14138_, _10779_);
  and (_14140_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_14141_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_14142_, _14141_, _14140_);
  and (_14143_, _14142_, _04847_);
  and (_14144_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_14145_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_14146_, _14145_, _14144_);
  and (_14147_, _14146_, _10786_);
  or (_14148_, _14147_, _14143_);
  and (_14149_, _14148_, _04870_);
  or (_14150_, _14149_, _14139_);
  and (_14151_, _14150_, _10795_);
  or (_14152_, _14151_, _14129_);
  and (_14153_, _14152_, _04851_);
  or (_14154_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_14155_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_14156_, _14155_, _10786_);
  and (_14157_, _14156_, _14154_);
  or (_14158_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_14159_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_14160_, _14159_, _04847_);
  and (_14161_, _14160_, _14158_);
  or (_14162_, _14161_, _14157_);
  and (_14163_, _14162_, _10779_);
  or (_14165_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_14166_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_14167_, _14166_, _10786_);
  and (_14168_, _14167_, _14165_);
  or (_14169_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_14170_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_14171_, _14170_, _04847_);
  and (_14172_, _14171_, _14169_);
  or (_14173_, _14172_, _14168_);
  and (_14174_, _14173_, _04870_);
  or (_14175_, _14174_, _14163_);
  and (_14176_, _14175_, _04880_);
  and (_14177_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_14178_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_14179_, _14178_, _14177_);
  and (_14180_, _14179_, _04847_);
  and (_14181_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_14182_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_14183_, _14182_, _14181_);
  and (_14184_, _14183_, _10786_);
  or (_14186_, _14184_, _14180_);
  and (_14187_, _14186_, _10779_);
  and (_14188_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_14189_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_14190_, _14189_, _14188_);
  and (_14191_, _14190_, _04847_);
  and (_14192_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_14193_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_14194_, _14193_, _14192_);
  and (_14195_, _14194_, _10786_);
  or (_14196_, _14195_, _14191_);
  and (_14197_, _14196_, _04870_);
  or (_14198_, _14197_, _14187_);
  and (_14199_, _14198_, _10795_);
  or (_14200_, _14199_, _14176_);
  and (_14201_, _14200_, _10777_);
  or (_14202_, _14201_, _14153_);
  and (_14203_, _14202_, _04853_);
  or (_14204_, _14203_, _14107_);
  or (_14205_, _14204_, _11038_);
  and (_14207_, _14205_, _14011_);
  or (_14208_, _14207_, _03372_);
  and (_14209_, _14208_, _13821_);
  or (_14210_, _14209_, _04902_);
  or (_14211_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_14212_, _14211_, _23049_);
  and (_27326_[5], _14212_, _14210_);
  and (_14213_, _09610_, _23830_);
  and (_14214_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_05986_, _14214_, _14213_);
  nand (_14215_, _26621_, _26473_);
  nor (_14216_, _14215_, _23729_);
  and (_14217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nor (_14218_, _26802_, _26742_);
  nor (_14219_, _14218_, _26659_);
  nand (_14220_, _14219_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_14221_, _01776_, _01743_);
  nor (_14222_, _14221_, _26659_);
  and (_14223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_14224_, _26660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_14225_, _14224_, _14223_);
  nand (_14226_, _14225_, _14222_);
  or (_14227_, _14226_, _14220_);
  and (_14228_, _14227_, _14217_);
  and (_14229_, _14228_, _14215_);
  or (_14230_, _14229_, _26624_);
  or (_14231_, _14230_, _14216_);
  nand (_14232_, _26624_, _25160_);
  and (_14233_, _14232_, _23049_);
  and (_05987_, _14233_, _14231_);
  and (_14234_, _10419_, _26340_);
  and (_14235_, _14234_, _25886_);
  not (_14236_, _14234_);
  and (_14237_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or (_05990_, _14237_, _14235_);
  and (_14238_, _26472_, _25536_);
  nand (_14239_, _14238_, _23729_);
  or (_14240_, _14238_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_14241_, _14240_, _26499_);
  and (_14242_, _14241_, _14239_);
  nor (_14244_, _26499_, _25417_);
  or (_14245_, _14244_, _14242_);
  and (_05997_, _14245_, _23049_);
  and (_14246_, _14234_, _23830_);
  and (_14247_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_05999_, _14247_, _14246_);
  and (_14248_, _10640_, _26723_);
  and (_14249_, _14248_, _10638_);
  or (_14250_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_14251_, _10647_, _26725_);
  and (_14252_, _14251_, _23049_);
  and (_06001_, _14252_, _14250_);
  and (_14253_, _04041_, _26170_);
  and (_14254_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_06008_, _14254_, _14253_);
  and (_14255_, _10029_, _23830_);
  and (_14256_, _10031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or (_06018_, _14256_, _14255_);
  and (_14257_, _10724_, _26242_);
  and (_14258_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_26988_, _14258_, _14257_);
  and (_14259_, _09998_, _25927_);
  and (_14260_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_27038_, _14260_, _14259_);
  and (_14261_, _04041_, _25927_);
  and (_14262_, _04044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_27208_, _14262_, _14261_);
  and (_14263_, _09956_, _26170_);
  and (_14264_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_06050_, _14264_, _14263_);
  and (_14265_, _09903_, _26185_);
  and (_14266_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or (_06053_, _14266_, _14265_);
  and (_14267_, _09886_, _26242_);
  and (_14268_, _09888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or (_06065_, _14268_, _14267_);
  not (_14269_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_14270_, _14219_, _14269_);
  nor (_14271_, _14225_, _26659_);
  nand (_14272_, _14271_, _14221_);
  or (_14274_, _14272_, _14270_);
  and (_14275_, _14274_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_14276_, _14275_, _04209_);
  and (_14277_, _26621_, _25536_);
  or (_14278_, _14277_, _14276_);
  nand (_14279_, _14277_, _23729_);
  and (_14280_, _14279_, _14278_);
  or (_14281_, _14280_, _26624_);
  nand (_14282_, _26624_, _25417_);
  and (_14283_, _14282_, _23049_);
  and (_06068_, _14283_, _14281_);
  and (_14284_, _10463_, _26170_);
  and (_14285_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_06075_, _14285_, _14284_);
  and (_14286_, _10463_, _25927_);
  and (_14287_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_06079_, _14287_, _14286_);
  and (_14288_, _26423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_14289_, _26422_, _23768_);
  or (_06082_, _14289_, _14288_);
  and (_14290_, _14234_, _26242_);
  and (_14291_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_06090_, _14291_, _14290_);
  and (_14292_, _01371_, _26185_);
  and (_14293_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_27234_, _14293_, _14292_);
  and (_14294_, _14234_, _26185_);
  and (_14295_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_06094_, _14295_, _14294_);
  nor (_14296_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _02500_);
  or (_14297_, _14270_, _14226_);
  and (_14298_, _14297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_14299_, _14298_, _14296_);
  and (_14300_, _26621_, _26136_);
  or (_14301_, _14300_, _14299_);
  nand (_14302_, _14300_, _23729_);
  and (_14303_, _14302_, _14301_);
  or (_14304_, _14303_, _26624_);
  nand (_14305_, _26624_, _25362_);
  and (_14306_, _14305_, _23049_);
  and (_06100_, _14306_, _14304_);
  and (_14307_, _09732_, _23768_);
  and (_14308_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or (_06105_, _14308_, _14307_);
  and (_14309_, _06946_, _26170_);
  and (_14310_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or (_06108_, _14310_, _14309_);
  and (_14311_, _09672_, _25927_);
  and (_14312_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or (_06116_, _14312_, _14311_);
  nand (_14313_, _26621_, _25224_);
  nor (_14314_, _14313_, _23729_);
  or (_14315_, _14271_, _14222_);
  or (_14316_, _14315_, _14220_);
  nand (_14317_, _14316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_14318_, _14317_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_14319_, _14318_, _14313_);
  or (_14320_, _14319_, _26624_);
  or (_14321_, _14320_, _14314_);
  nand (_14322_, _26624_, _25279_);
  and (_14323_, _14322_, _23049_);
  and (_06123_, _14323_, _14321_);
  and (_14324_, _09610_, _26185_);
  and (_14325_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_06126_, _14325_, _14324_);
  and (_14326_, _06946_, _25927_);
  and (_14327_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or (_06128_, _14327_, _14326_);
  and (_14328_, _09998_, _26085_);
  and (_14329_, _10000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_06145_, _14329_, _14328_);
  and (_14330_, _06946_, _23768_);
  and (_14331_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or (_27205_, _14331_, _14330_);
  and (_14332_, _10419_, _26421_);
  and (_14333_, _14332_, _23830_);
  not (_14334_, _14332_);
  and (_14335_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_27014_, _14335_, _14333_);
  and (_14336_, _09956_, _26185_);
  and (_14337_, _09960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_27037_, _14337_, _14336_);
  and (_14338_, _14332_, _26185_);
  and (_14339_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_06177_, _14339_, _14338_);
  and (_14340_, _09852_, _26170_);
  and (_14341_, _09855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_06183_, _14341_, _14340_);
  and (_14342_, _09610_, _26170_);
  and (_14343_, _09612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_06186_, _14343_, _14342_);
  and (_14344_, _14332_, _26085_);
  and (_14345_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_06188_, _14345_, _14344_);
  and (_14346_, _09780_, _25886_);
  and (_14347_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_06197_, _14347_, _14346_);
  and (_14348_, _09732_, _23830_);
  and (_14349_, _09734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or (_06205_, _14349_, _14348_);
  and (_14350_, _09672_, _26085_);
  and (_14351_, _09675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or (_06211_, _14351_, _14350_);
  and (_14352_, _10455_, _25927_);
  and (_14353_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_26972_, _14353_, _14352_);
  and (_14354_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_14355_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_14356_, _25943_, _14355_);
  or (_14357_, _14356_, _14354_);
  and (_26914_[15], _14357_, _23049_);
  and (_14358_, _09600_, _25927_);
  and (_14359_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or (_27033_, _14359_, _14358_);
  and (_14360_, _02849_, _25886_);
  and (_14361_, _02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or (_06220_, _14361_, _14360_);
  and (_14362_, _09903_, _26242_);
  and (_14363_, _09905_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or (_06227_, _14363_, _14362_);
  and (_14364_, _09600_, _25886_);
  and (_14365_, _09603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or (_06241_, _14365_, _14364_);
  and (_14366_, _10375_, _26242_);
  and (_14367_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or (_06278_, _14367_, _14366_);
  and (_06282_, _24685_, _23049_);
  and (_06284_, _24784_, _23049_);
  and (_06288_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _23049_);
  and (_06291_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _23049_);
  and (_06295_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _23049_);
  and (_14368_, _10670_, _26242_);
  and (_14369_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_27017_, _14369_, _14368_);
  and (_14370_, _10768_, _23768_);
  and (_14371_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or (_06310_, _14371_, _14370_);
  and (_14372_, _14332_, _25886_);
  and (_14373_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_06321_, _14373_, _14372_);
  or (_14374_, _23752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_14375_, _10598_, rst);
  and (_06331_, _14375_, _14374_);
  and (_14376_, _10419_, _26150_);
  and (_14377_, _14376_, _26085_);
  not (_14378_, _14376_);
  and (_14379_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_27013_, _14379_, _14377_);
  and (_06348_, _00479_, _23049_);
  nor (_06350_, _00583_, rst);
  and (_06351_, _00525_, _23049_);
  and (_06358_, _00635_, _23049_);
  and (_06375_, _00684_, _23049_);
  and (_06379_, _00800_, _23049_);
  and (_06381_, _00739_, _23049_);
  and (_14380_, _10419_, _23775_);
  and (_14381_, _14380_, _25886_);
  not (_14382_, _14380_);
  and (_14383_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_06391_, _14383_, _14381_);
  and (_14384_, _10419_, _26213_);
  and (_14385_, _14384_, _25886_);
  not (_14386_, _14384_);
  and (_14387_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_27002_, _14387_, _14385_);
  and (_14388_, _10419_, _26190_);
  and (_14389_, _14388_, _26085_);
  not (_14390_, _14388_);
  and (_14391_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or (_27000_, _14391_, _14389_);
  and (_14392_, _10419_, _25914_);
  and (_14393_, _14392_, _26085_);
  not (_14394_, _14392_);
  and (_14395_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_06406_, _14395_, _14393_);
  and (_14396_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  and (_14397_, _02019_, _23768_);
  or (_06409_, _14397_, _14396_);
  and (_14398_, _26273_, _26072_);
  and (_14399_, _14398_, _26185_);
  not (_14400_, _14398_);
  and (_14401_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_06421_, _14401_, _14399_);
  and (_14402_, _14398_, _25927_);
  and (_14403_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or (_06423_, _14403_, _14402_);
  and (_14404_, _26273_, _25932_);
  and (_14405_, _14404_, _25886_);
  not (_14406_, _14404_);
  and (_14407_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_06426_, _14407_, _14405_);
  and (_14408_, _26340_, _26273_);
  and (_14409_, _14408_, _26185_);
  not (_14410_, _14408_);
  and (_14411_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_06433_, _14411_, _14409_);
  and (_14412_, _26301_, _23830_);
  and (_14413_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_06440_, _14413_, _14412_);
  and (_14414_, _04825_, _26242_);
  and (_14415_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_26983_, _14415_, _14414_);
  and (_14416_, _05799_, _26185_);
  and (_14417_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_26979_, _14417_, _14416_);
  and (_14418_, _05799_, _26170_);
  and (_14419_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_06472_, _14419_, _14418_);
  and (_14420_, _26294_, _26185_);
  and (_14421_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_26975_, _14421_, _14420_);
  and (_14422_, _12650_, _26242_);
  and (_14423_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_06476_, _14423_, _14422_);
  and (_14424_, _05557_, _23830_);
  and (_14425_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_06482_, _14425_, _14424_);
  and (_14426_, _10455_, _23830_);
  and (_14427_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_06504_, _14427_, _14426_);
  and (_14428_, _09224_, _23768_);
  and (_14429_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_06511_, _14429_, _14428_);
  and (_14430_, _10420_, _23830_);
  and (_14431_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_06522_, _14431_, _14430_);
  and (_14432_, _14234_, _25927_);
  and (_14433_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_06523_, _14433_, _14432_);
  and (_14434_, _06946_, _26085_);
  and (_14435_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or (_06525_, _14435_, _14434_);
  and (_14436_, _14234_, _23768_);
  and (_14437_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or (_06530_, _14437_, _14436_);
  and (_14438_, _09176_, _25927_);
  and (_14439_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_06536_, _14439_, _14438_);
  and (_14440_, _10419_, _26224_);
  and (_14441_, _14440_, _26242_);
  not (_14442_, _14440_);
  and (_14443_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_27012_, _14443_, _14441_);
  and (_14444_, _06946_, _23830_);
  and (_14445_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or (_06540_, _14445_, _14444_);
  and (_14446_, _10419_, _26283_);
  and (_14447_, _14446_, _26170_);
  not (_14448_, _14446_);
  and (_14449_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_06543_, _14449_, _14447_);
  and (_14450_, _10419_, _26258_);
  and (_14451_, _14450_, _26242_);
  not (_14452_, _14450_);
  and (_14453_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_06547_, _14453_, _14451_);
  and (_14454_, _06946_, _25886_);
  and (_14455_, _06948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or (_06549_, _14455_, _14454_);
  and (_14456_, _10419_, _26374_);
  and (_14457_, _14456_, _26170_);
  not (_14458_, _14456_);
  and (_14459_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_06553_, _14459_, _14457_);
  and (_14460_, _14408_, _25927_);
  and (_14461_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_06561_, _14461_, _14460_);
  and (_14462_, _12650_, _25927_);
  and (_14463_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_06563_, _14463_, _14462_);
  and (_14464_, _26275_, _26185_);
  and (_14465_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_06568_, _14465_, _14464_);
  nand (_14466_, _01826_, _23215_);
  and (_14467_, _14466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_14468_, _25905_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_14469_, _14468_, _26475_);
  and (_14470_, _14469_, _01826_);
  or (_14471_, _14470_, _14467_);
  and (_14472_, _14471_, _25618_);
  nand (_14473_, _01834_, _25160_);
  or (_14474_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_14475_, _14474_, _25128_);
  and (_14476_, _14475_, _14473_);
  and (_14477_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_14478_, _14477_, rst);
  or (_14479_, _14478_, _14476_);
  or (_06571_, _14479_, _14472_);
  and (_14480_, _02102_, _26170_);
  and (_14481_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or (_06579_, _14481_, _14480_);
  nor (_14482_, _01574_, _00243_);
  nand (_14483_, _14482_, _23729_);
  or (_14484_, _14482_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_14485_, _14484_, _25618_);
  and (_14486_, _14485_, _14483_);
  nand (_14487_, _01578_, _25332_);
  or (_14488_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_14489_, _14488_, _25128_);
  and (_14490_, _14489_, _14487_);
  and (_14491_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_14492_, _14491_, rst);
  or (_14493_, _14492_, _14490_);
  or (_06582_, _14493_, _14486_);
  and (_14494_, _26294_, _23768_);
  and (_14495_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_06584_, _14495_, _14494_);
  and (_14496_, _10455_, _23768_);
  and (_14497_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_06594_, _14497_, _14496_);
  and (_14498_, _14376_, _26242_);
  and (_14499_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_06596_, _14499_, _14498_);
  and (_14500_, _14376_, _26185_);
  and (_14501_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_06598_, _14501_, _14500_);
  and (_14502_, _04047_, _26170_);
  and (_14503_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or (_06603_, _14503_, _14502_);
  nor (_14504_, _01574_, _01411_);
  nand (_14505_, _14504_, _23729_);
  or (_14506_, _14504_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_14507_, _14506_, _25618_);
  and (_14508_, _14507_, _14505_);
  nand (_14509_, _01578_, _25279_);
  or (_14510_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_14511_, _14510_, _25128_);
  and (_14512_, _14511_, _14509_);
  and (_14513_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_14514_, _14513_, rst);
  or (_14515_, _14514_, _14512_);
  or (_06629_, _14515_, _14508_);
  nor (_14516_, _00404_, _26556_);
  nand (_14517_, _14516_, _23729_);
  or (_14518_, _14516_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_14519_, _14518_, _25618_);
  and (_14520_, _14519_, _14517_);
  nand (_14521_, _00410_, _23824_);
  or (_14522_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_14523_, _14522_, _25128_);
  and (_14524_, _14523_, _14521_);
  and (_14525_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_14526_, _14525_, rst);
  or (_14527_, _14526_, _14524_);
  or (_06632_, _14527_, _14520_);
  and (_14528_, _10768_, _25927_);
  and (_14529_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_06635_, _14529_, _14528_);
  and (_14530_, _04047_, _25927_);
  and (_14531_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or (_27199_, _14531_, _14530_);
  and (_14532_, _04047_, _23768_);
  and (_14533_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or (_06639_, _14533_, _14532_);
  and (_14534_, _14384_, _23830_);
  and (_14535_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or (_06648_, _14535_, _14534_);
  and (_14536_, _14404_, _23830_);
  and (_14537_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_06654_, _14537_, _14536_);
  and (_14538_, _14332_, _26170_);
  and (_14539_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_06658_, _14539_, _14538_);
  and (_14540_, _04825_, _25886_);
  and (_14541_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or (_06660_, _14541_, _14540_);
  and (_14542_, _00249_, _25224_);
  or (_14543_, _14542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_14544_, _14543_, _25618_);
  nand (_14545_, _14542_, _23729_);
  and (_14546_, _14545_, _14544_);
  nand (_14547_, _00257_, _25279_);
  or (_14548_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_14549_, _14548_, _25128_);
  and (_14550_, _14549_, _14547_);
  and (_14551_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_14552_, _14551_, rst);
  or (_14553_, _14552_, _14550_);
  or (_06669_, _14553_, _14546_);
  and (_14554_, _14332_, _25927_);
  and (_14555_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_06671_, _14555_, _14554_);
  and (_14556_, _14332_, _23768_);
  and (_14557_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_06678_, _14557_, _14556_);
  and (_14558_, _26273_, _26150_);
  and (_14559_, _14558_, _26085_);
  not (_14560_, _14558_);
  and (_14561_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or (_06688_, _14561_, _14559_);
  and (_14562_, _04047_, _25886_);
  and (_14563_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or (_06696_, _14563_, _14562_);
  and (_14564_, _04047_, _26085_);
  and (_14565_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or (_27201_, _14565_, _14564_);
  and (_14566_, _04047_, _23830_);
  and (_14567_, _04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or (_27200_, _14567_, _14566_);
  and (_14568_, _14558_, _23830_);
  and (_14569_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or (_06701_, _14569_, _14568_);
  and (_14570_, _14558_, _26170_);
  and (_14571_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_06703_, _14571_, _14570_);
  and (_14572_, _14376_, _25927_);
  and (_14573_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_06723_, _14573_, _14572_);
  and (_14574_, _12650_, _26085_);
  and (_14575_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_06726_, _14575_, _14574_);
  and (_14577_, _12650_, _25886_);
  and (_14578_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or (_06728_, _14578_, _14577_);
  and (_14579_, _14376_, _23768_);
  and (_14580_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_06730_, _14580_, _14579_);
  and (_14581_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  and (_14582_, _00418_, _25927_);
  or (_06737_, _14582_, _14581_);
  and (_14583_, _09224_, _26242_);
  and (_14584_, _09226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_06742_, _14584_, _14583_);
  and (_14585_, _26176_, _23830_);
  and (_14586_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_06744_, _14586_, _14585_);
  and (_14587_, _09176_, _25886_);
  and (_14588_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_06752_, _14588_, _14587_);
  and (_14589_, _10455_, _26242_);
  and (_14590_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_06754_, _14590_, _14589_);
  and (_06756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _23049_);
  and (_14591_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _23049_);
  and (_06762_, _14591_, _26657_);
  and (_14592_, _05557_, _25927_);
  and (_14593_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_06765_, _14593_, _14592_);
  and (_14594_, _09053_, _25927_);
  and (_14595_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_06769_, _14595_, _14594_);
  and (_14596_, _26294_, _25886_);
  and (_14597_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_06776_, _14597_, _14596_);
  and (_14598_, _05799_, _26085_);
  and (_14599_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_06779_, _14599_, _14598_);
  and (_14600_, _05799_, _23768_);
  and (_14601_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_06788_, _14601_, _14600_);
  and (_14603_, _04194_, _25886_);
  and (_14604_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_06790_, _14604_, _14603_);
  and (_14605_, _14376_, _23830_);
  and (_14606_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_06795_, _14606_, _14605_);
  and (_14607_, _14376_, _25886_);
  and (_14608_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_06801_, _14608_, _14607_);
  and (_14609_, _04194_, _26170_);
  and (_14610_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_27198_, _14610_, _14609_);
  and (_14611_, _14376_, _26170_);
  and (_14612_, _14378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_06807_, _14612_, _14611_);
  and (_14613_, _02102_, _25927_);
  and (_14614_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_26980_, _14614_, _14613_);
  and (_14615_, _02102_, _26185_);
  and (_14616_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_06820_, _14616_, _14615_);
  and (_14617_, _04825_, _26170_);
  and (_14618_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_06825_, _14618_, _14617_);
  and (_14619_, _04825_, _23768_);
  and (_14620_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_06827_, _14620_, _14619_);
  and (_14621_, _04194_, _25927_);
  and (_14622_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_06846_, _14622_, _14621_);
  and (_14623_, _04825_, _26085_);
  and (_14624_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_06851_, _14624_, _14623_);
  and (_14625_, _26275_, _26085_);
  and (_14626_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_06856_, _14626_, _14625_);
  and (_14627_, _26275_, _26170_);
  and (_14628_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_06858_, _14628_, _14627_);
  and (_14629_, _26273_, _23847_);
  and (_14630_, _14629_, _25886_);
  not (_14631_, _14629_);
  and (_14632_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_26984_, _14632_, _14630_);
  and (_14633_, _12650_, _23768_);
  and (_14634_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or (_26986_, _14634_, _14633_);
  and (_14635_, _14440_, _25886_);
  and (_14636_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or (_06870_, _14636_, _14635_);
  and (_14637_, _14629_, _26185_);
  and (_14638_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_26985_, _14638_, _14637_);
  and (_14639_, _26421_, _26273_);
  and (_14640_, _14639_, _26170_);
  not (_14641_, _14639_);
  and (_14642_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or (_06876_, _14642_, _14640_);
  and (_14643_, _14440_, _26170_);
  and (_14644_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_06880_, _14644_, _14643_);
  and (_14645_, _14440_, _25927_);
  and (_14646_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_06883_, _14646_, _14645_);
  and (_14647_, _04194_, _26185_);
  and (_14648_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_06887_, _14648_, _14647_);
  and (_14649_, _04194_, _26085_);
  and (_14650_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_06891_, _14650_, _14649_);
  and (_14651_, _14404_, _23768_);
  and (_14652_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_06893_, _14652_, _14651_);
  and (_14653_, _14404_, _26185_);
  and (_14654_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_06897_, _14654_, _14653_);
  and (_14655_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_14656_, _04300_, _25927_);
  or (_06900_, _14656_, _14655_);
  and (_14657_, _26273_, _23220_);
  and (_14658_, _14657_, _23830_);
  not (_14659_, _14657_);
  and (_14660_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_26998_, _14660_, _14658_);
  and (_14661_, _04194_, _23830_);
  and (_14662_, _04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_06904_, _14662_, _14661_);
  and (_14663_, _12650_, _26170_);
  and (_14664_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or (_26987_, _14664_, _14663_);
  and (_14665_, _26273_, _26202_);
  and (_14666_, _14665_, _26170_);
  not (_14667_, _14665_);
  and (_14668_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_06910_, _14668_, _14666_);
  and (_14669_, _14440_, _26085_);
  and (_14670_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_06914_, _14670_, _14669_);
  and (_14671_, _14392_, _25927_);
  and (_14672_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_06935_, _14672_, _14671_);
  or (_14673_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_14674_, _14673_, _25891_);
  nand (_14675_, _03204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_14676_, _14675_, _25891_);
  or (_14677_, _14676_, _03206_);
  and (_14678_, _14677_, _14674_);
  or (_14679_, _14678_, _25903_);
  nand (_14680_, _25903_, _25417_);
  and (_14681_, _14680_, _23049_);
  and (_06939_, _14681_, _14679_);
  and (_14682_, _14440_, _23830_);
  and (_14683_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_06944_, _14683_, _14682_);
  and (_14684_, _14388_, _26242_);
  and (_14685_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_06945_, _14685_, _14684_);
  and (_14686_, _06836_, _26170_);
  and (_14687_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or (_06950_, _14687_, _14686_);
  and (_14688_, _14456_, _25927_);
  and (_14689_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_06952_, _14689_, _14688_);
  and (_14690_, _14450_, _25927_);
  and (_14691_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_27006_, _14691_, _14690_);
  and (_14692_, _14456_, _26185_);
  and (_14693_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_06960_, _14693_, _14692_);
  and (_14694_, _06836_, _25886_);
  and (_14695_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or (_27197_, _14695_, _14694_);
  and (_14696_, _14450_, _26185_);
  and (_14697_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_06963_, _14697_, _14696_);
  and (_14698_, _14446_, _26085_);
  and (_14699_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_06966_, _14699_, _14698_);
  and (_14700_, _14450_, _23830_);
  and (_14701_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_06969_, _14701_, _14700_);
  and (_14702_, _10419_, _23847_);
  and (_14703_, _14702_, _23830_);
  not (_14704_, _14702_);
  and (_14705_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or (_06972_, _14705_, _14703_);
  and (_14706_, _14446_, _23830_);
  and (_14707_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_06975_, _14707_, _14706_);
  and (_14708_, _14446_, _25927_);
  and (_14709_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_06977_, _14709_, _14708_);
  and (_14710_, _14440_, _23768_);
  and (_14711_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or (_27011_, _14711_, _14710_);
  and (_14712_, _14440_, _26185_);
  and (_14713_, _14442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_06981_, _14713_, _14712_);
  and (_14714_, _14446_, _25886_);
  and (_14715_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_27010_, _14715_, _14714_);
  and (_14717_, _09176_, _26085_);
  and (_14718_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_06992_, _14718_, _14717_);
  and (_14719_, _00016_, _25927_);
  and (_14720_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_06994_, _14720_, _14719_);
  and (_14721_, _14234_, _26170_);
  and (_14722_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_06996_, _14722_, _14721_);
  and (_14723_, _14332_, _26242_);
  and (_14724_, _14334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_06998_, _14724_, _14723_);
  and (_14725_, _14234_, _26085_);
  and (_14726_, _14236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or (_07000_, _14726_, _14725_);
  and (_14727_, _05557_, _23768_);
  and (_14728_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_07002_, _14728_, _14727_);
  and (_14729_, _10768_, _23830_);
  and (_14730_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or (_07007_, _14730_, _14729_);
  and (_14731_, _26190_, _23848_);
  and (_14732_, _14731_, _25886_);
  not (_14733_, _14731_);
  and (_14734_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_07011_, _14734_, _14732_);
  and (_14735_, _01371_, _26085_);
  and (_14736_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_07013_, _14736_, _14735_);
  and (_14737_, _10670_, _25886_);
  and (_14738_, _10673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_07018_, _14738_, _14737_);
  and (_14739_, _10483_, _26085_);
  and (_14740_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_07020_, _14740_, _14739_);
  and (_14741_, _26351_, _23768_);
  and (_14742_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_07022_, _14742_, _14741_);
  and (_14743_, _06836_, _23830_);
  and (_14744_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or (_07042_, _14744_, _14743_);
  and (_14745_, _10483_, _26170_);
  and (_14746_, _10486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_27018_, _14746_, _14745_);
  and (_14747_, _10420_, _25886_);
  and (_14748_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_07045_, _14748_, _14747_);
  and (_14749_, _06836_, _26242_);
  and (_14750_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_07047_, _14750_, _14749_);
  nand (_14752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _23049_);
  nor (_07049_, _14752_, t2ex_i);
  and (_14753_, _10375_, _23768_);
  and (_14754_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or (_07050_, _14754_, _14753_);
  and (_14755_, _10420_, _26185_);
  and (_14756_, _10423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_07052_, _14756_, _14755_);
  and (_14757_, _14446_, _26242_);
  and (_14758_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_07055_, _14758_, _14757_);
  nor (_14759_, t2_i, rst);
  and (_07057_, _14759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_14760_, _10375_, _23830_);
  and (_14761_, _10378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or (_07059_, _14761_, _14760_);
  and (_14762_, _06836_, _26185_);
  and (_14763_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or (_07063_, _14763_, _14762_);
  and (_14764_, _14446_, _26185_);
  and (_14765_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_07065_, _14765_, _14764_);
  and (_14766_, _09566_, _23830_);
  and (_14767_, _09568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_07067_, _14767_, _14766_);
  nand (_14768_, _09682_, _25417_);
  or (_14769_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_14770_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_14771_, _14770_, _14769_);
  or (_14772_, _14771_, _09682_);
  and (_14773_, _14772_, _23049_);
  and (_07069_, _14773_, _14768_);
  and (_14774_, _09667_, _25927_);
  and (_14775_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_07071_, _14775_, _14774_);
  nand (_14776_, _09679_, _25417_);
  and (_14777_, _09723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_14778_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_14779_, _14778_, _14777_);
  or (_14780_, _14779_, _09679_);
  and (_14781_, _14780_, _09684_);
  and (_14782_, _14781_, _14776_);
  and (_14783_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_14784_, _14783_, _14782_);
  and (_07072_, _14784_, _23049_);
  and (_14785_, _06836_, _26085_);
  and (_14786_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or (_07078_, _14786_, _14785_);
  and (_14787_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_14788_, _26261_, _26242_);
  or (_07086_, _14788_, _14787_);
  and (_14789_, _09756_, _25927_);
  and (_14790_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_07090_, _14790_, _14789_);
  and (_14791_, _23782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_14792_, _26170_, _23780_);
  or (_07093_, _14792_, _14791_);
  and (_14793_, _14702_, _26242_);
  and (_14794_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_27009_, _14794_, _14793_);
  and (_14795_, _09176_, _26185_);
  and (_14796_, _09178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_07100_, _14796_, _14795_);
  and (_14797_, _14702_, _26185_);
  and (_14798_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or (_07101_, _14798_, _14797_);
  and (_14799_, _14702_, _26085_);
  and (_14800_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or (_07135_, _14800_, _14799_);
  and (_14801_, _04055_, _26085_);
  and (_14802_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_07140_, _14802_, _14801_);
  and (_14803_, _04055_, _23830_);
  and (_14804_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_07151_, _14804_, _14803_);
  and (_14805_, _26275_, _25927_);
  and (_14806_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_07153_, _14806_, _14805_);
  and (_14807_, _09170_, _23768_);
  and (_14808_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or (_07156_, _14808_, _14807_);
  and (_14809_, _09170_, _26170_);
  and (_14810_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  or (_07163_, _14810_, _14809_);
  and (_14811_, _04055_, _25886_);
  and (_14812_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_07167_, _14812_, _14811_);
  and (_14813_, _04055_, _26170_);
  and (_14814_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_07170_, _14814_, _14813_);
  and (_14815_, _09170_, _23830_);
  and (_14816_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or (_07177_, _14816_, _14815_);
  and (_14817_, _14446_, _23768_);
  and (_14818_, _14448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_07179_, _14818_, _14817_);
  and (_14819_, _10562_, _25886_);
  and (_14820_, _10565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_07187_, _14820_, _14819_);
  nand (_14821_, _09682_, _25362_);
  not (_14822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_14823_, _09724_, _14822_);
  and (_14824_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_14825_, _14824_, _14823_);
  or (_14826_, _14825_, _09682_);
  and (_14827_, _14826_, _23049_);
  and (_07189_, _14827_, _14821_);
  nand (_14828_, _09682_, _25332_);
  not (_14829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_14830_, _09724_, _14829_);
  and (_14831_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_14832_, _14831_, _14830_);
  or (_14833_, _14832_, _09682_);
  and (_14834_, _14833_, _23049_);
  and (_07198_, _14834_, _14828_);
  nand (_14835_, _09682_, _23824_);
  or (_14836_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_14837_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_14838_, _14837_, _14836_);
  or (_14839_, _14838_, _09682_);
  and (_14840_, _14839_, _23049_);
  and (_07203_, _14840_, _14835_);
  and (_14841_, _14731_, _26170_);
  and (_14842_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_07214_, _14842_, _14841_);
  and (_14843_, _06836_, _23768_);
  and (_14844_, _06838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or (_07237_, _14844_, _14843_);
  and (_14845_, _09170_, _26085_);
  and (_14846_, _09172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or (_07240_, _14846_, _14845_);
  nand (_14847_, _09679_, _25332_);
  nor (_14848_, _09686_, _09350_);
  and (_14849_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_14850_, _14849_, _14848_);
  or (_14851_, _14850_, _09679_);
  and (_14852_, _14851_, _09684_);
  and (_14853_, _14852_, _14847_);
  and (_14854_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_14855_, _14854_, _14853_);
  and (_07244_, _14855_, _23049_);
  and (_14856_, _14702_, _26170_);
  and (_14857_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_07247_, _14857_, _14856_);
  and (_14858_, _07645_, _26185_);
  and (_14859_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_07254_, _14859_, _14858_);
  and (_14860_, _09053_, _23830_);
  and (_14861_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_07255_, _14861_, _14860_);
  and (_14862_, _04055_, _26242_);
  and (_14863_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_27196_, _14863_, _14862_);
  and (_14864_, _14702_, _25927_);
  and (_14865_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_27008_, _14865_, _14864_);
  and (_14866_, _04055_, _26185_);
  and (_14867_, _04057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_07267_, _14867_, _14866_);
  and (_14868_, _14702_, _23768_);
  and (_14869_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or (_07269_, _14869_, _14868_);
  and (_14870_, _09053_, _25886_);
  and (_14871_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_07272_, _14871_, _14870_);
  and (_14872_, _14731_, _25927_);
  and (_14873_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_07275_, _14873_, _14872_);
  and (_14874_, _14629_, _26170_);
  and (_14875_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_07277_, _14875_, _14874_);
  or (_14876_, _09684_, _25258_);
  and (_14877_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_14878_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_14879_, _14878_, _14877_);
  or (_14880_, _14879_, _09682_);
  and (_14881_, _14880_, _23049_);
  and (_07279_, _14881_, _14876_);
  and (_14882_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_14883_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_14884_, _14883_, _14882_);
  or (_14885_, _14884_, _09682_);
  nand (_14886_, _09682_, _25279_);
  and (_14887_, _14886_, _23049_);
  and (_07282_, _14887_, _14885_);
  or (_14888_, _09724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_14889_, _09725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_14890_, _14889_, _14888_);
  or (_14891_, _14890_, _09682_);
  nand (_14892_, _09682_, _23761_);
  and (_14893_, _14892_, _23049_);
  and (_07284_, _14893_, _14891_);
  and (_14894_, _07645_, _26242_);
  and (_14895_, _07647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_07290_, _14895_, _14894_);
  and (_14896_, _09152_, _25927_);
  and (_14897_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_27153_, _14897_, _14896_);
  and (_14898_, _02329_, _25927_);
  and (_14899_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_07296_, _14899_, _14898_);
  and (_14900_, _09152_, _26170_);
  and (_14901_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_07304_, _14901_, _14900_);
  and (_14902_, _26275_, _26242_);
  and (_14903_, _26277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_07307_, _14903_, _14902_);
  and (_14904_, _09152_, _26085_);
  and (_14905_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_07314_, _14905_, _14904_);
  and (_14906_, _26150_, _23848_);
  and (_14907_, _14906_, _25927_);
  not (_14908_, _14906_);
  and (_14909_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_07319_, _14909_, _14907_);
  nand (_14910_, _09679_, _25279_);
  nor (_14911_, _09686_, _09059_);
  and (_14912_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_14913_, _14912_, _14911_);
  or (_14914_, _14913_, _09679_);
  and (_14915_, _14914_, _09684_);
  and (_14916_, _14915_, _14910_);
  and (_14917_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_14918_, _14917_, _14916_);
  and (_07327_, _14918_, _23049_);
  nand (_14919_, _09679_, _23824_);
  not (_14920_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_14921_, _09686_, _14920_);
  and (_14922_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_14923_, _14922_, _14921_);
  or (_14924_, _14923_, _09679_);
  and (_14925_, _14924_, _09684_);
  and (_14926_, _14925_, _14919_);
  and (_14927_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_14928_, _14927_, _14926_);
  and (_07331_, _14928_, _23049_);
  nand (_14929_, _09679_, _25160_);
  not (_14930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor (_14931_, _09686_, _14930_);
  and (_14932_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_14933_, _14932_, _14931_);
  or (_14934_, _14933_, _09679_);
  and (_14935_, _14934_, _09684_);
  and (_14936_, _14935_, _14929_);
  and (_14937_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_14938_, _14937_, _14936_);
  and (_07334_, _14938_, _23049_);
  and (_14939_, _09723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_14940_, _09686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_14941_, _14940_, _14939_);
  nor (_14942_, _14941_, _09679_);
  and (_14943_, _09679_, _25258_);
  or (_14944_, _14943_, _14942_);
  and (_14945_, _14944_, _09684_);
  and (_14946_, _09682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_14947_, _14946_, _14945_);
  and (_07336_, _14947_, _23049_);
  and (_14948_, _14906_, _25886_);
  and (_14949_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_07357_, _14949_, _14948_);
  and (_14950_, _14702_, _25886_);
  and (_14951_, _14704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or (_07359_, _14951_, _14950_);
  and (_14952_, _04085_, _23830_);
  and (_14953_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_07364_, _14953_, _14952_);
  and (_14954_, _04085_, _25886_);
  and (_14955_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_07367_, _14955_, _14954_);
  and (_14956_, _14906_, _26170_);
  and (_14957_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_07369_, _14957_, _14956_);
  and (_14958_, _09152_, _26185_);
  and (_14959_, _09154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_07382_, _14959_, _14958_);
  and (_14960_, _09140_, _23768_);
  and (_14961_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or (_07392_, _14961_, _14960_);
  and (_14962_, _14450_, _26170_);
  and (_14963_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_07397_, _14963_, _14962_);
  and (_14964_, _14450_, _25886_);
  and (_14965_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_27007_, _14965_, _14964_);
  and (_14966_, _09667_, _26185_);
  and (_14967_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_27029_, _14967_, _14966_);
  and (_14968_, _09667_, _23830_);
  and (_14969_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_07410_, _14969_, _14968_);
  and (_14970_, _00256_, _25126_);
  not (_14971_, _14970_);
  or (_14972_, _14971_, _25053_);
  or (_14973_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_14974_, _14973_, _25128_);
  and (_14975_, _14974_, _14972_);
  and (_14976_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_14977_, _25627_, _25617_);
  and (_14978_, _14977_, _25536_);
  nand (_14979_, _14978_, _23729_);
  or (_14980_, _14978_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_14981_, _14980_, _25618_);
  and (_14982_, _14981_, _14979_);
  or (_14983_, _14982_, _14976_);
  or (_14984_, _14983_, _14975_);
  and (_07414_, _14984_, _23049_);
  and (_14985_, _09667_, _25886_);
  and (_14986_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_07416_, _14986_, _14985_);
  and (_14987_, _09140_, _25927_);
  and (_14988_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or (_07422_, _14988_, _14987_);
  and (_14989_, _04085_, _26242_);
  and (_14990_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_07427_, _14990_, _14989_);
  and (_14991_, _26175_, _26072_);
  and (_14992_, _14991_, _25886_);
  not (_14993_, _14991_);
  and (_14994_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_07429_, _14994_, _14992_);
  and (_14995_, _09140_, _23830_);
  and (_14996_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  or (_07431_, _14996_, _14995_);
  and (_14997_, _04085_, _26185_);
  and (_14998_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_07433_, _14998_, _14997_);
  and (_14999_, _26175_, _25932_);
  and (_15000_, _14999_, _26242_);
  not (_15001_, _14999_);
  and (_15002_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_07438_, _15002_, _15000_);
  and (_15003_, _04085_, _26085_);
  and (_15004_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_27195_, _15004_, _15003_);
  and (_15005_, _09140_, _26185_);
  and (_15006_, _09142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or (_27156_, _15006_, _15005_);
  and (_15007_, _14999_, _25927_);
  and (_15008_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_07458_, _15008_, _15007_);
  and (_15009_, _26340_, _26175_);
  and (_15010_, _15009_, _26185_);
  not (_15011_, _15009_);
  and (_15012_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_07463_, _15012_, _15010_);
  and (_15013_, _14450_, _26085_);
  and (_15014_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or (_07465_, _15014_, _15013_);
  and (_15015_, _15009_, _25927_);
  and (_15016_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_07469_, _15016_, _15015_);
  and (_15017_, _26421_, _26175_);
  and (_15018_, _15017_, _26185_);
  not (_15019_, _15017_);
  and (_15020_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_07472_, _15020_, _15018_);
  and (_15021_, _04198_, _26085_);
  and (_15022_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_07474_, _15022_, _15021_);
  and (_15023_, _15017_, _26170_);
  and (_15024_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_07477_, _15024_, _15023_);
  and (_15025_, _04198_, _26242_);
  and (_15026_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_07480_, _15026_, _15025_);
  and (_15027_, _14906_, _26242_);
  and (_15028_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_27266_, _15028_, _15027_);
  and (_15029_, _26175_, _26150_);
  and (_15031_, _15029_, _26242_);
  not (_15032_, _15029_);
  and (_15033_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_26959_, _15033_, _15031_);
  and (_15034_, _04198_, _26185_);
  and (_15035_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or (_27193_, _15035_, _15034_);
  and (_15036_, _14456_, _25886_);
  and (_15037_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_07489_, _15037_, _15036_);
  and (_15038_, _14456_, _26085_);
  and (_15039_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_07493_, _15039_, _15038_);
  and (_15040_, _15029_, _25927_);
  and (_15041_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_07497_, _15041_, _15040_);
  and (_15042_, _14456_, _23830_);
  and (_15043_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_07499_, _15043_, _15042_);
  and (_15044_, _26224_, _26175_);
  and (_15045_, _15044_, _23830_);
  not (_15046_, _15044_);
  and (_15047_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_07502_, _15047_, _15045_);
  and (_15048_, _15044_, _26170_);
  and (_15049_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_07504_, _15049_, _15048_);
  and (_15050_, _26175_, _23847_);
  and (_15051_, _15050_, _25927_);
  not (_15052_, _15050_);
  and (_15053_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_07507_, _15053_, _15051_);
  and (_15054_, _26258_, _26175_);
  and (_15055_, _15054_, _26185_);
  not (_15056_, _15054_);
  and (_15057_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_07514_, _15057_, _15055_);
  and (_15058_, _15054_, _23830_);
  and (_15059_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_07516_, _15059_, _15058_);
  and (_15060_, _09756_, _23768_);
  and (_15061_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_07519_, _15061_, _15060_);
  and (_15062_, _15054_, _23768_);
  and (_15063_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_07521_, _15063_, _15062_);
  and (_15064_, _26374_, _26175_);
  and (_15065_, _15064_, _26185_);
  not (_15066_, _15064_);
  and (_15067_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_07524_, _15067_, _15065_);
  and (_15069_, _09756_, _26170_);
  and (_15070_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_07530_, _15070_, _15069_);
  and (_15071_, _26446_, _26185_);
  and (_15072_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_07532_, _15072_, _15071_);
  and (_15073_, _14456_, _26242_);
  and (_15074_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_07535_, _15074_, _15073_);
  and (_15075_, _00049_, _23768_);
  and (_15076_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_07547_, _15076_, _15075_);
  and (_15077_, _04085_, _25927_);
  and (_15078_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_07549_, _15078_, _15077_);
  and (_15079_, _14450_, _23768_);
  and (_15080_, _14452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or (_07551_, _15080_, _15079_);
  and (_15081_, _26283_, _26175_);
  and (_15083_, _15081_, _26185_);
  not (_15084_, _15081_);
  and (_15085_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_07554_, _15085_, _15083_);
  and (_15086_, _15081_, _25886_);
  and (_15087_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_26956_, _15087_, _15086_);
  and (_15088_, _04085_, _23768_);
  and (_15089_, _04087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_27194_, _15089_, _15088_);
  and (_15090_, _15050_, _26085_);
  and (_15091_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_26954_, _15091_, _15090_);
  and (_15092_, _15081_, _23768_);
  and (_15093_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_07581_, _15093_, _15092_);
  and (_15094_, _14380_, _26185_);
  and (_15095_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_07583_, _15095_, _15094_);
  and (_15096_, _14991_, _26085_);
  and (_15097_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_07597_, _15097_, _15096_);
  and (_15098_, _14380_, _26085_);
  and (_15099_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_07600_, _15099_, _15098_);
  and (_15100_, _14380_, _23830_);
  and (_15101_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_07602_, _15101_, _15100_);
  and (_15102_, _04092_, _26242_);
  and (_15103_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or (_07828_, _15103_, _15102_);
  and (_15104_, _04092_, _26185_);
  and (_15105_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or (_07832_, _15105_, _15104_);
  and (_15106_, _14380_, _26242_);
  and (_15107_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_27004_, _15107_, _15106_);
  and (_15108_, _14456_, _23768_);
  and (_15109_, _14458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_27005_, _15109_, _15108_);
  and (_15110_, _15044_, _26185_);
  and (_15111_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_07844_, _15111_, _15110_);
  and (_15112_, _04198_, _25927_);
  and (_15113_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or (_07846_, _15113_, _15112_);
  and (_15114_, _26215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  and (_15115_, _26242_, _26214_);
  or (_07849_, _15115_, _15114_);
  and (_15116_, _15050_, _25886_);
  and (_15117_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_07851_, _15117_, _15116_);
  and (_15118_, _14384_, _26242_);
  and (_15119_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_07854_, _15119_, _15118_);
  and (_15120_, _14384_, _26185_);
  and (_15121_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_07857_, _15121_, _15120_);
  and (_15122_, _15064_, _25886_);
  and (_15123_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_07896_, _15123_, _15122_);
  and (_15124_, _15050_, _26242_);
  and (_15125_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_26955_, _15125_, _15124_);
  and (_15126_, _14999_, _26170_);
  and (_15127_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_26963_, _15127_, _15126_);
  and (_15128_, _15009_, _26170_);
  and (_15129_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_07904_, _15129_, _15128_);
  and (_15130_, _15017_, _25886_);
  and (_15131_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_07906_, _15131_, _15130_);
  and (_15132_, _04825_, _23830_);
  and (_15133_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or (_07909_, _15133_, _15132_);
  and (_15134_, _15064_, _26242_);
  and (_15135_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_07912_, _15135_, _15134_);
  and (_15136_, _15064_, _23768_);
  and (_15137_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_07913_, _15137_, _15136_);
  and (_15138_, _15081_, _26242_);
  and (_15139_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_07915_, _15139_, _15138_);
  and (_15140_, _15029_, _23830_);
  and (_15141_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_07919_, _15141_, _15140_);
  and (_15142_, _15009_, _25886_);
  and (_15143_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_07925_, _15143_, _15142_);
  and (_15144_, _04301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_15145_, _04300_, _23768_);
  or (_07929_, _15145_, _15144_);
  and (_15146_, _26355_, _26190_);
  and (_15147_, _15146_, _26185_);
  not (_15148_, _15146_);
  and (_15149_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_07932_, _15149_, _15147_);
  and (_15150_, _02329_, _26170_);
  and (_15152_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_27276_, _15152_, _15150_);
  and (_15153_, _26615_, _26242_);
  and (_15154_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_07936_, _15154_, _15153_);
  and (_15155_, _26615_, _25927_);
  and (_15156_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_07939_, _15156_, _15155_);
  and (_15157_, _26308_, _25886_);
  and (_15158_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_07942_, _15158_, _15157_);
  and (_15159_, _26185_, _23849_);
  and (_15160_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_07946_, _15160_, _15159_);
  and (_15161_, _12650_, _23830_);
  and (_15162_, _12652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or (_07947_, _15162_, _15161_);
  and (_15163_, _26329_, _23768_);
  and (_15164_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_07949_, _15164_, _15163_);
  and (_15166_, _01989_, _25886_);
  and (_15167_, _01991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_07952_, _15167_, _15166_);
  and (_15168_, _04198_, _26170_);
  and (_15169_, _04200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or (_27192_, _15169_, _15168_);
  and (_15170_, _14384_, _26085_);
  and (_15171_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or (_08188_, _15171_, _15170_);
  and (_15172_, _10404_, _26185_);
  and (_15173_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_27256_, _15173_, _15172_);
  and (_15174_, _02519_, _26085_);
  and (_15175_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_08195_, _15175_, _15174_);
  and (_15176_, _14380_, _23768_);
  and (_15177_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_27003_, _15177_, _15176_);
  and (_15178_, _14380_, _26170_);
  and (_15179_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_08198_, _15179_, _15178_);
  and (_15181_, _14380_, _25927_);
  and (_15182_, _14382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_08201_, _15182_, _15181_);
  and (_15183_, _04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_15184_, _04120_, _25927_);
  or (_08207_, _15184_, _15183_);
  and (_15185_, _04092_, _25927_);
  and (_15186_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or (_08209_, _15186_, _15185_);
  and (_15187_, _04092_, _23768_);
  and (_15188_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or (_08213_, _15188_, _15187_);
  and (_15189_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  and (_15190_, _04143_, _23830_);
  or (_08221_, _15190_, _15189_);
  and (_15191_, _10475_, _26242_);
  and (_15192_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_27247_, _15192_, _15191_);
  nand (_15193_, _22830_, _22738_);
  or (_15194_, _22738_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_15195_, _15194_, _23049_);
  and (_26896_[0], _15195_, _15193_);
  and (_15196_, _01873_, _22992_);
  or (_15197_, _15196_, _23023_);
  and (_15198_, _22992_, _22989_);
  and (_15199_, _24164_, _23022_);
  or (_15200_, _15199_, _15198_);
  and (_15201_, _22992_, _24143_);
  or (_15202_, _15201_, _15200_);
  or (_15203_, _15202_, _15197_);
  not (_15204_, _23055_);
  and (_15205_, _01873_, _22982_);
  or (_15206_, _15205_, _15204_);
  or (_15207_, _15206_, _15203_);
  and (_15208_, _15207_, _01913_);
  nor (_15209_, _23055_, _23040_);
  and (_15210_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_15211_, _15210_, _15209_);
  and (_15212_, _15211_, _23049_);
  or (_26904_[1], _15212_, _15208_);
  or (_15213_, _09643_, _09629_);
  or (_15214_, _15213_, _09646_);
  or (_15215_, _15214_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_15216_, _15215_, _09661_);
  nor (_15217_, _09659_, _22942_);
  or (_15218_, _15217_, rst);
  or (_26895_[0], _15218_, _15216_);
  and (_26893_[0], _23046_, _23049_);
  and (_26893_[1], _25119_, _23049_);
  and (_15219_, _02512_, _23768_);
  and (_15220_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_08308_, _15220_, _15219_);
  and (_15221_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  and (_15222_, _02010_, _26085_);
  or (_08310_, _15222_, _15221_);
  and (_15223_, _02512_, _25927_);
  and (_15224_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_08313_, _15224_, _15223_);
  and (_15225_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  and (_15226_, _02010_, _26185_);
  or (_08316_, _15226_, _15225_);
  and (_15227_, _02329_, _23830_);
  and (_15228_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_08328_, _15228_, _15227_);
  and (_15229_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  and (_15230_, _02010_, _26242_);
  or (_08348_, _15230_, _15229_);
  and (_15231_, _26258_, _25938_);
  and (_15232_, _15231_, _23768_);
  not (_15233_, _15231_);
  and (_15234_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_08360_, _15234_, _15232_);
  and (_15235_, _15231_, _25927_);
  and (_15236_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_27237_, _15236_, _15235_);
  and (_15237_, _00049_, _26242_);
  and (_15238_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_08389_, _15238_, _15237_);
  or (_15239_, _22804_, _00137_);
  or (_15241_, _22738_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_15242_, _15241_, _23049_);
  and (_26896_[3], _15242_, _15239_);
  nand (_15243_, _08650_, _01913_);
  not (_15244_, _22862_);
  or (_15245_, _05550_, _15244_);
  and (_26894_[1], _15245_, _15243_);
  or (_15246_, _22777_, _00137_);
  or (_15247_, _22738_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_15248_, _15247_, _23049_);
  and (_26896_[2], _15248_, _15246_);
  and (_15249_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_15250_, _04820_, _26185_);
  or (_08400_, _15250_, _15249_);
  nand (_26894_[0], _08653_, _01913_);
  and (_15251_, _01871_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_15252_, _01907_, _23004_);
  and (_15253_, _22982_, _22862_);
  or (_15254_, _15253_, _22977_);
  and (_15255_, _15205_, _22836_);
  not (_15257_, _24154_);
  nand (_15258_, _15257_, _24144_);
  or (_15259_, _15258_, _15255_);
  or (_15260_, _15259_, _15254_);
  or (_15261_, _15260_, _15252_);
  or (_15262_, _15261_, _01897_);
  and (_15263_, _15262_, _01913_);
  or (_26899_[1], _15263_, _15251_);
  nand (_15264_, _22855_, _22738_);
  or (_15265_, _22738_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_15266_, _15265_, _23049_);
  and (_26896_[1], _15266_, _15264_);
  and (_15267_, _02011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  and (_15268_, _02010_, _25886_);
  or (_08411_, _15268_, _15267_);
  nor (_15269_, _25074_, _25060_);
  nand (_15270_, _15269_, _25098_);
  and (_15271_, _24151_, _22972_);
  and (_15272_, _15271_, _23007_);
  or (_15273_, _15272_, _01894_);
  or (_15274_, _15273_, _15270_);
  nand (_15275_, _25092_, _25073_);
  or (_15276_, _25087_, _25100_);
  or (_15277_, _15276_, _08639_);
  or (_15278_, _15277_, _15275_);
  or (_15279_, _15278_, _15274_);
  or (_15280_, _03988_, _23021_);
  and (_15281_, _24164_, _23007_);
  or (_15282_, _15281_, _23031_);
  or (_15283_, _15282_, _01907_);
  or (_15284_, _15283_, _15280_);
  and (_15285_, _22972_, _23007_);
  and (_15286_, _15285_, _22989_);
  or (_15287_, _15286_, _22998_);
  or (_15288_, _15287_, _25111_);
  or (_15289_, _25083_, _25080_);
  and (_15290_, _23030_, _24143_);
  or (_15291_, _15290_, _08640_);
  or (_15292_, _15291_, _15289_);
  or (_15293_, _15292_, _15288_);
  or (_15294_, _15293_, _15284_);
  or (_15295_, _15294_, _15279_);
  and (_15296_, _15295_, _22739_);
  and (_15297_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15298_, _24148_, _22944_);
  and (_15299_, _15204_, _08647_);
  or (_15300_, _08643_, _15299_);
  or (_15301_, _15300_, _15298_);
  or (_15302_, _15301_, _15297_);
  or (_15303_, _15302_, _15296_);
  and (_26905_, _15303_, _23049_);
  and (_15304_, _01660_, _02503_);
  nand (_15305_, _15304_, _10271_);
  and (_15306_, _15305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_15307_, _05692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_15308_, _01660_, _01664_);
  or (_15309_, _15308_, _05698_);
  and (_15310_, _15309_, _15307_);
  nor (_15311_, _15310_, _00071_);
  or (_15312_, _15311_, _15306_);
  and (_15313_, _15312_, _00070_);
  nor (_15314_, _00070_, _25362_);
  or (_15315_, _15314_, _15313_);
  and (_08463_, _15315_, _23049_);
  and (_15316_, _26351_, _26170_);
  and (_15317_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_27273_, _15317_, _15316_);
  and (_15318_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_15319_, _04820_, _26242_);
  or (_08478_, _15319_, _15318_);
  and (_15320_, _26615_, _25886_);
  and (_15321_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_08481_, _15321_, _15320_);
  and (_15322_, _02512_, _26185_);
  and (_15323_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_08507_, _15323_, _15322_);
  and (_15324_, _02512_, _26242_);
  and (_15325_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_08511_, _15325_, _15324_);
  and (_15326_, _02512_, _26085_);
  and (_15327_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_08513_, _15327_, _15326_);
  nand (_15328_, _22883_, _22738_);
  or (_15329_, _22738_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_15330_, _15329_, _23049_);
  and (_26896_[5], _15330_, _15328_);
  or (_15331_, _22934_, _00137_);
  or (_15332_, _22738_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_15333_, _15332_, _23049_);
  and (_26896_[6], _15333_, _15331_);
  nand (_15334_, _00069_, _25332_);
  nor (_15335_, _15305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_15336_, _15305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_15337_, _09311_, _01667_);
  and (_15338_, _15337_, _01654_);
  nand (_15339_, _15338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_15340_, _15339_, _00071_);
  or (_15341_, _15340_, _15336_);
  or (_15342_, _15341_, _15335_);
  or (_15343_, _15342_, _00069_);
  and (_15344_, _15343_, _23049_);
  and (_08524_, _15344_, _15334_);
  and (_15345_, _26414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_15346_, _26413_, _23830_);
  or (_08537_, _15346_, _15345_);
  and (_15347_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_15348_, _04820_, _25886_);
  or (_08557_, _15348_, _15347_);
  and (_15349_, _15231_, _26185_);
  and (_15350_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_27241_, _15350_, _15349_);
  and (_15351_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_15352_, _04820_, _23830_);
  or (_27075_, _15352_, _15351_);
  and (_15353_, _15231_, _26242_);
  and (_15354_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_08582_, _15354_, _15353_);
  and (_15355_, _01371_, _26170_);
  and (_15356_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_08588_, _15356_, _15355_);
  and (_15357_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_15358_, _10259_, _26242_);
  or (_08591_, _15358_, _15357_);
  and (_15359_, _02519_, _26170_);
  and (_15360_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_08609_, _15360_, _15359_);
  and (_15361_, _25927_, _23231_);
  and (_15362_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_08612_, _15362_, _15361_);
  and (_15363_, _26185_, _26073_);
  and (_15364_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_08615_, _15364_, _15363_);
  or (_15365_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _22734_);
  and (_15366_, _15365_, _23049_);
  and (_15367_, _15366_, _08655_);
  and (_15368_, _22995_, _24143_);
  or (_15369_, _15368_, _01908_);
  or (_15370_, _15205_, _15196_);
  and (_15371_, _01899_, _22990_);
  and (_15372_, _15285_, _23052_);
  or (_15373_, _15372_, _15371_);
  or (_15374_, _15373_, _15370_);
  and (_15375_, _22994_, _22989_);
  or (_15376_, _15375_, _01874_);
  or (_15377_, _09032_, _03526_);
  or (_15378_, _15377_, _15376_);
  or (_15379_, _15378_, _15374_);
  or (_15380_, _15379_, _15369_);
  or (_15381_, _23018_, _22997_);
  and (_15382_, _15381_, _23052_);
  and (_15383_, _01873_, _23010_);
  or (_15384_, _15383_, _15253_);
  or (_15385_, _15384_, _15200_);
  or (_15386_, _15385_, _15382_);
  and (_15387_, _01898_, _23007_);
  or (_15388_, _15387_, _23034_);
  and (_15389_, _22989_, _22982_);
  or (_15390_, _25082_, _15389_);
  or (_15391_, _15390_, _15388_);
  or (_15392_, _23012_, _22977_);
  or (_15393_, _15392_, _15391_);
  or (_15394_, _15393_, _15386_);
  or (_15395_, _15394_, _15380_);
  and (_15396_, _15395_, _01913_);
  or (_26898_[0], _15396_, _15367_);
  and (_15397_, _14629_, _26242_);
  and (_15398_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_08622_, _15398_, _15397_);
  and (_15399_, _15146_, _23830_);
  and (_15400_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_27278_, _15400_, _15399_);
  and (_15401_, _15231_, _26085_);
  and (_15402_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_27240_, _15402_, _15401_);
  and (_15403_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_15404_, _10259_, _26185_);
  or (_08661_, _15404_, _15403_);
  and (_15405_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_15406_, _10259_, _26085_);
  or (_08665_, _15406_, _15405_);
  and (_15407_, _14906_, _26185_);
  and (_15408_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_08667_, _15408_, _15407_);
  and (_15409_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_15410_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_15411_, _15410_, _15409_);
  and (_15412_, _15411_, _04847_);
  and (_15413_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_15414_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_15415_, _15414_, _15413_);
  and (_15416_, _15415_, _10786_);
  or (_15417_, _15416_, _15412_);
  or (_15418_, _15417_, _10779_);
  and (_15419_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_15420_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_15421_, _15420_, _15419_);
  and (_15422_, _15421_, _04847_);
  and (_15423_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_15424_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_15425_, _15424_, _15423_);
  and (_15426_, _15425_, _10786_);
  or (_15427_, _15426_, _15422_);
  or (_15428_, _15427_, _04870_);
  and (_15429_, _15428_, _10795_);
  and (_15430_, _15429_, _15418_);
  or (_15431_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_15432_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_15433_, _15432_, _15431_);
  and (_15434_, _15433_, _04847_);
  or (_15435_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_15436_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_15437_, _15436_, _15435_);
  and (_15438_, _15437_, _10786_);
  or (_15439_, _15438_, _15434_);
  or (_15440_, _15439_, _10779_);
  or (_15441_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_15442_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_15443_, _15442_, _15441_);
  and (_15444_, _15443_, _04847_);
  or (_15445_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_15446_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_15447_, _15446_, _15445_);
  and (_15448_, _15447_, _10786_);
  or (_15449_, _15448_, _15444_);
  or (_15450_, _15449_, _04870_);
  and (_15451_, _15450_, _04880_);
  and (_15452_, _15451_, _15440_);
  or (_15453_, _15452_, _15430_);
  or (_15454_, _15453_, _10777_);
  and (_15455_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_15456_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_15457_, _15456_, _15455_);
  and (_15458_, _15457_, _04847_);
  and (_15459_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_15460_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_15461_, _15460_, _15459_);
  and (_15462_, _15461_, _10786_);
  or (_15463_, _15462_, _15458_);
  or (_15464_, _15463_, _10779_);
  and (_15465_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_15466_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_15467_, _15466_, _15465_);
  and (_15468_, _15467_, _04847_);
  and (_15469_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_15470_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_15471_, _15470_, _15469_);
  and (_15472_, _15471_, _10786_);
  or (_15473_, _15472_, _15468_);
  or (_15474_, _15473_, _04870_);
  and (_15475_, _15474_, _10795_);
  and (_15476_, _15475_, _15464_);
  or (_15477_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_15478_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_15479_, _15478_, _10786_);
  and (_15480_, _15479_, _15477_);
  or (_15481_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_15482_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_15483_, _15482_, _04847_);
  and (_15484_, _15483_, _15481_);
  or (_15485_, _15484_, _15480_);
  or (_15486_, _15485_, _10779_);
  or (_15487_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_15488_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_15489_, _15488_, _10786_);
  and (_15490_, _15489_, _15487_);
  or (_15491_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_15492_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_15493_, _15492_, _04847_);
  and (_15494_, _15493_, _15491_);
  or (_15495_, _15494_, _15490_);
  or (_15496_, _15495_, _04870_);
  and (_15497_, _15496_, _04880_);
  and (_15498_, _15497_, _15486_);
  or (_15499_, _15498_, _15476_);
  or (_15500_, _15499_, _04851_);
  and (_15501_, _15500_, _10849_);
  and (_15502_, _15501_, _15454_);
  and (_15503_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_15504_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_15505_, _15504_, _15503_);
  and (_15506_, _15505_, _04847_);
  and (_15507_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_15508_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_15509_, _15508_, _15507_);
  and (_15510_, _15509_, _10786_);
  or (_15511_, _15510_, _15506_);
  and (_15512_, _15511_, _04870_);
  and (_15513_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_15514_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_15515_, _15514_, _15513_);
  and (_15516_, _15515_, _04847_);
  and (_15517_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_15518_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_15519_, _15518_, _15517_);
  and (_15520_, _15519_, _10786_);
  or (_15521_, _15520_, _15516_);
  and (_15522_, _15521_, _10779_);
  or (_15523_, _15522_, _04880_);
  or (_15524_, _15523_, _15512_);
  or (_15525_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_15526_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_15527_, _15526_, _10786_);
  and (_15528_, _15527_, _15525_);
  or (_15529_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_15530_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_15531_, _15530_, _04847_);
  and (_15532_, _15531_, _15529_);
  or (_15533_, _15532_, _15528_);
  and (_15534_, _15533_, _04870_);
  or (_15535_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_15536_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_15537_, _15536_, _10786_);
  and (_15538_, _15537_, _15535_);
  or (_15539_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_15540_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_15541_, _15540_, _04847_);
  and (_15542_, _15541_, _15539_);
  or (_15543_, _15542_, _15538_);
  and (_15544_, _15543_, _10779_);
  or (_15545_, _15544_, _10795_);
  or (_15546_, _15545_, _15534_);
  and (_15547_, _15546_, _15524_);
  or (_15548_, _15547_, _04851_);
  and (_15549_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_15550_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_15551_, _15550_, _15549_);
  and (_15552_, _15551_, _04847_);
  and (_15553_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_15554_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_15555_, _15554_, _15553_);
  and (_15556_, _15555_, _10786_);
  or (_15557_, _15556_, _15552_);
  and (_15558_, _15557_, _04870_);
  and (_15559_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_15560_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_15561_, _15560_, _15559_);
  and (_15562_, _15561_, _04847_);
  and (_15563_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_15564_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_15565_, _15564_, _15563_);
  and (_15566_, _15565_, _10786_);
  or (_15567_, _15566_, _15562_);
  and (_15568_, _15567_, _10779_);
  or (_15569_, _15568_, _04880_);
  or (_15570_, _15569_, _15558_);
  or (_15571_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_15572_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_15573_, _15572_, _15571_);
  and (_15574_, _15573_, _04847_);
  or (_15575_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_15576_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_15577_, _15576_, _15575_);
  and (_15578_, _15577_, _10786_);
  or (_15579_, _15578_, _15574_);
  and (_15580_, _15579_, _04870_);
  or (_15581_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_15582_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_15583_, _15582_, _15581_);
  and (_15584_, _15583_, _04847_);
  or (_15585_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_15586_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_15587_, _15586_, _15585_);
  and (_15588_, _15587_, _10786_);
  or (_15589_, _15588_, _15584_);
  and (_15590_, _15589_, _10779_);
  or (_15591_, _15590_, _10795_);
  or (_15592_, _15591_, _15580_);
  and (_15593_, _15592_, _15570_);
  or (_15594_, _15593_, _10777_);
  and (_15595_, _15594_, _04853_);
  and (_15596_, _15595_, _15548_);
  or (_15597_, _15596_, _15502_);
  or (_15598_, _15597_, _04858_);
  and (_15599_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and (_15600_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_15601_, _15600_, _15599_);
  and (_15602_, _15601_, _04847_);
  and (_15603_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  and (_15604_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_15605_, _15604_, _15603_);
  and (_15606_, _15605_, _10786_);
  or (_15607_, _15606_, _15602_);
  and (_15608_, _15607_, _04870_);
  and (_15609_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and (_15610_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_15611_, _15610_, _15609_);
  and (_15612_, _15611_, _04847_);
  and (_15613_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and (_15614_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_15615_, _15614_, _15613_);
  and (_15617_, _15615_, _10786_);
  or (_15618_, _15617_, _15612_);
  and (_15619_, _15618_, _10779_);
  or (_15620_, _15619_, _04880_);
  or (_15621_, _15620_, _15608_);
  or (_15622_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_15623_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and (_15624_, _15623_, _15622_);
  and (_15625_, _15624_, _04847_);
  or (_15626_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_15627_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  and (_15628_, _15627_, _15626_);
  and (_15629_, _15628_, _10786_);
  or (_15630_, _15629_, _15625_);
  and (_15631_, _15630_, _04870_);
  or (_15632_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_15633_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and (_15634_, _15633_, _15632_);
  and (_15635_, _15634_, _04847_);
  or (_15636_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_15638_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and (_15639_, _15638_, _15636_);
  and (_15640_, _15639_, _10786_);
  or (_15641_, _15640_, _15635_);
  and (_15642_, _15641_, _10779_);
  or (_15643_, _15642_, _10795_);
  or (_15644_, _15643_, _15631_);
  and (_15645_, _15644_, _15621_);
  or (_15646_, _15645_, _04851_);
  and (_15647_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_15648_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_15649_, _15648_, _15647_);
  and (_15650_, _15649_, _04847_);
  and (_15651_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_15652_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_15653_, _15652_, _15651_);
  and (_15654_, _15653_, _10786_);
  or (_15655_, _15654_, _15650_);
  and (_15656_, _15655_, _04870_);
  and (_15657_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_15658_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_15659_, _15658_, _15657_);
  and (_15660_, _15659_, _04847_);
  and (_15661_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_15662_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_15663_, _15662_, _15661_);
  and (_15664_, _15663_, _10786_);
  or (_15665_, _15664_, _15660_);
  and (_15666_, _15665_, _10779_);
  or (_15667_, _15666_, _04880_);
  or (_15668_, _15667_, _15656_);
  or (_15669_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_15670_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_15671_, _15670_, _15669_);
  and (_15672_, _15671_, _04847_);
  or (_15673_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_15674_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_15675_, _15674_, _15673_);
  and (_15676_, _15675_, _10786_);
  or (_15677_, _15676_, _15672_);
  and (_15678_, _15677_, _04870_);
  or (_15679_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_15680_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_15681_, _15680_, _15679_);
  and (_15682_, _15681_, _04847_);
  or (_15683_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_15684_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_15685_, _15684_, _15683_);
  and (_15686_, _15685_, _10786_);
  or (_15687_, _15686_, _15682_);
  and (_15688_, _15687_, _10779_);
  or (_15689_, _15688_, _10795_);
  or (_15690_, _15689_, _15678_);
  and (_15691_, _15690_, _15668_);
  or (_15692_, _15691_, _10777_);
  and (_15693_, _15692_, _04853_);
  and (_15694_, _15693_, _15646_);
  and (_15695_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_15696_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_15697_, _15696_, _15695_);
  and (_15698_, _15697_, _10786_);
  and (_15699_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_15700_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_15701_, _15700_, _15699_);
  and (_15702_, _15701_, _04847_);
  or (_15703_, _15702_, _15698_);
  or (_15704_, _15703_, _10779_);
  and (_15705_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_15706_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_15707_, _15706_, _15705_);
  and (_15708_, _15707_, _10786_);
  and (_15709_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_15710_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_15711_, _15710_, _15709_);
  and (_15712_, _15711_, _04847_);
  or (_15713_, _15712_, _15708_);
  or (_15714_, _15713_, _04870_);
  and (_15715_, _15714_, _10795_);
  and (_15716_, _15715_, _15704_);
  or (_15717_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_15718_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_15719_, _15718_, _04847_);
  and (_15720_, _15719_, _15717_);
  or (_15721_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_15722_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_15723_, _15722_, _10786_);
  and (_15724_, _15723_, _15721_);
  or (_15725_, _15724_, _15720_);
  or (_15726_, _15725_, _10779_);
  or (_15727_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_15728_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_15729_, _15728_, _04847_);
  and (_15730_, _15729_, _15727_);
  or (_15731_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_15732_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_15733_, _15732_, _10786_);
  and (_15734_, _15733_, _15731_);
  or (_15735_, _15734_, _15730_);
  or (_15736_, _15735_, _04870_);
  and (_15737_, _15736_, _04880_);
  and (_15738_, _15737_, _15726_);
  or (_15739_, _15738_, _15716_);
  and (_15740_, _15739_, _10777_);
  and (_15741_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_15742_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_15743_, _15742_, _04847_);
  or (_15744_, _15743_, _15741_);
  and (_15745_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_15746_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_15747_, _15746_, _10786_);
  or (_15748_, _15747_, _15745_);
  and (_15749_, _15748_, _15744_);
  or (_15750_, _15749_, _10779_);
  and (_15751_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_15752_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_15753_, _15752_, _04847_);
  or (_15754_, _15753_, _15751_);
  and (_15755_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_15756_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_15757_, _15756_, _10786_);
  or (_15759_, _15757_, _15755_);
  and (_15760_, _15759_, _15754_);
  or (_15761_, _15760_, _04870_);
  and (_15762_, _15761_, _10795_);
  and (_15763_, _15762_, _15750_);
  or (_15764_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_15765_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_15766_, _15765_, _15764_);
  or (_15767_, _15766_, _10786_);
  or (_15768_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_15769_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_15770_, _15769_, _15768_);
  or (_15771_, _15770_, _04847_);
  and (_15772_, _15771_, _15767_);
  or (_15773_, _15772_, _10779_);
  or (_15774_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_15775_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_15776_, _15775_, _15774_);
  or (_15777_, _15776_, _10786_);
  or (_15778_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_15779_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_15780_, _15779_, _15778_);
  or (_15781_, _15780_, _04847_);
  and (_15782_, _15781_, _15777_);
  or (_15783_, _15782_, _04870_);
  and (_15784_, _15783_, _04880_);
  and (_15785_, _15784_, _15773_);
  or (_15786_, _15785_, _15763_);
  and (_15787_, _15786_, _04851_);
  or (_15788_, _15787_, _15740_);
  and (_15789_, _15788_, _10849_);
  or (_15790_, _15789_, _15694_);
  or (_15791_, _15790_, _11038_);
  and (_15792_, _15791_, _15598_);
  or (_15793_, _15792_, _25445_);
  and (_15794_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_15795_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_15796_, _15795_, _15794_);
  and (_15797_, _15796_, _04847_);
  and (_15798_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_15799_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_15800_, _15799_, _15798_);
  and (_15801_, _15800_, _10786_);
  or (_15802_, _15801_, _15797_);
  or (_15803_, _15802_, _10779_);
  and (_15804_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_15805_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_15806_, _15805_, _15804_);
  and (_15807_, _15806_, _04847_);
  and (_15808_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_15809_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_15810_, _15809_, _15808_);
  and (_15811_, _15810_, _10786_);
  or (_15812_, _15811_, _15807_);
  or (_15813_, _15812_, _04870_);
  and (_15814_, _15813_, _10795_);
  and (_15815_, _15814_, _15803_);
  or (_15816_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_15817_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_15818_, _15817_, _15816_);
  and (_15819_, _15818_, _04847_);
  or (_15820_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_15821_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_15822_, _15821_, _15820_);
  and (_15823_, _15822_, _10786_);
  or (_15824_, _15823_, _15819_);
  or (_15825_, _15824_, _10779_);
  or (_15826_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_15827_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_15828_, _15827_, _15826_);
  and (_15829_, _15828_, _04847_);
  or (_15830_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_15831_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_15832_, _15831_, _15830_);
  and (_15833_, _15832_, _10786_);
  or (_15834_, _15833_, _15829_);
  or (_15835_, _15834_, _04870_);
  and (_15836_, _15835_, _04880_);
  and (_15837_, _15836_, _15825_);
  or (_15838_, _15837_, _15815_);
  and (_15840_, _15838_, _04851_);
  and (_15841_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_15842_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_15843_, _15842_, _15841_);
  and (_15844_, _15843_, _04847_);
  and (_15845_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_15846_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_15847_, _15846_, _15845_);
  and (_15848_, _15847_, _10786_);
  or (_15849_, _15848_, _15844_);
  or (_15850_, _15849_, _10779_);
  and (_15851_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_15852_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_15853_, _15852_, _15851_);
  and (_15854_, _15853_, _04847_);
  and (_15855_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_15856_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_15857_, _15856_, _15855_);
  and (_15858_, _15857_, _10786_);
  or (_15859_, _15858_, _15854_);
  or (_15860_, _15859_, _04870_);
  and (_15861_, _15860_, _10795_);
  and (_15862_, _15861_, _15850_);
  or (_15863_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_15864_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_15865_, _15864_, _10786_);
  and (_15866_, _15865_, _15863_);
  or (_15867_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_15868_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_15869_, _15868_, _04847_);
  and (_15870_, _15869_, _15867_);
  or (_15871_, _15870_, _15866_);
  or (_15872_, _15871_, _10779_);
  or (_15873_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_15874_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_15875_, _15874_, _10786_);
  and (_15876_, _15875_, _15873_);
  or (_15877_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_15878_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_15879_, _15878_, _04847_);
  and (_15880_, _15879_, _15877_);
  or (_15881_, _15880_, _15876_);
  or (_15882_, _15881_, _04870_);
  and (_15883_, _15882_, _04880_);
  and (_15884_, _15883_, _15872_);
  or (_15885_, _15884_, _15862_);
  and (_15886_, _15885_, _10777_);
  or (_15887_, _15886_, _15840_);
  and (_15888_, _15887_, _10849_);
  and (_15889_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_15890_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_15891_, _15890_, _15889_);
  and (_15892_, _15891_, _04847_);
  and (_15893_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_15894_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_15895_, _15894_, _15893_);
  and (_15896_, _15895_, _10786_);
  or (_15897_, _15896_, _15892_);
  and (_15898_, _15897_, _04870_);
  and (_15899_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_15900_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_15901_, _15900_, _15899_);
  and (_15902_, _15901_, _04847_);
  and (_15903_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_15904_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_15905_, _15904_, _15903_);
  and (_15906_, _15905_, _10786_);
  or (_15907_, _15906_, _15902_);
  and (_15908_, _15907_, _10779_);
  or (_15909_, _15908_, _15898_);
  and (_15910_, _15909_, _10795_);
  or (_15911_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_15912_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_15913_, _15912_, _10786_);
  and (_15914_, _15913_, _15911_);
  or (_15915_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_15916_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_15917_, _15916_, _04847_);
  and (_15918_, _15917_, _15915_);
  or (_15919_, _15918_, _15914_);
  and (_15920_, _15919_, _04870_);
  or (_15921_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_15922_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_15923_, _15922_, _10786_);
  and (_15924_, _15923_, _15921_);
  or (_15925_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_15926_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_15927_, _15926_, _04847_);
  and (_15928_, _15927_, _15925_);
  or (_15929_, _15928_, _15924_);
  and (_15930_, _15929_, _10779_);
  or (_15931_, _15930_, _15920_);
  and (_15932_, _15931_, _04880_);
  or (_15933_, _15932_, _15910_);
  and (_15934_, _15933_, _10777_);
  and (_15935_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_15936_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_15937_, _15936_, _15935_);
  and (_15938_, _15937_, _04847_);
  and (_15939_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_15940_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_15941_, _15940_, _15939_);
  and (_15942_, _15941_, _10786_);
  or (_15943_, _15942_, _15938_);
  and (_15944_, _15943_, _04870_);
  and (_15945_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_15946_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_15947_, _15946_, _15945_);
  and (_15948_, _15947_, _04847_);
  and (_15949_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_15950_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_15951_, _15950_, _15949_);
  and (_15952_, _15951_, _10786_);
  or (_15953_, _15952_, _15948_);
  and (_15954_, _15953_, _10779_);
  or (_15955_, _15954_, _15944_);
  and (_15956_, _15955_, _10795_);
  or (_15957_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_15958_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_15959_, _15958_, _15957_);
  and (_15960_, _15959_, _04847_);
  or (_15961_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_15962_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_15963_, _15962_, _15961_);
  and (_15964_, _15963_, _10786_);
  or (_15965_, _15964_, _15960_);
  and (_15966_, _15965_, _04870_);
  or (_15967_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_15968_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_15969_, _15968_, _15967_);
  and (_15970_, _15969_, _04847_);
  or (_15971_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_15972_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_15973_, _15972_, _15971_);
  and (_15974_, _15973_, _10786_);
  or (_15975_, _15974_, _15970_);
  and (_15976_, _15975_, _10779_);
  or (_15977_, _15976_, _15966_);
  and (_15978_, _15977_, _04880_);
  or (_15979_, _15978_, _15956_);
  and (_15980_, _15979_, _04851_);
  or (_15981_, _15980_, _15934_);
  and (_15982_, _15981_, _04853_);
  or (_15983_, _15982_, _15888_);
  or (_15984_, _15983_, _04858_);
  and (_15985_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_15986_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_15987_, _15986_, _15985_);
  and (_15988_, _15987_, _04847_);
  and (_15989_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_15991_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_15992_, _15991_, _15989_);
  and (_15993_, _15992_, _10786_);
  or (_15994_, _15993_, _15988_);
  or (_15995_, _15994_, _10779_);
  and (_15996_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_15997_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_15998_, _15997_, _15996_);
  and (_15999_, _15998_, _04847_);
  and (_16000_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_16001_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_16002_, _16001_, _16000_);
  and (_16003_, _16002_, _10786_);
  or (_16004_, _16003_, _15999_);
  or (_16005_, _16004_, _04870_);
  and (_16006_, _16005_, _10795_);
  and (_16007_, _16006_, _15995_);
  or (_16008_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_16009_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_16010_, _16009_, _10786_);
  and (_16011_, _16010_, _16008_);
  or (_16012_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_16013_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_16014_, _16013_, _04847_);
  and (_16015_, _16014_, _16012_);
  or (_16016_, _16015_, _16011_);
  or (_16017_, _16016_, _10779_);
  or (_16018_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_16019_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_16020_, _16019_, _10786_);
  and (_16021_, _16020_, _16018_);
  or (_16022_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_16023_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_16024_, _16023_, _04847_);
  and (_16025_, _16024_, _16022_);
  or (_16026_, _16025_, _16021_);
  or (_16027_, _16026_, _04870_);
  and (_16028_, _16027_, _04880_);
  and (_16029_, _16028_, _16017_);
  or (_16030_, _16029_, _16007_);
  and (_16031_, _16030_, _10777_);
  and (_16032_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_16033_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_16034_, _16033_, _16032_);
  and (_16035_, _16034_, _04847_);
  and (_16036_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_16037_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_16038_, _16037_, _16036_);
  and (_16039_, _16038_, _10786_);
  or (_16040_, _16039_, _16035_);
  or (_16041_, _16040_, _10779_);
  and (_16042_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_16043_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_16044_, _16043_, _16042_);
  and (_16045_, _16044_, _04847_);
  and (_16046_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_16047_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_16048_, _16047_, _16046_);
  and (_16049_, _16048_, _10786_);
  or (_16050_, _16049_, _16045_);
  or (_16051_, _16050_, _04870_);
  and (_16052_, _16051_, _10795_);
  and (_16053_, _16052_, _16041_);
  or (_16054_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_16055_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_16056_, _16055_, _16054_);
  and (_16057_, _16056_, _04847_);
  or (_16058_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_16059_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_16060_, _16059_, _16058_);
  and (_16061_, _16060_, _10786_);
  or (_16062_, _16061_, _16057_);
  or (_16063_, _16062_, _10779_);
  or (_16064_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_16065_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_16066_, _16065_, _16064_);
  and (_16067_, _16066_, _04847_);
  or (_16068_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_16069_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_16070_, _16069_, _16068_);
  and (_16071_, _16070_, _10786_);
  or (_16072_, _16071_, _16067_);
  or (_16073_, _16072_, _04870_);
  and (_16074_, _16073_, _04880_);
  and (_16075_, _16074_, _16063_);
  or (_16076_, _16075_, _16053_);
  and (_16077_, _16076_, _04851_);
  or (_16078_, _16077_, _16031_);
  and (_16079_, _16078_, _10849_);
  or (_16080_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_16081_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_16082_, _16081_, _16080_);
  and (_16083_, _16082_, _04847_);
  or (_16084_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_16085_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_16086_, _16085_, _16084_);
  and (_16087_, _16086_, _10786_);
  or (_16088_, _16087_, _16083_);
  and (_16089_, _16088_, _10779_);
  or (_16090_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_16091_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_16092_, _16091_, _16090_);
  and (_16093_, _16092_, _04847_);
  or (_16094_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_16095_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_16096_, _16095_, _16094_);
  and (_16097_, _16096_, _10786_);
  or (_16098_, _16097_, _16093_);
  and (_16099_, _16098_, _04870_);
  or (_16100_, _16099_, _16089_);
  and (_16101_, _16100_, _04880_);
  and (_16102_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_16103_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_16104_, _16103_, _16102_);
  and (_16105_, _16104_, _04847_);
  and (_16106_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_16107_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_16108_, _16107_, _16106_);
  and (_16109_, _16108_, _10786_);
  or (_16110_, _16109_, _16105_);
  and (_16111_, _16110_, _10779_);
  and (_16112_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_16113_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_16114_, _16113_, _16112_);
  and (_16115_, _16114_, _04847_);
  and (_16116_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_16117_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_16118_, _16117_, _16116_);
  and (_16119_, _16118_, _10786_);
  or (_16120_, _16119_, _16115_);
  and (_16121_, _16120_, _04870_);
  or (_16122_, _16121_, _16111_);
  and (_16123_, _16122_, _10795_);
  or (_16124_, _16123_, _16101_);
  and (_16125_, _16124_, _04851_);
  or (_16126_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_16127_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_16128_, _16127_, _10786_);
  and (_16129_, _16128_, _16126_);
  or (_16130_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_16131_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_16132_, _16131_, _04847_);
  and (_16133_, _16132_, _16130_);
  or (_16134_, _16133_, _16129_);
  and (_16135_, _16134_, _10779_);
  or (_16136_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_16137_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_16138_, _16137_, _10786_);
  and (_16139_, _16138_, _16136_);
  or (_16140_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_16141_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_16142_, _16141_, _04847_);
  and (_16143_, _16142_, _16140_);
  or (_16144_, _16143_, _16139_);
  and (_16145_, _16144_, _04870_);
  or (_16146_, _16145_, _16135_);
  and (_16147_, _16146_, _04880_);
  and (_16148_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_16149_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_16150_, _16149_, _16148_);
  and (_16151_, _16150_, _04847_);
  and (_16152_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_16153_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_16154_, _16153_, _16152_);
  and (_16155_, _16154_, _10786_);
  or (_16156_, _16155_, _16151_);
  and (_16157_, _16156_, _10779_);
  and (_16158_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_16159_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_16160_, _16159_, _16158_);
  and (_16161_, _16160_, _04847_);
  and (_16162_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_16163_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_16164_, _16163_, _16162_);
  and (_16165_, _16164_, _10786_);
  or (_16166_, _16165_, _16161_);
  and (_16167_, _16166_, _04870_);
  or (_16168_, _16167_, _16157_);
  and (_16169_, _16168_, _10795_);
  or (_16170_, _16169_, _16147_);
  and (_16171_, _16170_, _10777_);
  or (_16172_, _16171_, _16125_);
  and (_16173_, _16172_, _04853_);
  or (_16174_, _16173_, _16079_);
  or (_16175_, _16174_, _11038_);
  and (_16176_, _16175_, _15984_);
  or (_16177_, _16176_, _03372_);
  and (_16178_, _16177_, _15793_);
  or (_16179_, _16178_, _04902_);
  or (_16180_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_16181_, _16180_, _23049_);
  and (_08669_, _16181_, _16179_);
  and (_16182_, _09128_, _25927_);
  and (_16183_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  or (_08672_, _16183_, _16182_);
  and (_16184_, _26185_, _26151_);
  and (_16185_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_08675_, _16185_, _16184_);
  and (_16186_, _14558_, _25927_);
  and (_16187_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or (_08677_, _16187_, _16186_);
  and (_16188_, _26151_, _23768_);
  and (_16189_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_27245_, _16189_, _16188_);
  and (_16190_, _26284_, _23830_);
  and (_16191_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_08680_, _16191_, _16190_);
  and (_16192_, _26284_, _25927_);
  and (_16193_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_08682_, _16193_, _16192_);
  and (_16194_, _26225_, _25927_);
  and (_16195_, _26228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_08684_, _16195_, _16194_);
  and (_16196_, _00016_, _23830_);
  and (_16197_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_08686_, _16197_, _16196_);
  and (_16198_, _15146_, _23768_);
  and (_16199_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_08688_, _16199_, _16198_);
  and (_16200_, _26351_, _26185_);
  and (_16201_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_08691_, _16201_, _16200_);
  and (_16202_, _03115_, _23830_);
  and (_16203_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_08693_, _16203_, _16202_);
  and (_16204_, _09053_, _26185_);
  and (_16205_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_08694_, _16205_, _16204_);
  and (_16206_, _14906_, _23768_);
  and (_16207_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_08696_, _16207_, _16206_);
  and (_16208_, _26283_, _23848_);
  and (_16209_, _16208_, _23830_);
  not (_16210_, _16208_);
  and (_16211_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_08699_, _16211_, _16209_);
  and (_16212_, _14388_, _26185_);
  and (_16213_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or (_08701_, _16213_, _16212_);
  and (_16214_, _26329_, _26185_);
  and (_16215_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_27261_, _16215_, _16214_);
  and (_16216_, _02519_, _25886_);
  and (_16217_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_08705_, _16217_, _16216_);
  and (_16218_, _04092_, _23830_);
  and (_16219_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or (_08707_, _16219_, _16218_);
  and (_16220_, _26242_, _25939_);
  and (_16221_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_08709_, _16221_, _16220_);
  and (_16222_, _14731_, _26185_);
  and (_16223_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_08713_, _16223_, _16222_);
  and (_16224_, _14731_, _26085_);
  and (_16225_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_08721_, _16225_, _16224_);
  and (_16226_, _14906_, _26085_);
  and (_16227_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_08724_, _16227_, _16226_);
  and (_16228_, _14558_, _23768_);
  and (_16229_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or (_08733_, _16229_, _16228_);
  and (_16230_, _14731_, _23768_);
  and (_16231_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_08735_, _16231_, _16230_);
  and (_16232_, _26341_, _25927_);
  and (_16233_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_08739_, _16233_, _16232_);
  and (_16234_, _15231_, _26170_);
  and (_16235_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_08741_, _16235_, _16234_);
  and (_16236_, _01568_, _26242_);
  and (_16237_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_08743_, _16237_, _16236_);
  and (_16238_, _01604_, _23830_);
  and (_16239_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_27236_, _16239_, _16238_);
  and (_16240_, _00049_, _25886_);
  and (_16241_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_08746_, _16241_, _16240_);
  and (_16242_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  and (_16243_, _04143_, _26185_);
  or (_08748_, _16243_, _16242_);
  and (_16244_, _04092_, _25886_);
  and (_16245_, _04094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or (_08751_, _16245_, _16244_);
  and (_16246_, _14384_, _26170_);
  and (_16247_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_08753_, _16247_, _16246_);
  and (_16248_, _10455_, _25886_);
  and (_16249_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_08755_, _16249_, _16248_);
  and (_16250_, _14384_, _25927_);
  and (_16251_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_08757_, _16251_, _16250_);
  and (_16252_, _14731_, _23830_);
  and (_16253_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_08759_, _16253_, _16252_);
  and (_16254_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  and (_16255_, _06369_, _25927_);
  or (_08761_, _16255_, _16254_);
  and (_16256_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_16257_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_16258_, _16257_, _16256_);
  and (_16259_, _16258_, _04847_);
  and (_16260_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_16261_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_16262_, _16261_, _16260_);
  and (_16263_, _16262_, _10786_);
  or (_16264_, _16263_, _16259_);
  or (_16265_, _16264_, _10779_);
  and (_16266_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_16267_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_16268_, _16267_, _16266_);
  and (_16269_, _16268_, _04847_);
  and (_16270_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_16271_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_16272_, _16271_, _16270_);
  and (_16273_, _16272_, _10786_);
  or (_16274_, _16273_, _16269_);
  or (_16275_, _16274_, _04870_);
  and (_16276_, _16275_, _10795_);
  and (_16277_, _16276_, _16265_);
  or (_16278_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_16279_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_16280_, _16279_, _16278_);
  and (_16281_, _16280_, _04847_);
  or (_16282_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_16283_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_16284_, _16283_, _16282_);
  and (_16285_, _16284_, _10786_);
  or (_16286_, _16285_, _16281_);
  or (_16287_, _16286_, _10779_);
  or (_16288_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_16289_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_16290_, _16289_, _16288_);
  and (_16291_, _16290_, _04847_);
  or (_16292_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_16293_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_16294_, _16293_, _16292_);
  and (_16295_, _16294_, _10786_);
  or (_16296_, _16295_, _16291_);
  or (_16297_, _16296_, _04870_);
  and (_16298_, _16297_, _04880_);
  and (_16299_, _16298_, _16287_);
  or (_16300_, _16299_, _16277_);
  and (_16301_, _16300_, _04851_);
  and (_16302_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_16303_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_16304_, _16303_, _16302_);
  and (_16305_, _16304_, _04847_);
  and (_16306_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_16307_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_16308_, _16307_, _16306_);
  and (_16309_, _16308_, _10786_);
  or (_16310_, _16309_, _16305_);
  or (_16311_, _16310_, _10779_);
  and (_16312_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_16313_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_16314_, _16313_, _16312_);
  and (_16315_, _16314_, _04847_);
  and (_16316_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_16317_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_16318_, _16317_, _16316_);
  and (_16319_, _16318_, _10786_);
  or (_16320_, _16319_, _16315_);
  or (_16321_, _16320_, _04870_);
  and (_16322_, _16321_, _10795_);
  and (_16323_, _16322_, _16311_);
  or (_16324_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_16325_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_16326_, _16325_, _10786_);
  and (_16327_, _16326_, _16324_);
  or (_16328_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_16329_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_16330_, _16329_, _04847_);
  and (_16331_, _16330_, _16328_);
  or (_16332_, _16331_, _16327_);
  or (_16333_, _16332_, _10779_);
  or (_16334_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_16335_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_16336_, _16335_, _10786_);
  and (_16337_, _16336_, _16334_);
  or (_16338_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_16339_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_16340_, _16339_, _04847_);
  and (_16341_, _16340_, _16338_);
  or (_16342_, _16341_, _16337_);
  or (_16343_, _16342_, _04870_);
  and (_16344_, _16343_, _04880_);
  and (_16345_, _16344_, _16333_);
  or (_16346_, _16345_, _16323_);
  and (_16347_, _16346_, _10777_);
  or (_16348_, _16347_, _16301_);
  and (_16349_, _16348_, _10849_);
  and (_16350_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_16351_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_16352_, _16351_, _16350_);
  and (_16353_, _16352_, _04847_);
  and (_16354_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_16355_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_16356_, _16355_, _16354_);
  and (_16357_, _16356_, _10786_);
  or (_16358_, _16357_, _16353_);
  and (_16359_, _16358_, _04870_);
  and (_16360_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_16361_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_16362_, _16361_, _16360_);
  and (_16363_, _16362_, _04847_);
  and (_16364_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_16365_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_16366_, _16365_, _16364_);
  and (_16367_, _16366_, _10786_);
  or (_16368_, _16367_, _16363_);
  and (_16369_, _16368_, _10779_);
  or (_16370_, _16369_, _16359_);
  and (_16371_, _16370_, _10795_);
  or (_16372_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_16373_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_16374_, _16373_, _10786_);
  and (_16375_, _16374_, _16372_);
  or (_16376_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_16377_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_16378_, _16377_, _04847_);
  and (_16379_, _16378_, _16376_);
  or (_16380_, _16379_, _16375_);
  and (_16381_, _16380_, _04870_);
  or (_16382_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_16383_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_16384_, _16383_, _10786_);
  and (_16385_, _16384_, _16382_);
  or (_16386_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_16387_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_16388_, _16387_, _04847_);
  and (_16389_, _16388_, _16386_);
  or (_16390_, _16389_, _16385_);
  and (_16391_, _16390_, _10779_);
  or (_16392_, _16391_, _16381_);
  and (_16393_, _16392_, _04880_);
  or (_16394_, _16393_, _16371_);
  and (_16395_, _16394_, _10777_);
  and (_16396_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_16397_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_16398_, _16397_, _16396_);
  and (_16399_, _16398_, _04847_);
  and (_16400_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_16401_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_16402_, _16401_, _16400_);
  and (_16403_, _16402_, _10786_);
  or (_16404_, _16403_, _16399_);
  and (_16405_, _16404_, _04870_);
  and (_16406_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_16407_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_16408_, _16407_, _16406_);
  and (_16409_, _16408_, _04847_);
  and (_16410_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_16411_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_16412_, _16411_, _16410_);
  and (_16413_, _16412_, _10786_);
  or (_16414_, _16413_, _16409_);
  and (_16415_, _16414_, _10779_);
  or (_16416_, _16415_, _16405_);
  and (_16417_, _16416_, _10795_);
  or (_16418_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_16419_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_16420_, _16419_, _16418_);
  and (_16421_, _16420_, _04847_);
  or (_16422_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_16423_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_16424_, _16423_, _16422_);
  and (_16425_, _16424_, _10786_);
  or (_16426_, _16425_, _16421_);
  and (_16427_, _16426_, _04870_);
  or (_16428_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_16429_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_16430_, _16429_, _16428_);
  and (_16431_, _16430_, _04847_);
  or (_16432_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_16433_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_16434_, _16433_, _16432_);
  and (_16435_, _16434_, _10786_);
  or (_16436_, _16435_, _16431_);
  and (_16437_, _16436_, _10779_);
  or (_16438_, _16437_, _16427_);
  and (_16439_, _16438_, _04880_);
  or (_16440_, _16439_, _16417_);
  and (_16441_, _16440_, _04851_);
  or (_16442_, _16441_, _16395_);
  and (_16443_, _16442_, _04853_);
  or (_16444_, _16443_, _16349_);
  or (_16445_, _16444_, _04858_);
  and (_16446_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_16447_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_16448_, _16447_, _16446_);
  and (_16449_, _16448_, _04847_);
  and (_16450_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_16451_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_16452_, _16451_, _16450_);
  and (_16453_, _16452_, _10786_);
  or (_16455_, _16453_, _16449_);
  or (_16456_, _16455_, _10779_);
  and (_16457_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_16458_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_16459_, _16458_, _16457_);
  and (_16460_, _16459_, _04847_);
  and (_16461_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_16462_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_16463_, _16462_, _16461_);
  and (_16464_, _16463_, _10786_);
  or (_16465_, _16464_, _16460_);
  or (_16466_, _16465_, _04870_);
  and (_16467_, _16466_, _10795_);
  and (_16468_, _16467_, _16456_);
  or (_16469_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_16470_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_16471_, _16470_, _10786_);
  and (_16472_, _16471_, _16469_);
  or (_16473_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_16474_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_16475_, _16474_, _04847_);
  and (_16476_, _16475_, _16473_);
  or (_16477_, _16476_, _16472_);
  or (_16478_, _16477_, _10779_);
  or (_16479_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_16480_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_16481_, _16480_, _10786_);
  and (_16482_, _16481_, _16479_);
  or (_16483_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_16484_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_16485_, _16484_, _04847_);
  and (_16486_, _16485_, _16483_);
  or (_16487_, _16486_, _16482_);
  or (_16488_, _16487_, _04870_);
  and (_16489_, _16488_, _04880_);
  and (_16490_, _16489_, _16478_);
  or (_16491_, _16490_, _16468_);
  and (_16492_, _16491_, _10777_);
  and (_16493_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_16494_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_16495_, _16494_, _16493_);
  and (_16496_, _16495_, _04847_);
  and (_16497_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_16498_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_16499_, _16498_, _16497_);
  and (_16500_, _16499_, _10786_);
  or (_16501_, _16500_, _16496_);
  or (_16502_, _16501_, _10779_);
  and (_16503_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_16504_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_16505_, _16504_, _16503_);
  and (_16506_, _16505_, _04847_);
  and (_16507_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_16508_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_16509_, _16508_, _16507_);
  and (_16510_, _16509_, _10786_);
  or (_16511_, _16510_, _16506_);
  or (_16512_, _16511_, _04870_);
  and (_16513_, _16512_, _10795_);
  and (_16514_, _16513_, _16502_);
  or (_16515_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_16516_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_16517_, _16516_, _16515_);
  and (_16518_, _16517_, _04847_);
  or (_16519_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_16520_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_16521_, _16520_, _16519_);
  and (_16522_, _16521_, _10786_);
  or (_16523_, _16522_, _16518_);
  or (_16524_, _16523_, _10779_);
  or (_16525_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_16526_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_16527_, _16526_, _16525_);
  and (_16528_, _16527_, _04847_);
  or (_16529_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_16530_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_16531_, _16530_, _16529_);
  and (_16532_, _16531_, _10786_);
  or (_16533_, _16532_, _16528_);
  or (_16534_, _16533_, _04870_);
  and (_16535_, _16534_, _04880_);
  and (_16536_, _16535_, _16524_);
  or (_16537_, _16536_, _16514_);
  and (_16538_, _16537_, _04851_);
  or (_16539_, _16538_, _16492_);
  and (_16540_, _16539_, _10849_);
  or (_16541_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_16542_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_16543_, _16542_, _16541_);
  and (_16544_, _16543_, _04847_);
  or (_16545_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_16546_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_16547_, _16546_, _16545_);
  and (_16548_, _16547_, _10786_);
  or (_16549_, _16548_, _16544_);
  and (_16550_, _16549_, _10779_);
  or (_16551_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_16552_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_16553_, _16552_, _16551_);
  and (_16554_, _16553_, _04847_);
  or (_16555_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_16556_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_16557_, _16556_, _16555_);
  and (_16558_, _16557_, _10786_);
  or (_16559_, _16558_, _16554_);
  and (_16560_, _16559_, _04870_);
  or (_16561_, _16560_, _16550_);
  and (_16562_, _16561_, _04880_);
  and (_16563_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_16564_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_16565_, _16564_, _16563_);
  and (_16566_, _16565_, _04847_);
  and (_16567_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_16568_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_16569_, _16568_, _16567_);
  and (_16570_, _16569_, _10786_);
  or (_16571_, _16570_, _16566_);
  and (_16572_, _16571_, _10779_);
  and (_16573_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_16574_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_16575_, _16574_, _16573_);
  and (_16576_, _16575_, _04847_);
  and (_16577_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_16578_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_16579_, _16578_, _16577_);
  and (_16580_, _16579_, _10786_);
  or (_16581_, _16580_, _16576_);
  and (_16582_, _16581_, _04870_);
  or (_16583_, _16582_, _16572_);
  and (_16584_, _16583_, _10795_);
  or (_16585_, _16584_, _16562_);
  and (_16586_, _16585_, _04851_);
  or (_16587_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_16588_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_16589_, _16588_, _10786_);
  and (_16590_, _16589_, _16587_);
  or (_16591_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_16592_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_16593_, _16592_, _04847_);
  and (_16594_, _16593_, _16591_);
  or (_16595_, _16594_, _16590_);
  and (_16596_, _16595_, _10779_);
  or (_16597_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_16598_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_16599_, _16598_, _10786_);
  and (_16600_, _16599_, _16597_);
  or (_16601_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_16602_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_16603_, _16602_, _04847_);
  and (_16604_, _16603_, _16601_);
  or (_16606_, _16604_, _16600_);
  and (_16607_, _16606_, _04870_);
  or (_16608_, _16607_, _16596_);
  and (_16609_, _16608_, _04880_);
  and (_16610_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_16611_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_16612_, _16611_, _16610_);
  and (_16613_, _16612_, _04847_);
  and (_16614_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_16615_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_16616_, _16615_, _16614_);
  and (_16617_, _16616_, _10786_);
  or (_16618_, _16617_, _16613_);
  and (_16619_, _16618_, _10779_);
  and (_16620_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_16621_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_16622_, _16621_, _16620_);
  and (_16623_, _16622_, _04847_);
  and (_16624_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_16625_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_16626_, _16625_, _16624_);
  and (_16627_, _16626_, _10786_);
  or (_16628_, _16627_, _16623_);
  and (_16629_, _16628_, _04870_);
  or (_16630_, _16629_, _16619_);
  and (_16631_, _16630_, _10795_);
  or (_16632_, _16631_, _16609_);
  and (_16633_, _16632_, _10777_);
  or (_16634_, _16633_, _16586_);
  and (_16635_, _16634_, _04853_);
  or (_16636_, _16635_, _16540_);
  or (_16637_, _16636_, _11038_);
  and (_16638_, _16637_, _16445_);
  or (_16639_, _16638_, _25445_);
  and (_16640_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_16641_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_16642_, _16641_, _16640_);
  and (_16643_, _16642_, _04847_);
  and (_16644_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_16645_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_16647_, _16645_, _16644_);
  and (_16648_, _16647_, _10786_);
  or (_16649_, _16648_, _16643_);
  and (_16650_, _16649_, _04870_);
  and (_16651_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_16652_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_16653_, _16652_, _16651_);
  and (_16654_, _16653_, _04847_);
  and (_16655_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_16656_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_16657_, _16656_, _16655_);
  and (_16658_, _16657_, _10786_);
  or (_16659_, _16658_, _16654_);
  and (_16660_, _16659_, _10779_);
  or (_16661_, _16660_, _16650_);
  and (_16662_, _16661_, _10795_);
  or (_16663_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_16664_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_16665_, _16664_, _10786_);
  and (_16666_, _16665_, _16663_);
  or (_16667_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_16668_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_16669_, _16668_, _04847_);
  and (_16670_, _16669_, _16667_);
  or (_16671_, _16670_, _16666_);
  and (_16672_, _16671_, _04870_);
  or (_16673_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_16674_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_16675_, _16674_, _10786_);
  and (_16676_, _16675_, _16673_);
  or (_16677_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_16678_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_16679_, _16678_, _04847_);
  and (_16680_, _16679_, _16677_);
  or (_16681_, _16680_, _16676_);
  and (_16682_, _16681_, _10779_);
  or (_16683_, _16682_, _16672_);
  and (_16684_, _16683_, _04880_);
  or (_16685_, _16684_, _16662_);
  and (_16686_, _16685_, _10777_);
  and (_16687_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_16688_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_16689_, _16688_, _16687_);
  and (_16690_, _16689_, _04847_);
  and (_16691_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_16692_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_16693_, _16692_, _16691_);
  and (_16694_, _16693_, _10786_);
  or (_16695_, _16694_, _16690_);
  and (_16696_, _16695_, _04870_);
  and (_16697_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_16698_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_16699_, _16698_, _16697_);
  and (_16700_, _16699_, _04847_);
  and (_16701_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_16702_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_16703_, _16702_, _16701_);
  and (_16704_, _16703_, _10786_);
  or (_16705_, _16704_, _16700_);
  and (_16706_, _16705_, _10779_);
  or (_16707_, _16706_, _16696_);
  and (_16708_, _16707_, _10795_);
  or (_16709_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_16710_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_16711_, _16710_, _16709_);
  and (_16712_, _16711_, _04847_);
  or (_16713_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_16714_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_16715_, _16714_, _16713_);
  and (_16716_, _16715_, _10786_);
  or (_16717_, _16716_, _16712_);
  and (_16718_, _16717_, _04870_);
  or (_16719_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_16720_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_16721_, _16720_, _16719_);
  and (_16722_, _16721_, _04847_);
  or (_16723_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_16724_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_16725_, _16724_, _16723_);
  and (_16726_, _16725_, _10786_);
  or (_16727_, _16726_, _16722_);
  and (_16728_, _16727_, _10779_);
  or (_16729_, _16728_, _16718_);
  and (_16730_, _16729_, _04880_);
  or (_16731_, _16730_, _16708_);
  and (_16732_, _16731_, _04851_);
  or (_16733_, _16732_, _16686_);
  and (_16734_, _16733_, _04853_);
  and (_16735_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_16736_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_16737_, _16736_, _16735_);
  and (_16738_, _16737_, _04847_);
  and (_16739_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_16740_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_16741_, _16740_, _16739_);
  and (_16742_, _16741_, _10786_);
  or (_16743_, _16742_, _16738_);
  or (_16744_, _16743_, _10779_);
  and (_16745_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_16746_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_16747_, _16746_, _16745_);
  and (_16748_, _16747_, _04847_);
  and (_16749_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_16750_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_16751_, _16750_, _16749_);
  and (_16752_, _16751_, _10786_);
  or (_16753_, _16752_, _16748_);
  or (_16754_, _16753_, _04870_);
  and (_16755_, _16754_, _10795_);
  and (_16756_, _16755_, _16744_);
  or (_16757_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_16758_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_16759_, _16758_, _16757_);
  and (_16760_, _16759_, _04847_);
  or (_16761_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_16762_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_16763_, _16762_, _16761_);
  and (_16764_, _16763_, _10786_);
  or (_16765_, _16764_, _16760_);
  or (_16766_, _16765_, _10779_);
  or (_16767_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_16768_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_16769_, _16768_, _16767_);
  and (_16770_, _16769_, _04847_);
  or (_16771_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_16772_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_16773_, _16772_, _16771_);
  and (_16774_, _16773_, _10786_);
  or (_16775_, _16774_, _16770_);
  or (_16776_, _16775_, _04870_);
  and (_16777_, _16776_, _04880_);
  and (_16778_, _16777_, _16766_);
  or (_16779_, _16778_, _16756_);
  and (_16780_, _16779_, _04851_);
  and (_16781_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_16782_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_16783_, _16782_, _16781_);
  and (_16784_, _16783_, _04847_);
  and (_16785_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_16786_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_16787_, _16786_, _16785_);
  and (_16788_, _16787_, _10786_);
  or (_16789_, _16788_, _16784_);
  or (_16790_, _16789_, _10779_);
  and (_16791_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_16792_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_16793_, _16792_, _16791_);
  and (_16794_, _16793_, _04847_);
  and (_16795_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_16796_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_16797_, _16796_, _16795_);
  and (_16798_, _16797_, _10786_);
  or (_16799_, _16798_, _16794_);
  or (_16800_, _16799_, _04870_);
  and (_16801_, _16800_, _10795_);
  and (_16802_, _16801_, _16790_);
  or (_16803_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_16804_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_16805_, _16804_, _10786_);
  and (_16806_, _16805_, _16803_);
  or (_16807_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_16808_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_16809_, _16808_, _04847_);
  and (_16810_, _16809_, _16807_);
  or (_16811_, _16810_, _16806_);
  or (_16812_, _16811_, _10779_);
  or (_16813_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_16814_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_16815_, _16814_, _10786_);
  and (_16816_, _16815_, _16813_);
  or (_16817_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_16818_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_16819_, _16818_, _04847_);
  and (_16820_, _16819_, _16817_);
  or (_16821_, _16820_, _16816_);
  or (_16822_, _16821_, _04870_);
  and (_16823_, _16822_, _04880_);
  and (_16824_, _16823_, _16812_);
  or (_16825_, _16824_, _16802_);
  and (_16826_, _16825_, _10777_);
  or (_16827_, _16826_, _16780_);
  and (_16828_, _16827_, _10849_);
  or (_16829_, _16828_, _16734_);
  or (_16830_, _16829_, _04858_);
  and (_16831_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_16832_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_16833_, _16832_, _16831_);
  and (_16834_, _16833_, _10786_);
  and (_16835_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_16836_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_16837_, _16836_, _16835_);
  and (_16838_, _16837_, _04847_);
  or (_16839_, _16838_, _16834_);
  or (_16840_, _16839_, _10779_);
  and (_16841_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_16842_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_16843_, _16842_, _16841_);
  and (_16844_, _16843_, _10786_);
  and (_16845_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_16846_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_16847_, _16846_, _16845_);
  and (_16848_, _16847_, _04847_);
  or (_16849_, _16848_, _16844_);
  or (_16850_, _16849_, _04870_);
  and (_16851_, _16850_, _10795_);
  and (_16852_, _16851_, _16840_);
  or (_16853_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_16854_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_16855_, _16854_, _04847_);
  and (_16856_, _16855_, _16853_);
  or (_16857_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_16858_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_16859_, _16858_, _10786_);
  and (_16860_, _16859_, _16857_);
  or (_16861_, _16860_, _16856_);
  or (_16862_, _16861_, _10779_);
  or (_16863_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_16864_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_16865_, _16864_, _04847_);
  and (_16866_, _16865_, _16863_);
  or (_16867_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_16868_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_16869_, _16868_, _10786_);
  and (_16870_, _16869_, _16867_);
  or (_16871_, _16870_, _16866_);
  or (_16872_, _16871_, _04870_);
  and (_16873_, _16872_, _04880_);
  and (_16874_, _16873_, _16862_);
  or (_16875_, _16874_, _16852_);
  and (_16876_, _16875_, _10777_);
  and (_16877_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_16878_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_16879_, _16878_, _04847_);
  or (_16880_, _16879_, _16877_);
  and (_16881_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_16882_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_16883_, _16882_, _10786_);
  or (_16884_, _16883_, _16881_);
  and (_16885_, _16884_, _16880_);
  or (_16886_, _16885_, _10779_);
  and (_16887_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_16888_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_16889_, _16888_, _04847_);
  or (_16890_, _16889_, _16887_);
  and (_16891_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_16892_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_16893_, _16892_, _10786_);
  or (_16894_, _16893_, _16891_);
  and (_16895_, _16894_, _16890_);
  or (_16896_, _16895_, _04870_);
  and (_16897_, _16896_, _10795_);
  and (_16898_, _16897_, _16886_);
  or (_16899_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_16900_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_16901_, _16900_, _16899_);
  or (_16902_, _16901_, _10786_);
  or (_16903_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_16904_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_16905_, _16904_, _16903_);
  or (_16906_, _16905_, _04847_);
  and (_16907_, _16906_, _16902_);
  or (_16908_, _16907_, _10779_);
  or (_16909_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_16910_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_16911_, _16910_, _16909_);
  or (_16912_, _16911_, _10786_);
  or (_16913_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_16914_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_16915_, _16914_, _16913_);
  or (_16916_, _16915_, _04847_);
  and (_16917_, _16916_, _16912_);
  or (_16918_, _16917_, _04870_);
  and (_16919_, _16918_, _04880_);
  and (_16920_, _16919_, _16908_);
  or (_16921_, _16920_, _16898_);
  and (_16922_, _16921_, _04851_);
  or (_16923_, _16922_, _16876_);
  and (_16924_, _16923_, _10849_);
  and (_16925_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_16926_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_16928_, _16926_, _16925_);
  and (_16929_, _16928_, _04847_);
  and (_16930_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_16931_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_16932_, _16931_, _16930_);
  and (_16933_, _16932_, _10786_);
  or (_16934_, _16933_, _16929_);
  and (_16935_, _16934_, _04870_);
  and (_16936_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_16937_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_16938_, _16937_, _16936_);
  and (_16939_, _16938_, _04847_);
  and (_16940_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_16941_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_16942_, _16941_, _16940_);
  and (_16943_, _16942_, _10786_);
  or (_16944_, _16943_, _16939_);
  and (_16945_, _16944_, _10779_);
  or (_16946_, _16945_, _16935_);
  and (_16947_, _16946_, _10795_);
  or (_16949_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_16950_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_16951_, _16950_, _16949_);
  and (_16952_, _16951_, _04847_);
  or (_16953_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_16954_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_16955_, _16954_, _16953_);
  and (_16956_, _16955_, _10786_);
  or (_16957_, _16956_, _16952_);
  and (_16958_, _16957_, _04870_);
  or (_16959_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_16960_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_16961_, _16960_, _16959_);
  and (_16962_, _16961_, _04847_);
  or (_16963_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_16964_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_16965_, _16964_, _16963_);
  and (_16966_, _16965_, _10786_);
  or (_16967_, _16966_, _16962_);
  and (_16968_, _16967_, _10779_);
  or (_16969_, _16968_, _16958_);
  and (_16970_, _16969_, _04880_);
  or (_16971_, _16970_, _16947_);
  and (_16972_, _16971_, _04851_);
  and (_16973_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  and (_16974_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_16975_, _16974_, _16973_);
  and (_16976_, _16975_, _04847_);
  and (_16977_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  and (_16978_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_16979_, _16978_, _16977_);
  and (_16980_, _16979_, _10786_);
  or (_16981_, _16980_, _16976_);
  and (_16982_, _16981_, _04870_);
  and (_16983_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  and (_16984_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_16985_, _16984_, _16983_);
  and (_16986_, _16985_, _04847_);
  and (_16987_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  and (_16988_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_16989_, _16988_, _16987_);
  and (_16990_, _16989_, _10786_);
  or (_16991_, _16990_, _16986_);
  and (_16992_, _16991_, _10779_);
  or (_16993_, _16992_, _16982_);
  and (_16994_, _16993_, _10795_);
  or (_16995_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_16996_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  and (_16997_, _16996_, _16995_);
  and (_16998_, _16997_, _04847_);
  or (_16999_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_17000_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  and (_17001_, _17000_, _16999_);
  and (_17002_, _17001_, _10786_);
  or (_17003_, _17002_, _16998_);
  and (_17004_, _17003_, _04870_);
  or (_17005_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_17006_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and (_17007_, _17006_, _17005_);
  and (_17008_, _17007_, _04847_);
  or (_17009_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_17010_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  and (_17011_, _17010_, _17009_);
  and (_17012_, _17011_, _10786_);
  or (_17013_, _17012_, _17008_);
  and (_17014_, _17013_, _10779_);
  or (_17015_, _17014_, _17004_);
  and (_17016_, _17015_, _04880_);
  or (_17017_, _17016_, _16994_);
  and (_17018_, _17017_, _10777_);
  or (_17019_, _17018_, _16972_);
  and (_17020_, _17019_, _04853_);
  or (_17021_, _17020_, _16924_);
  or (_17022_, _17021_, _11038_);
  and (_17023_, _17022_, _16830_);
  or (_17024_, _17023_, _03372_);
  and (_17025_, _17024_, _16639_);
  or (_17026_, _17025_, _04902_);
  or (_17027_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_17028_, _17027_, _23049_);
  and (_08768_, _17028_, _17026_);
  and (_17029_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_17030_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_17031_, _17030_, _17029_);
  and (_17032_, _17031_, _04847_);
  and (_17033_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_17034_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_17035_, _17034_, _17033_);
  and (_17036_, _17035_, _10786_);
  or (_17037_, _17036_, _17032_);
  or (_17038_, _17037_, _10779_);
  and (_17039_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_17040_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_17041_, _17040_, _17039_);
  and (_17042_, _17041_, _04847_);
  and (_17043_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_17044_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_17045_, _17044_, _17043_);
  and (_17046_, _17045_, _10786_);
  or (_17047_, _17046_, _17042_);
  or (_17048_, _17047_, _04870_);
  and (_17049_, _17048_, _10795_);
  and (_17050_, _17049_, _17038_);
  or (_17051_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_17052_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_17053_, _17052_, _17051_);
  and (_17054_, _17053_, _04847_);
  or (_17055_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_17056_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_17057_, _17056_, _17055_);
  and (_17058_, _17057_, _10786_);
  or (_17059_, _17058_, _17054_);
  or (_17060_, _17059_, _10779_);
  or (_17061_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_17062_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_17063_, _17062_, _17061_);
  and (_17064_, _17063_, _04847_);
  or (_17065_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_17066_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_17067_, _17066_, _17065_);
  and (_17069_, _17067_, _10786_);
  or (_17070_, _17069_, _17064_);
  or (_17071_, _17070_, _04870_);
  and (_17072_, _17071_, _04880_);
  and (_17073_, _17072_, _17060_);
  or (_17074_, _17073_, _17050_);
  and (_17075_, _17074_, _04851_);
  and (_17076_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_17077_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_17078_, _17077_, _17076_);
  and (_17079_, _17078_, _04847_);
  and (_17080_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_17081_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_17082_, _17081_, _17080_);
  and (_17083_, _17082_, _10786_);
  or (_17084_, _17083_, _17079_);
  or (_17085_, _17084_, _10779_);
  and (_17086_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_17087_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_17088_, _17087_, _17086_);
  and (_17090_, _17088_, _04847_);
  and (_17091_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_17092_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_17093_, _17092_, _17091_);
  and (_17094_, _17093_, _10786_);
  or (_17095_, _17094_, _17090_);
  or (_17096_, _17095_, _04870_);
  and (_17097_, _17096_, _10795_);
  and (_17098_, _17097_, _17085_);
  or (_17099_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_17100_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_17101_, _17100_, _10786_);
  and (_17102_, _17101_, _17099_);
  or (_17103_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_17104_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_17105_, _17104_, _04847_);
  and (_17106_, _17105_, _17103_);
  or (_17107_, _17106_, _17102_);
  or (_17108_, _17107_, _10779_);
  or (_17109_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_17110_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_17111_, _17110_, _10786_);
  and (_17112_, _17111_, _17109_);
  or (_17113_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_17114_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_17115_, _17114_, _04847_);
  and (_17116_, _17115_, _17113_);
  or (_17117_, _17116_, _17112_);
  or (_17118_, _17117_, _04870_);
  and (_17119_, _17118_, _04880_);
  and (_17120_, _17119_, _17108_);
  or (_17121_, _17120_, _17098_);
  and (_17122_, _17121_, _10777_);
  or (_17123_, _17122_, _17075_);
  and (_17124_, _17123_, _10849_);
  and (_17125_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_17126_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_17127_, _17126_, _17125_);
  and (_17128_, _17127_, _04847_);
  and (_17129_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_17130_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_17131_, _17130_, _17129_);
  and (_17132_, _17131_, _10786_);
  or (_17133_, _17132_, _17128_);
  and (_17134_, _17133_, _04870_);
  and (_17135_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_17136_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_17137_, _17136_, _17135_);
  and (_17138_, _17137_, _04847_);
  and (_17139_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_17140_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_17141_, _17140_, _17139_);
  and (_17142_, _17141_, _10786_);
  or (_17143_, _17142_, _17138_);
  and (_17144_, _17143_, _10779_);
  or (_17145_, _17144_, _17134_);
  and (_17146_, _17145_, _10795_);
  or (_17147_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_17148_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_17149_, _17148_, _10786_);
  and (_17150_, _17149_, _17147_);
  or (_17151_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_17152_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_17153_, _17152_, _04847_);
  and (_17154_, _17153_, _17151_);
  or (_17155_, _17154_, _17150_);
  and (_17156_, _17155_, _04870_);
  or (_17157_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_17158_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_17159_, _17158_, _10786_);
  and (_17160_, _17159_, _17157_);
  or (_17161_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_17162_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_17163_, _17162_, _04847_);
  and (_17164_, _17163_, _17161_);
  or (_17165_, _17164_, _17160_);
  and (_17166_, _17165_, _10779_);
  or (_17167_, _17166_, _17156_);
  and (_17168_, _17167_, _04880_);
  or (_17169_, _17168_, _17146_);
  and (_17170_, _17169_, _10777_);
  and (_17171_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_17172_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_17173_, _17172_, _17171_);
  and (_17174_, _17173_, _04847_);
  and (_17175_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_17176_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_17177_, _17176_, _17175_);
  and (_17178_, _17177_, _10786_);
  or (_17179_, _17178_, _17174_);
  and (_17180_, _17179_, _04870_);
  and (_17181_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_17182_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_17183_, _17182_, _17181_);
  and (_17184_, _17183_, _04847_);
  and (_17185_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_17186_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_17187_, _17186_, _17185_);
  and (_17188_, _17187_, _10786_);
  or (_17189_, _17188_, _17184_);
  and (_17190_, _17189_, _10779_);
  or (_17191_, _17190_, _17180_);
  and (_17192_, _17191_, _10795_);
  or (_17193_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_17194_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_17195_, _17194_, _17193_);
  and (_17196_, _17195_, _04847_);
  or (_17197_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_17198_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_17199_, _17198_, _17197_);
  and (_17200_, _17199_, _10786_);
  or (_17201_, _17200_, _17196_);
  and (_17202_, _17201_, _04870_);
  or (_17203_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_17204_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_17205_, _17204_, _17203_);
  and (_17206_, _17205_, _04847_);
  or (_17207_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_17208_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_17209_, _17208_, _17207_);
  and (_17210_, _17209_, _10786_);
  or (_17211_, _17210_, _17206_);
  and (_17212_, _17211_, _10779_);
  or (_17213_, _17212_, _17202_);
  and (_17214_, _17213_, _04880_);
  or (_17215_, _17214_, _17192_);
  and (_17216_, _17215_, _04851_);
  or (_17217_, _17216_, _17170_);
  and (_17218_, _17217_, _04853_);
  or (_17219_, _17218_, _17124_);
  or (_17220_, _17219_, _04858_);
  and (_17221_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_17222_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_17223_, _17222_, _17221_);
  and (_17224_, _17223_, _04847_);
  and (_17225_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_17226_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_17227_, _17226_, _17225_);
  and (_17228_, _17227_, _10786_);
  or (_17229_, _17228_, _17224_);
  or (_17230_, _17229_, _10779_);
  and (_17231_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_17232_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_17233_, _17232_, _17231_);
  and (_17234_, _17233_, _04847_);
  and (_17235_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_17236_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_17237_, _17236_, _17235_);
  and (_17238_, _17237_, _10786_);
  or (_17239_, _17238_, _17234_);
  or (_17240_, _17239_, _04870_);
  and (_17241_, _17240_, _10795_);
  and (_17242_, _17241_, _17230_);
  or (_17243_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_17244_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_17245_, _17244_, _10786_);
  and (_17246_, _17245_, _17243_);
  or (_17247_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_17248_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_17249_, _17248_, _04847_);
  and (_17250_, _17249_, _17247_);
  or (_17251_, _17250_, _17246_);
  or (_17252_, _17251_, _10779_);
  or (_17253_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_17254_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_17255_, _17254_, _10786_);
  and (_17256_, _17255_, _17253_);
  or (_17257_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_17258_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_17259_, _17258_, _04847_);
  and (_17260_, _17259_, _17257_);
  or (_17261_, _17260_, _17256_);
  or (_17262_, _17261_, _04870_);
  and (_17263_, _17262_, _04880_);
  and (_17264_, _17263_, _17252_);
  or (_17265_, _17264_, _17242_);
  and (_17266_, _17265_, _10777_);
  and (_17267_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_17268_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_17269_, _17268_, _17267_);
  and (_17270_, _17269_, _04847_);
  and (_17271_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_17272_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_17273_, _17272_, _17271_);
  and (_17274_, _17273_, _10786_);
  or (_17275_, _17274_, _17270_);
  or (_17276_, _17275_, _10779_);
  and (_17277_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_17278_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_17279_, _17278_, _17277_);
  and (_17280_, _17279_, _04847_);
  and (_17281_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_17282_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_17283_, _17282_, _17281_);
  and (_17284_, _17283_, _10786_);
  or (_17285_, _17284_, _17280_);
  or (_17286_, _17285_, _04870_);
  and (_17287_, _17286_, _10795_);
  and (_17288_, _17287_, _17276_);
  or (_17289_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_17290_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_17291_, _17290_, _17289_);
  and (_17292_, _17291_, _04847_);
  or (_17293_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_17294_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_17295_, _17294_, _17293_);
  and (_17296_, _17295_, _10786_);
  or (_17297_, _17296_, _17292_);
  or (_17298_, _17297_, _10779_);
  or (_17299_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_17300_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_17301_, _17300_, _17299_);
  and (_17302_, _17301_, _04847_);
  or (_17303_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_17304_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_17305_, _17304_, _17303_);
  and (_17306_, _17305_, _10786_);
  or (_17307_, _17306_, _17302_);
  or (_17308_, _17307_, _04870_);
  and (_17309_, _17308_, _04880_);
  and (_17310_, _17309_, _17298_);
  or (_17311_, _17310_, _17288_);
  and (_17312_, _17311_, _04851_);
  or (_17313_, _17312_, _17266_);
  and (_17314_, _17313_, _10849_);
  or (_17315_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_17316_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_17317_, _17316_, _17315_);
  and (_17318_, _17317_, _04847_);
  or (_17319_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_17320_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_17321_, _17320_, _17319_);
  and (_17322_, _17321_, _10786_);
  or (_17323_, _17322_, _17318_);
  and (_17324_, _17323_, _10779_);
  or (_17325_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_17326_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_17327_, _17326_, _17325_);
  and (_17328_, _17327_, _04847_);
  or (_17329_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_17330_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_17331_, _17330_, _17329_);
  and (_17332_, _17331_, _10786_);
  or (_17333_, _17332_, _17328_);
  and (_17334_, _17333_, _04870_);
  or (_17335_, _17334_, _17324_);
  and (_17336_, _17335_, _04880_);
  and (_17337_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_17338_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_17339_, _17338_, _17337_);
  and (_17340_, _17339_, _04847_);
  and (_17341_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_17342_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_17343_, _17342_, _17341_);
  and (_17344_, _17343_, _10786_);
  or (_17345_, _17344_, _17340_);
  and (_17346_, _17345_, _10779_);
  and (_17347_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_17348_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_17349_, _17348_, _17347_);
  and (_17350_, _17349_, _04847_);
  and (_17351_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_17352_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_17353_, _17352_, _17351_);
  and (_17354_, _17353_, _10786_);
  or (_17355_, _17354_, _17350_);
  and (_17356_, _17355_, _04870_);
  or (_17357_, _17356_, _17346_);
  and (_17358_, _17357_, _10795_);
  or (_17359_, _17358_, _17336_);
  and (_17360_, _17359_, _04851_);
  or (_17361_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_17362_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_17363_, _17362_, _10786_);
  and (_17364_, _17363_, _17361_);
  or (_17365_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_17366_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_17367_, _17366_, _04847_);
  and (_17368_, _17367_, _17365_);
  or (_17369_, _17368_, _17364_);
  and (_17370_, _17369_, _10779_);
  or (_17371_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_17372_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_17373_, _17372_, _10786_);
  and (_17374_, _17373_, _17371_);
  or (_17375_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_17376_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_17377_, _17376_, _04847_);
  and (_17378_, _17377_, _17375_);
  or (_17379_, _17378_, _17374_);
  and (_17380_, _17379_, _04870_);
  or (_17381_, _17380_, _17370_);
  and (_17382_, _17381_, _04880_);
  and (_17383_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_17384_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_17385_, _17384_, _17383_);
  and (_17386_, _17385_, _04847_);
  and (_17387_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_17388_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_17389_, _17388_, _17387_);
  and (_17390_, _17389_, _10786_);
  or (_17391_, _17390_, _17386_);
  and (_17392_, _17391_, _10779_);
  and (_17393_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_17394_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_17395_, _17394_, _17393_);
  and (_17396_, _17395_, _04847_);
  and (_17397_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_17398_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_17399_, _17398_, _17397_);
  and (_17401_, _17399_, _10786_);
  or (_17402_, _17401_, _17396_);
  and (_17403_, _17402_, _04870_);
  or (_17404_, _17403_, _17392_);
  and (_17405_, _17404_, _10795_);
  or (_17406_, _17405_, _17382_);
  and (_17407_, _17406_, _10777_);
  or (_17408_, _17407_, _17360_);
  and (_17409_, _17408_, _04853_);
  or (_17410_, _17409_, _17314_);
  or (_17411_, _17410_, _11038_);
  and (_17412_, _17411_, _17220_);
  or (_17413_, _17412_, _25445_);
  and (_17414_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_17415_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_17416_, _17415_, _17414_);
  and (_17417_, _17416_, _04847_);
  and (_17418_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_17419_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_17420_, _17419_, _17418_);
  and (_17421_, _17420_, _10786_);
  or (_17422_, _17421_, _17417_);
  or (_17423_, _17422_, _10779_);
  and (_17424_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_17425_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_17426_, _17425_, _17424_);
  and (_17427_, _17426_, _04847_);
  and (_17428_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_17429_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_17430_, _17429_, _17428_);
  and (_17432_, _17430_, _10786_);
  or (_17433_, _17432_, _17427_);
  or (_17434_, _17433_, _04870_);
  and (_17435_, _17434_, _10795_);
  and (_17436_, _17435_, _17423_);
  or (_17437_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_17438_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_17439_, _17438_, _17437_);
  and (_17440_, _17439_, _04847_);
  or (_17441_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_17442_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_17443_, _17442_, _17441_);
  and (_17444_, _17443_, _10786_);
  or (_17445_, _17444_, _17440_);
  or (_17446_, _17445_, _10779_);
  or (_17447_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_17448_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_17449_, _17448_, _17447_);
  and (_17450_, _17449_, _04847_);
  or (_17451_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_17453_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_17454_, _17453_, _17451_);
  and (_17455_, _17454_, _10786_);
  or (_17456_, _17455_, _17450_);
  or (_17457_, _17456_, _04870_);
  and (_17458_, _17457_, _04880_);
  and (_17459_, _17458_, _17446_);
  or (_17460_, _17459_, _17436_);
  and (_17461_, _17460_, _04851_);
  and (_17462_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_17463_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_17464_, _17463_, _17462_);
  and (_17465_, _17464_, _04847_);
  and (_17466_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_17467_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_17468_, _17467_, _17466_);
  and (_17469_, _17468_, _10786_);
  or (_17470_, _17469_, _17465_);
  or (_17471_, _17470_, _10779_);
  and (_17472_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_17473_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_17474_, _17473_, _17472_);
  and (_17475_, _17474_, _04847_);
  and (_17476_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_17477_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_17478_, _17477_, _17476_);
  and (_17479_, _17478_, _10786_);
  or (_17480_, _17479_, _17475_);
  or (_17481_, _17480_, _04870_);
  and (_17482_, _17481_, _10795_);
  and (_17483_, _17482_, _17471_);
  or (_17484_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_17485_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_17486_, _17485_, _10786_);
  and (_17487_, _17486_, _17484_);
  or (_17488_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_17489_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_17490_, _17489_, _04847_);
  and (_17491_, _17490_, _17488_);
  or (_17492_, _17491_, _17487_);
  or (_17493_, _17492_, _10779_);
  or (_17494_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_17495_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_17496_, _17495_, _10786_);
  and (_17497_, _17496_, _17494_);
  or (_17498_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_17499_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_17500_, _17499_, _04847_);
  and (_17501_, _17500_, _17498_);
  or (_17502_, _17501_, _17497_);
  or (_17503_, _17502_, _04870_);
  and (_17504_, _17503_, _04880_);
  and (_17505_, _17504_, _17493_);
  or (_17506_, _17505_, _17483_);
  and (_17507_, _17506_, _10777_);
  or (_17508_, _17507_, _17461_);
  and (_17509_, _17508_, _10849_);
  and (_17510_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_17511_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_17512_, _17511_, _17510_);
  and (_17513_, _17512_, _04847_);
  and (_17514_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_17515_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_17516_, _17515_, _17514_);
  and (_17517_, _17516_, _10786_);
  or (_17518_, _17517_, _17513_);
  and (_17519_, _17518_, _04870_);
  and (_17520_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_17521_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_17522_, _17521_, _17520_);
  and (_17523_, _17522_, _04847_);
  and (_17524_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_17525_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_17526_, _17525_, _17524_);
  and (_17527_, _17526_, _10786_);
  or (_17528_, _17527_, _17523_);
  and (_17529_, _17528_, _10779_);
  or (_17530_, _17529_, _17519_);
  and (_17531_, _17530_, _10795_);
  or (_17532_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_17533_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_17534_, _17533_, _10786_);
  and (_17535_, _17534_, _17532_);
  or (_17536_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_17537_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_17538_, _17537_, _04847_);
  and (_17539_, _17538_, _17536_);
  or (_17540_, _17539_, _17535_);
  and (_17541_, _17540_, _04870_);
  or (_17542_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_17543_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_17544_, _17543_, _10786_);
  and (_17545_, _17544_, _17542_);
  or (_17546_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_17547_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_17548_, _17547_, _04847_);
  and (_17549_, _17548_, _17546_);
  or (_17550_, _17549_, _17545_);
  and (_17551_, _17550_, _10779_);
  or (_17552_, _17551_, _17541_);
  and (_17553_, _17552_, _04880_);
  or (_17554_, _17553_, _17531_);
  and (_17555_, _17554_, _10777_);
  and (_17556_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_17557_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_17558_, _17557_, _17556_);
  and (_17559_, _17558_, _04847_);
  and (_17560_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_17561_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_17562_, _17561_, _17560_);
  and (_17563_, _17562_, _10786_);
  or (_17564_, _17563_, _17559_);
  and (_17565_, _17564_, _04870_);
  and (_17566_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_17567_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_17568_, _17567_, _17566_);
  and (_17569_, _17568_, _04847_);
  and (_17570_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_17571_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_17572_, _17571_, _17570_);
  and (_17573_, _17572_, _10786_);
  or (_17574_, _17573_, _17569_);
  and (_17575_, _17574_, _10779_);
  or (_17576_, _17575_, _17565_);
  and (_17577_, _17576_, _10795_);
  or (_17578_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_17579_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_17580_, _17579_, _17578_);
  and (_17581_, _17580_, _04847_);
  or (_17582_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_17583_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_17584_, _17583_, _17582_);
  and (_17585_, _17584_, _10786_);
  or (_17586_, _17585_, _17581_);
  and (_17587_, _17586_, _04870_);
  or (_17588_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_17589_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_17590_, _17589_, _17588_);
  and (_17591_, _17590_, _04847_);
  or (_17592_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_17593_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_17594_, _17593_, _17592_);
  and (_17595_, _17594_, _10786_);
  or (_17596_, _17595_, _17591_);
  and (_17597_, _17596_, _10779_);
  or (_17598_, _17597_, _17587_);
  and (_17599_, _17598_, _04880_);
  or (_17600_, _17599_, _17577_);
  and (_17601_, _17600_, _04851_);
  or (_17602_, _17601_, _17555_);
  and (_17603_, _17602_, _04853_);
  or (_17604_, _17603_, _17509_);
  or (_17605_, _17604_, _04858_);
  and (_17606_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_17607_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_17608_, _17607_, _17606_);
  and (_17609_, _17608_, _04847_);
  and (_17610_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_17611_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_17612_, _17611_, _17610_);
  and (_17613_, _17612_, _10786_);
  or (_17614_, _17613_, _17609_);
  or (_17615_, _17614_, _10779_);
  and (_17616_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_17617_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_17618_, _17617_, _17616_);
  and (_17619_, _17618_, _04847_);
  and (_17620_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_17621_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_17622_, _17621_, _17620_);
  and (_17623_, _17622_, _10786_);
  or (_17624_, _17623_, _17619_);
  or (_17625_, _17624_, _04870_);
  and (_17626_, _17625_, _10795_);
  and (_17627_, _17626_, _17615_);
  or (_17628_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_17629_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_17630_, _17629_, _10786_);
  and (_17631_, _17630_, _17628_);
  or (_17632_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_17633_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_17634_, _17633_, _04847_);
  and (_17635_, _17634_, _17632_);
  or (_17636_, _17635_, _17631_);
  or (_17637_, _17636_, _10779_);
  or (_17638_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_17639_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_17640_, _17639_, _10786_);
  and (_17641_, _17640_, _17638_);
  or (_17642_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_17643_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_17644_, _17643_, _04847_);
  and (_17645_, _17644_, _17642_);
  or (_17646_, _17645_, _17641_);
  or (_17647_, _17646_, _04870_);
  and (_17648_, _17647_, _04880_);
  and (_17649_, _17648_, _17637_);
  or (_17650_, _17649_, _17627_);
  and (_17651_, _17650_, _10777_);
  and (_17652_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_17653_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_17654_, _17653_, _17652_);
  and (_17655_, _17654_, _04847_);
  and (_17656_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_17657_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_17658_, _17657_, _17656_);
  and (_17659_, _17658_, _10786_);
  or (_17660_, _17659_, _17655_);
  or (_17661_, _17660_, _10779_);
  and (_17662_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_17663_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_17664_, _17663_, _17662_);
  and (_17665_, _17664_, _04847_);
  and (_17666_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_17667_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_17668_, _17667_, _17666_);
  and (_17669_, _17668_, _10786_);
  or (_17670_, _17669_, _17665_);
  or (_17671_, _17670_, _04870_);
  and (_17672_, _17671_, _10795_);
  and (_17673_, _17672_, _17661_);
  or (_17674_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_17675_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_17676_, _17675_, _17674_);
  and (_17677_, _17676_, _04847_);
  or (_17678_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_17679_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_17680_, _17679_, _17678_);
  and (_17681_, _17680_, _10786_);
  or (_17682_, _17681_, _17677_);
  or (_17683_, _17682_, _10779_);
  or (_17684_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_17685_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_17686_, _17685_, _17684_);
  and (_17687_, _17686_, _04847_);
  or (_17688_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_17689_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_17690_, _17689_, _17688_);
  and (_17691_, _17690_, _10786_);
  or (_17692_, _17691_, _17687_);
  or (_17693_, _17692_, _04870_);
  and (_17694_, _17693_, _04880_);
  and (_17695_, _17694_, _17683_);
  or (_17696_, _17695_, _17673_);
  and (_17697_, _17696_, _04851_);
  or (_17698_, _17697_, _17651_);
  and (_17699_, _17698_, _10849_);
  or (_17700_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_17701_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_17702_, _17701_, _17700_);
  and (_17703_, _17702_, _04847_);
  or (_17704_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_17705_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_17706_, _17705_, _17704_);
  and (_17707_, _17706_, _10786_);
  or (_17708_, _17707_, _17703_);
  and (_17709_, _17708_, _10779_);
  or (_17710_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_17711_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_17712_, _17711_, _17710_);
  and (_17713_, _17712_, _04847_);
  or (_17714_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_17715_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_17716_, _17715_, _17714_);
  and (_17717_, _17716_, _10786_);
  or (_17718_, _17717_, _17713_);
  and (_17719_, _17718_, _04870_);
  or (_17720_, _17719_, _17709_);
  and (_17721_, _17720_, _04880_);
  and (_17722_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_17723_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_17724_, _17723_, _17722_);
  and (_17725_, _17724_, _04847_);
  and (_17726_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_17727_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_17728_, _17727_, _17726_);
  and (_17729_, _17728_, _10786_);
  or (_17730_, _17729_, _17725_);
  and (_17731_, _17730_, _10779_);
  and (_17732_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_17733_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_17734_, _17733_, _17732_);
  and (_17735_, _17734_, _04847_);
  and (_17736_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_17737_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_17738_, _17737_, _17736_);
  and (_17739_, _17738_, _10786_);
  or (_17740_, _17739_, _17735_);
  and (_17741_, _17740_, _04870_);
  or (_17742_, _17741_, _17731_);
  and (_17743_, _17742_, _10795_);
  or (_17744_, _17743_, _17721_);
  and (_17745_, _17744_, _04851_);
  or (_17746_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_17747_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_17748_, _17747_, _10786_);
  and (_17749_, _17748_, _17746_);
  or (_17750_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_17751_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_17752_, _17751_, _04847_);
  and (_17753_, _17752_, _17750_);
  or (_17754_, _17753_, _17749_);
  and (_17755_, _17754_, _10779_);
  or (_17756_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_17757_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_17758_, _17757_, _10786_);
  and (_17759_, _17758_, _17756_);
  or (_17760_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_17761_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_17762_, _17761_, _04847_);
  and (_17763_, _17762_, _17760_);
  or (_17764_, _17763_, _17759_);
  and (_17765_, _17764_, _04870_);
  or (_17766_, _17765_, _17755_);
  and (_17767_, _17766_, _04880_);
  and (_17768_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_17769_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_17770_, _17769_, _17768_);
  and (_17771_, _17770_, _04847_);
  and (_17772_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_17773_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_17774_, _17773_, _17772_);
  and (_17775_, _17774_, _10786_);
  or (_17776_, _17775_, _17771_);
  and (_17777_, _17776_, _10779_);
  and (_17778_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_17779_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_17780_, _17779_, _17778_);
  and (_17781_, _17780_, _04847_);
  and (_17782_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_17783_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_17784_, _17783_, _17782_);
  and (_17785_, _17784_, _10786_);
  or (_17786_, _17785_, _17781_);
  and (_17787_, _17786_, _04870_);
  or (_17788_, _17787_, _17777_);
  and (_17789_, _17788_, _10795_);
  or (_17790_, _17789_, _17767_);
  and (_17791_, _17790_, _10777_);
  or (_17792_, _17791_, _17745_);
  and (_17793_, _17792_, _04853_);
  or (_17794_, _17793_, _17699_);
  or (_17795_, _17794_, _11038_);
  and (_17796_, _17795_, _17605_);
  or (_17797_, _17796_, _03372_);
  and (_17798_, _17797_, _17413_);
  or (_17799_, _17798_, _04902_);
  or (_17800_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_17801_, _17800_, _23049_);
  and (_08770_, _17801_, _17799_);
  and (_17802_, _10404_, _26242_);
  and (_17803_, _10406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_27257_, _17803_, _17802_);
  and (_17804_, _25939_, _25886_);
  and (_17805_, _25941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_08777_, _17805_, _17804_);
  and (_17806_, _01371_, _25886_);
  and (_17807_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_08781_, _17807_, _17806_);
  and (_17808_, _26242_, _26151_);
  and (_17809_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_08785_, _17809_, _17808_);
  and (_17810_, _03115_, _26085_);
  and (_17811_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_08789_, _17811_, _17810_);
  and (_17812_, _26329_, _26242_);
  and (_17813_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_08791_, _17813_, _17812_);
  and (_17814_, _14384_, _23768_);
  and (_17815_, _14386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or (_08797_, _17815_, _17814_);
  and (_17816_, _14629_, _25927_);
  and (_17817_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_08821_, _17817_, _17816_);
  and (_17818_, _04821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_17819_, _04820_, _26085_);
  or (_08825_, _17819_, _17818_);
  and (_17820_, _25927_, _23849_);
  and (_17821_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_08844_, _17821_, _17820_);
  and (_17822_, _25914_, _23848_);
  and (_17823_, _17822_, _26170_);
  not (_17824_, _17822_);
  and (_17825_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or (_08853_, _17825_, _17823_);
  and (_17826_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  and (_17827_, _10283_, _25927_);
  or (_27095_, _17827_, _17826_);
  and (_17828_, _00016_, _26085_);
  and (_17829_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_08865_, _17829_, _17828_);
  and (_17830_, _26375_, _23775_);
  and (_17831_, _17830_, _25927_);
  not (_17832_, _17830_);
  and (_17833_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_27303_, _17833_, _17831_);
  and (_17834_, _26375_, _26213_);
  and (_17835_, _17834_, _26085_);
  not (_17836_, _17834_);
  and (_17837_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_27302_, _17837_, _17835_);
  and (_17838_, _17834_, _26170_);
  and (_17839_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_08881_, _17839_, _17838_);
  and (_17840_, _26375_, _26190_);
  and (_17841_, _17840_, _26085_);
  not (_17842_, _17840_);
  and (_17843_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_08886_, _17843_, _17841_);
  and (_17844_, _17840_, _25886_);
  and (_17845_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_08889_, _17845_, _17844_);
  and (_17846_, _26375_, _25914_);
  and (_17847_, _17846_, _26185_);
  not (_17848_, _17846_);
  and (_17849_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_08893_, _17849_, _17847_);
  and (_17850_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_17851_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_17852_, _17851_, _17850_);
  and (_17853_, _17852_, _10786_);
  and (_17854_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_17855_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_17856_, _17855_, _17854_);
  and (_17857_, _17856_, _04847_);
  or (_17858_, _17857_, _17853_);
  or (_17859_, _17858_, _10779_);
  and (_17860_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_17861_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_17862_, _17861_, _17860_);
  and (_17863_, _17862_, _10786_);
  and (_17864_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_17865_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_17866_, _17865_, _17864_);
  and (_17867_, _17866_, _04847_);
  or (_17868_, _17867_, _17863_);
  or (_17869_, _17868_, _04870_);
  and (_17870_, _17869_, _10795_);
  and (_17871_, _17870_, _17859_);
  or (_17872_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_17873_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_17874_, _17873_, _04847_);
  and (_17875_, _17874_, _17872_);
  or (_17876_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_17877_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_17878_, _17877_, _10786_);
  and (_17879_, _17878_, _17876_);
  or (_17880_, _17879_, _17875_);
  or (_17881_, _17880_, _10779_);
  or (_17882_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_17883_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_17884_, _17883_, _04847_);
  and (_17885_, _17884_, _17882_);
  or (_17886_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_17887_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_17888_, _17887_, _10786_);
  and (_17889_, _17888_, _17886_);
  or (_17890_, _17889_, _17885_);
  or (_17891_, _17890_, _04870_);
  and (_17892_, _17891_, _04880_);
  and (_17893_, _17892_, _17881_);
  or (_17894_, _17893_, _17871_);
  or (_17895_, _17894_, _04851_);
  and (_17896_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_17897_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_17898_, _17897_, _04847_);
  or (_17899_, _17898_, _17896_);
  and (_17900_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_17901_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_17902_, _17901_, _10786_);
  or (_17903_, _17902_, _17900_);
  and (_17904_, _17903_, _17899_);
  or (_17905_, _17904_, _10779_);
  and (_17906_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_17907_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_17908_, _17907_, _04847_);
  or (_17909_, _17908_, _17906_);
  and (_17910_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_17911_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_17912_, _17911_, _10786_);
  or (_17913_, _17912_, _17910_);
  and (_17914_, _17913_, _17909_);
  or (_17915_, _17914_, _04870_);
  and (_17916_, _17915_, _10795_);
  and (_17917_, _17916_, _17905_);
  or (_17918_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_17919_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_17920_, _17919_, _17918_);
  or (_17921_, _17920_, _10786_);
  or (_17922_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_17923_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_17924_, _17923_, _17922_);
  or (_17925_, _17924_, _04847_);
  and (_17926_, _17925_, _17921_);
  or (_17927_, _17926_, _10779_);
  or (_17928_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_17929_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_17930_, _17929_, _17928_);
  or (_17931_, _17930_, _10786_);
  or (_17932_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_17933_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_17934_, _17933_, _17932_);
  or (_17935_, _17934_, _04847_);
  and (_17936_, _17935_, _17931_);
  or (_17937_, _17936_, _04870_);
  and (_17938_, _17937_, _04880_);
  and (_17939_, _17938_, _17927_);
  or (_17940_, _17939_, _17917_);
  or (_17941_, _17940_, _10777_);
  and (_17942_, _17941_, _10849_);
  and (_17943_, _17942_, _17895_);
  and (_17944_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_17945_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_17946_, _17945_, _17944_);
  and (_17947_, _17946_, _04847_);
  and (_17948_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_17949_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_17950_, _17949_, _17948_);
  and (_17951_, _17950_, _10786_);
  or (_17952_, _17951_, _17947_);
  and (_17953_, _17952_, _04870_);
  and (_17954_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_17955_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_17956_, _17955_, _17954_);
  and (_17957_, _17956_, _04847_);
  and (_17958_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_17959_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_17960_, _17959_, _17958_);
  and (_17961_, _17960_, _10786_);
  or (_17962_, _17961_, _17957_);
  and (_17963_, _17962_, _10779_);
  or (_17964_, _17963_, _17953_);
  and (_17965_, _17964_, _10795_);
  or (_17966_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_17967_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_17968_, _17967_, _17966_);
  and (_17969_, _17968_, _04847_);
  or (_17970_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_17971_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_17972_, _17971_, _17970_);
  and (_17973_, _17972_, _10786_);
  or (_17974_, _17973_, _17969_);
  and (_17975_, _17974_, _04870_);
  or (_17976_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_17977_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_17978_, _17977_, _17976_);
  and (_17979_, _17978_, _04847_);
  or (_17980_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_17981_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_17982_, _17981_, _17980_);
  and (_17983_, _17982_, _10786_);
  or (_17984_, _17983_, _17979_);
  and (_17985_, _17984_, _10779_);
  or (_17986_, _17985_, _17975_);
  and (_17987_, _17986_, _04880_);
  or (_17988_, _17987_, _17965_);
  and (_17989_, _17988_, _10777_);
  and (_17990_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_17991_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_17992_, _17991_, _17990_);
  and (_17993_, _17992_, _04847_);
  and (_17994_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_17995_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_17996_, _17995_, _17994_);
  and (_17997_, _17996_, _10786_);
  or (_17998_, _17997_, _17993_);
  and (_17999_, _17998_, _04870_);
  and (_18000_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_18001_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_18002_, _18001_, _18000_);
  and (_18003_, _18002_, _04847_);
  and (_18004_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_18005_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_18006_, _18005_, _18004_);
  and (_18007_, _18006_, _10786_);
  or (_18008_, _18007_, _18003_);
  and (_18009_, _18008_, _10779_);
  or (_18010_, _18009_, _17999_);
  and (_18011_, _18010_, _10795_);
  or (_18012_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_18013_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_18014_, _18013_, _18012_);
  and (_18015_, _18014_, _04847_);
  or (_18016_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_18017_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_18018_, _18017_, _18016_);
  and (_18019_, _18018_, _10786_);
  or (_18020_, _18019_, _18015_);
  and (_18021_, _18020_, _04870_);
  or (_18022_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_18023_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_18024_, _18023_, _18022_);
  and (_18025_, _18024_, _04847_);
  or (_18026_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_18027_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_18028_, _18027_, _18026_);
  and (_18029_, _18028_, _10786_);
  or (_18030_, _18029_, _18025_);
  and (_18031_, _18030_, _10779_);
  or (_18032_, _18031_, _18021_);
  and (_18033_, _18032_, _04880_);
  or (_18034_, _18033_, _18011_);
  and (_18035_, _18034_, _04851_);
  or (_18036_, _18035_, _17989_);
  and (_18037_, _18036_, _04853_);
  or (_18038_, _18037_, _17943_);
  or (_18039_, _18038_, _04858_);
  and (_18040_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_18041_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_18042_, _18041_, _18040_);
  and (_18043_, _18042_, _04847_);
  and (_18044_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_18045_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_18046_, _18045_, _18044_);
  and (_18047_, _18046_, _10786_);
  or (_18048_, _18047_, _18043_);
  or (_18049_, _18048_, _10779_);
  and (_18050_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_18051_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_18052_, _18051_, _18050_);
  and (_18053_, _18052_, _04847_);
  and (_18054_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_18055_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_18056_, _18055_, _18054_);
  and (_18057_, _18056_, _10786_);
  or (_18058_, _18057_, _18053_);
  or (_18059_, _18058_, _04870_);
  and (_18060_, _18059_, _10795_);
  and (_18061_, _18060_, _18049_);
  or (_18062_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_18063_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_18064_, _18063_, _10786_);
  and (_18065_, _18064_, _18062_);
  or (_18066_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_18067_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_18068_, _18067_, _04847_);
  and (_18069_, _18068_, _18066_);
  or (_18070_, _18069_, _18065_);
  or (_18071_, _18070_, _10779_);
  or (_18072_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_18073_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_18074_, _18073_, _10786_);
  and (_18075_, _18074_, _18072_);
  or (_18076_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_18077_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_18078_, _18077_, _04847_);
  and (_18079_, _18078_, _18076_);
  or (_18080_, _18079_, _18075_);
  or (_18081_, _18080_, _04870_);
  and (_18082_, _18081_, _04880_);
  and (_18083_, _18082_, _18071_);
  or (_18084_, _18083_, _18061_);
  and (_18085_, _18084_, _10777_);
  and (_18086_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_18087_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_18088_, _18087_, _18086_);
  and (_18089_, _18088_, _04847_);
  and (_18090_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_18091_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_18092_, _18091_, _18090_);
  and (_18093_, _18092_, _10786_);
  or (_18094_, _18093_, _18089_);
  or (_18095_, _18094_, _10779_);
  and (_18096_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_18097_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_18098_, _18097_, _18096_);
  and (_18099_, _18098_, _04847_);
  and (_18100_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_18101_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_18102_, _18101_, _18100_);
  and (_18103_, _18102_, _10786_);
  or (_18104_, _18103_, _18099_);
  or (_18105_, _18104_, _04870_);
  and (_18106_, _18105_, _10795_);
  and (_18107_, _18106_, _18095_);
  or (_18108_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_18109_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_18110_, _18109_, _18108_);
  and (_18111_, _18110_, _04847_);
  or (_18112_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_18113_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_18114_, _18113_, _18112_);
  and (_18115_, _18114_, _10786_);
  or (_18116_, _18115_, _18111_);
  or (_18117_, _18116_, _10779_);
  or (_18118_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_18119_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_18120_, _18119_, _18118_);
  and (_18121_, _18120_, _04847_);
  or (_18122_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_18123_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_18124_, _18123_, _18122_);
  and (_18125_, _18124_, _10786_);
  or (_18126_, _18125_, _18121_);
  or (_18127_, _18126_, _04870_);
  and (_18128_, _18127_, _04880_);
  and (_18129_, _18128_, _18117_);
  or (_18130_, _18129_, _18107_);
  and (_18131_, _18130_, _04851_);
  or (_18132_, _18131_, _18085_);
  and (_18133_, _18132_, _10849_);
  or (_18134_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_18135_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_18136_, _18135_, _18134_);
  and (_18137_, _18136_, _04847_);
  or (_18138_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_18139_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_18140_, _18139_, _18138_);
  and (_18141_, _18140_, _10786_);
  or (_18142_, _18141_, _18137_);
  and (_18143_, _18142_, _10779_);
  or (_18144_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_18145_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_18146_, _18145_, _18144_);
  and (_18147_, _18146_, _04847_);
  or (_18148_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_18149_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_18150_, _18149_, _18148_);
  and (_18151_, _18150_, _10786_);
  or (_18152_, _18151_, _18147_);
  and (_18153_, _18152_, _04870_);
  or (_18154_, _18153_, _18143_);
  and (_18155_, _18154_, _04880_);
  and (_18156_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_18157_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_18158_, _18157_, _18156_);
  and (_18159_, _18158_, _04847_);
  and (_18160_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_18161_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_18162_, _18161_, _18160_);
  and (_18163_, _18162_, _10786_);
  or (_18164_, _18163_, _18159_);
  and (_18165_, _18164_, _10779_);
  and (_18166_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_18167_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_18168_, _18167_, _18166_);
  and (_18169_, _18168_, _04847_);
  and (_18170_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_18171_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_18172_, _18171_, _18170_);
  and (_18173_, _18172_, _10786_);
  or (_18174_, _18173_, _18169_);
  and (_18175_, _18174_, _04870_);
  or (_18176_, _18175_, _18165_);
  and (_18177_, _18176_, _10795_);
  or (_18178_, _18177_, _18155_);
  and (_18179_, _18178_, _04851_);
  or (_18180_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_18181_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_18182_, _18181_, _10786_);
  and (_18183_, _18182_, _18180_);
  or (_18184_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_18185_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_18186_, _18185_, _04847_);
  and (_18187_, _18186_, _18184_);
  or (_18188_, _18187_, _18183_);
  and (_18189_, _18188_, _10779_);
  or (_18190_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_18191_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_18192_, _18191_, _10786_);
  and (_18193_, _18192_, _18190_);
  or (_18194_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_18195_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_18196_, _18195_, _04847_);
  and (_18197_, _18196_, _18194_);
  or (_18198_, _18197_, _18193_);
  and (_18199_, _18198_, _04870_);
  or (_18200_, _18199_, _18189_);
  and (_18201_, _18200_, _04880_);
  and (_18202_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_18203_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_18204_, _18203_, _18202_);
  and (_18205_, _18204_, _04847_);
  and (_18206_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_18207_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_18208_, _18207_, _18206_);
  and (_18209_, _18208_, _10786_);
  or (_18210_, _18209_, _18205_);
  and (_18211_, _18210_, _10779_);
  and (_18212_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_18213_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_18214_, _18213_, _18212_);
  and (_18215_, _18214_, _04847_);
  and (_18216_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_18217_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_18218_, _18217_, _18216_);
  and (_18219_, _18218_, _10786_);
  or (_18220_, _18219_, _18215_);
  and (_18221_, _18220_, _04870_);
  or (_18222_, _18221_, _18211_);
  and (_18223_, _18222_, _10795_);
  or (_18224_, _18223_, _18201_);
  and (_18225_, _18224_, _10777_);
  or (_18226_, _18225_, _18179_);
  and (_18227_, _18226_, _04853_);
  or (_18228_, _18227_, _18133_);
  or (_18229_, _18228_, _11038_);
  and (_18230_, _18229_, _18039_);
  or (_18231_, _18230_, _25445_);
  and (_18232_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_18233_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_18234_, _18233_, _18232_);
  and (_18235_, _18234_, _04847_);
  and (_18236_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_18237_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_18238_, _18237_, _18236_);
  and (_18239_, _18238_, _10786_);
  or (_18240_, _18239_, _18235_);
  or (_18241_, _18240_, _10779_);
  and (_18242_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_18243_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_18244_, _18243_, _18242_);
  and (_18245_, _18244_, _04847_);
  and (_18246_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_18247_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_18248_, _18247_, _18246_);
  and (_18249_, _18248_, _10786_);
  or (_18250_, _18249_, _18245_);
  or (_18251_, _18250_, _04870_);
  and (_18252_, _18251_, _10795_);
  and (_18253_, _18252_, _18241_);
  or (_18254_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_18255_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_18256_, _18255_, _18254_);
  and (_18257_, _18256_, _04847_);
  or (_18258_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_18259_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_18260_, _18259_, _18258_);
  and (_18261_, _18260_, _10786_);
  or (_18262_, _18261_, _18257_);
  or (_18263_, _18262_, _10779_);
  or (_18264_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_18265_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_18266_, _18265_, _18264_);
  and (_18267_, _18266_, _04847_);
  or (_18268_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_18269_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_18270_, _18269_, _18268_);
  and (_18271_, _18270_, _10786_);
  or (_18272_, _18271_, _18267_);
  or (_18273_, _18272_, _04870_);
  and (_18274_, _18273_, _04880_);
  and (_18275_, _18274_, _18263_);
  or (_18276_, _18275_, _18253_);
  and (_18277_, _18276_, _04851_);
  and (_18278_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_18279_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_18280_, _18279_, _18278_);
  and (_18281_, _18280_, _04847_);
  and (_18282_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_18283_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_18284_, _18283_, _18282_);
  and (_18285_, _18284_, _10786_);
  or (_18286_, _18285_, _18281_);
  or (_18287_, _18286_, _10779_);
  and (_18288_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_18289_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_18290_, _18289_, _18288_);
  and (_18291_, _18290_, _04847_);
  and (_18292_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_18293_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_18294_, _18293_, _18292_);
  and (_18295_, _18294_, _10786_);
  or (_18296_, _18295_, _18291_);
  or (_18297_, _18296_, _04870_);
  and (_18298_, _18297_, _10795_);
  and (_18299_, _18298_, _18287_);
  or (_18300_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_18301_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_18302_, _18301_, _10786_);
  and (_18303_, _18302_, _18300_);
  or (_18304_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_18305_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_18306_, _18305_, _04847_);
  and (_18307_, _18306_, _18304_);
  or (_18308_, _18307_, _18303_);
  or (_18309_, _18308_, _10779_);
  or (_18310_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_18311_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_18312_, _18311_, _10786_);
  and (_18313_, _18312_, _18310_);
  or (_18314_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_18315_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_18316_, _18315_, _04847_);
  and (_18317_, _18316_, _18314_);
  or (_18318_, _18317_, _18313_);
  or (_18319_, _18318_, _04870_);
  and (_18320_, _18319_, _04880_);
  and (_18321_, _18320_, _18309_);
  or (_18322_, _18321_, _18299_);
  and (_18323_, _18322_, _10777_);
  or (_18324_, _18323_, _18277_);
  and (_18325_, _18324_, _10849_);
  and (_18326_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_18327_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_18328_, _18327_, _18326_);
  and (_18329_, _18328_, _04847_);
  and (_18330_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_18331_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_18332_, _18331_, _18330_);
  and (_18333_, _18332_, _10786_);
  or (_18334_, _18333_, _18329_);
  and (_18335_, _18334_, _04870_);
  and (_18336_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_18337_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_18338_, _18337_, _18336_);
  and (_18339_, _18338_, _04847_);
  and (_18340_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_18341_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_18342_, _18341_, _18340_);
  and (_18343_, _18342_, _10786_);
  or (_18344_, _18343_, _18339_);
  and (_18345_, _18344_, _10779_);
  or (_18346_, _18345_, _18335_);
  and (_18347_, _18346_, _10795_);
  or (_18348_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_18349_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_18350_, _18349_, _10786_);
  and (_18351_, _18350_, _18348_);
  or (_18352_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_18353_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_18354_, _18353_, _04847_);
  and (_18355_, _18354_, _18352_);
  or (_18356_, _18355_, _18351_);
  and (_18357_, _18356_, _04870_);
  or (_18358_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_18359_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_18360_, _18359_, _10786_);
  and (_18361_, _18360_, _18358_);
  or (_18362_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_18363_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_18364_, _18363_, _04847_);
  and (_18365_, _18364_, _18362_);
  or (_18366_, _18365_, _18361_);
  and (_18367_, _18366_, _10779_);
  or (_18368_, _18367_, _18357_);
  and (_18369_, _18368_, _04880_);
  or (_18370_, _18369_, _18347_);
  and (_18371_, _18370_, _10777_);
  and (_18372_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_18373_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_18374_, _18373_, _18372_);
  and (_18375_, _18374_, _04847_);
  and (_18376_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_18377_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_18378_, _18377_, _18376_);
  and (_18379_, _18378_, _10786_);
  or (_18380_, _18379_, _18375_);
  and (_18381_, _18380_, _04870_);
  and (_18382_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_18383_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_18384_, _18383_, _18382_);
  and (_18385_, _18384_, _04847_);
  and (_18386_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_18387_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_18388_, _18387_, _18386_);
  and (_18389_, _18388_, _10786_);
  or (_18390_, _18389_, _18385_);
  and (_18391_, _18390_, _10779_);
  or (_18392_, _18391_, _18381_);
  and (_18393_, _18392_, _10795_);
  or (_18394_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_18395_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_18396_, _18395_, _18394_);
  and (_18397_, _18396_, _04847_);
  or (_18398_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_18399_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_18400_, _18399_, _18398_);
  and (_18401_, _18400_, _10786_);
  or (_18402_, _18401_, _18397_);
  and (_18403_, _18402_, _04870_);
  or (_18404_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_18405_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_18406_, _18405_, _18404_);
  and (_18407_, _18406_, _04847_);
  or (_18408_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_18409_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_18410_, _18409_, _18408_);
  and (_18411_, _18410_, _10786_);
  or (_18412_, _18411_, _18407_);
  and (_18413_, _18412_, _10779_);
  or (_18414_, _18413_, _18403_);
  and (_18415_, _18414_, _04880_);
  or (_18416_, _18415_, _18393_);
  and (_18417_, _18416_, _04851_);
  or (_18418_, _18417_, _18371_);
  and (_18419_, _18418_, _04853_);
  or (_18420_, _18419_, _18325_);
  or (_18421_, _18420_, _04858_);
  and (_18422_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_18423_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_18424_, _18423_, _18422_);
  and (_18425_, _18424_, _04847_);
  and (_18426_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_18427_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_18428_, _18427_, _18426_);
  and (_18429_, _18428_, _10786_);
  or (_18430_, _18429_, _18425_);
  or (_18431_, _18430_, _10779_);
  and (_18432_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_18433_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_18434_, _18433_, _18432_);
  and (_18435_, _18434_, _04847_);
  and (_18436_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_18437_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_18438_, _18437_, _18436_);
  and (_18439_, _18438_, _10786_);
  or (_18440_, _18439_, _18435_);
  or (_18441_, _18440_, _04870_);
  and (_18442_, _18441_, _10795_);
  and (_18443_, _18442_, _18431_);
  or (_18444_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_18445_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_18446_, _18445_, _10786_);
  and (_18447_, _18446_, _18444_);
  or (_18448_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_18449_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_18450_, _18449_, _04847_);
  and (_18451_, _18450_, _18448_);
  or (_18452_, _18451_, _18447_);
  or (_18453_, _18452_, _10779_);
  or (_18454_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_18455_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_18456_, _18455_, _10786_);
  and (_18457_, _18456_, _18454_);
  or (_18458_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_18459_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_18460_, _18459_, _04847_);
  and (_18461_, _18460_, _18458_);
  or (_18462_, _18461_, _18457_);
  or (_18463_, _18462_, _04870_);
  and (_18464_, _18463_, _04880_);
  and (_18465_, _18464_, _18453_);
  or (_18466_, _18465_, _18443_);
  and (_18467_, _18466_, _10777_);
  and (_18468_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_18469_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_18470_, _18469_, _18468_);
  and (_18471_, _18470_, _04847_);
  and (_18472_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_18473_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_18474_, _18473_, _18472_);
  and (_18475_, _18474_, _10786_);
  or (_18476_, _18475_, _18471_);
  or (_18477_, _18476_, _10779_);
  and (_18478_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_18479_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_18480_, _18479_, _18478_);
  and (_18481_, _18480_, _04847_);
  and (_18482_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_18483_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_18484_, _18483_, _18482_);
  and (_18485_, _18484_, _10786_);
  or (_18486_, _18485_, _18481_);
  or (_18487_, _18486_, _04870_);
  and (_18488_, _18487_, _10795_);
  and (_18489_, _18488_, _18477_);
  or (_18490_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_18491_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_18492_, _18491_, _18490_);
  and (_18493_, _18492_, _04847_);
  or (_18494_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_18495_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_18496_, _18495_, _18494_);
  and (_18497_, _18496_, _10786_);
  or (_18498_, _18497_, _18493_);
  or (_18499_, _18498_, _10779_);
  or (_18500_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_18501_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_18502_, _18501_, _18500_);
  and (_18503_, _18502_, _04847_);
  or (_18504_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_18505_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_18506_, _18505_, _18504_);
  and (_18507_, _18506_, _10786_);
  or (_18508_, _18507_, _18503_);
  or (_18509_, _18508_, _04870_);
  and (_18510_, _18509_, _04880_);
  and (_18511_, _18510_, _18499_);
  or (_18512_, _18511_, _18489_);
  and (_18513_, _18512_, _04851_);
  or (_18514_, _18513_, _18467_);
  and (_18515_, _18514_, _10849_);
  or (_18516_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_18517_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_18518_, _18517_, _18516_);
  and (_18519_, _18518_, _04847_);
  or (_18520_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_18521_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_18522_, _18521_, _18520_);
  and (_18523_, _18522_, _10786_);
  or (_18524_, _18523_, _18519_);
  and (_18525_, _18524_, _10779_);
  or (_18526_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_18527_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_18528_, _18527_, _18526_);
  and (_18529_, _18528_, _04847_);
  or (_18530_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_18531_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_18532_, _18531_, _18530_);
  and (_18533_, _18532_, _10786_);
  or (_18534_, _18533_, _18529_);
  and (_18535_, _18534_, _04870_);
  or (_18536_, _18535_, _18525_);
  and (_18537_, _18536_, _04880_);
  and (_18538_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_18539_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_18540_, _18539_, _18538_);
  and (_18541_, _18540_, _04847_);
  and (_18542_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_18543_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_18544_, _18543_, _18542_);
  and (_18545_, _18544_, _10786_);
  or (_18546_, _18545_, _18541_);
  and (_18547_, _18546_, _10779_);
  and (_18548_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_18549_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_18550_, _18549_, _18548_);
  and (_18551_, _18550_, _04847_);
  and (_18552_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_18553_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_18554_, _18553_, _18552_);
  and (_18555_, _18554_, _10786_);
  or (_18556_, _18555_, _18551_);
  and (_18557_, _18556_, _04870_);
  or (_18558_, _18557_, _18547_);
  and (_18559_, _18558_, _10795_);
  or (_18560_, _18559_, _18537_);
  and (_18561_, _18560_, _04851_);
  or (_18562_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_18563_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_18564_, _18563_, _10786_);
  and (_18565_, _18564_, _18562_);
  or (_18566_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_18567_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_18568_, _18567_, _04847_);
  and (_18569_, _18568_, _18566_);
  or (_18570_, _18569_, _18565_);
  and (_18571_, _18570_, _10779_);
  or (_18572_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_18573_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_18574_, _18573_, _10786_);
  and (_18575_, _18574_, _18572_);
  or (_18576_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_18577_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_18578_, _18577_, _04847_);
  and (_18579_, _18578_, _18576_);
  or (_18580_, _18579_, _18575_);
  and (_18581_, _18580_, _04870_);
  or (_18582_, _18581_, _18571_);
  and (_18583_, _18582_, _04880_);
  and (_18584_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_18585_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_18586_, _18585_, _18584_);
  and (_18587_, _18586_, _04847_);
  and (_18588_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_18589_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_18590_, _18589_, _18588_);
  and (_18591_, _18590_, _10786_);
  or (_18592_, _18591_, _18587_);
  and (_18593_, _18592_, _10779_);
  and (_18594_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_18595_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_18596_, _18595_, _18594_);
  and (_18597_, _18596_, _04847_);
  and (_18598_, _10780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_18599_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_18600_, _18599_, _18598_);
  and (_18601_, _18600_, _10786_);
  or (_18602_, _18601_, _18597_);
  and (_18603_, _18602_, _04870_);
  or (_18604_, _18603_, _18593_);
  and (_18605_, _18604_, _10795_);
  or (_18606_, _18605_, _18583_);
  and (_18607_, _18606_, _10777_);
  or (_18608_, _18607_, _18561_);
  and (_18609_, _18608_, _04853_);
  or (_18610_, _18609_, _18515_);
  or (_18611_, _18610_, _11038_);
  and (_18612_, _18611_, _18421_);
  or (_18613_, _18612_, _03372_);
  and (_18614_, _18613_, _18231_);
  or (_18615_, _18614_, _04902_);
  or (_18616_, _11760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_18617_, _18616_, _23049_);
  and (_08896_, _18617_, _18615_);
  and (_18618_, _17846_, _23830_);
  and (_18619_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_08898_, _18619_, _18618_);
  and (_18620_, _17822_, _25886_);
  and (_18621_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or (_08900_, _18621_, _18620_);
  and (_18622_, _10284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  and (_18623_, _10283_, _23768_);
  or (_08904_, _18623_, _18622_);
  and (_18624_, _05557_, _26170_);
  and (_18625_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_08908_, _18625_, _18624_);
  and (_18626_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  and (_18627_, _06369_, _23768_);
  or (_08910_, _18627_, _18626_);
  and (_18628_, _26355_, _26202_);
  and (_18629_, _18628_, _25886_);
  not (_18630_, _18628_);
  and (_18631_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_27298_, _18631_, _18629_);
  and (_18632_, _26355_, _23220_);
  and (_18633_, _18632_, _23830_);
  not (_18634_, _18632_);
  and (_18635_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_08920_, _18635_, _18633_);
  and (_18636_, _18632_, _23768_);
  and (_18637_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_08922_, _18637_, _18636_);
  and (_18638_, _26355_, _26072_);
  and (_18639_, _18638_, _26242_);
  not (_18640_, _18638_);
  and (_18641_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_08925_, _18641_, _18639_);
  and (_18642_, _18638_, _25886_);
  and (_18643_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_08929_, _18643_, _18642_);
  and (_18644_, _14392_, _26185_);
  and (_18645_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_08931_, _18645_, _18644_);
  and (_18646_, _14388_, _23768_);
  and (_18647_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or (_08933_, _18647_, _18646_);
  and (_18648_, _04096_, _25886_);
  and (_18649_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_08935_, _18649_, _18648_);
  and (_18650_, _26355_, _26340_);
  and (_18651_, _18650_, _26185_);
  not (_18652_, _18650_);
  and (_18653_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_08941_, _18653_, _18651_);
  and (_18654_, _15231_, _25886_);
  and (_18655_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_27238_, _18655_, _18654_);
  and (_18656_, _17822_, _23830_);
  and (_18657_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or (_08984_, _18657_, _18656_);
  and (_18658_, _17822_, _26242_);
  and (_18659_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or (_27249_, _18659_, _18658_);
  and (_18660_, _05557_, _25886_);
  and (_18661_, _05559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or (_08987_, _18661_, _18660_);
  and (_18662_, _17822_, _26185_);
  and (_18663_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or (_08990_, _18663_, _18662_);
  and (_18664_, _17822_, _26085_);
  and (_18665_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or (_08992_, _18665_, _18664_);
  and (_18666_, _09128_, _25886_);
  and (_18667_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  or (_08997_, _18667_, _18666_);
  and (_18668_, _09128_, _26085_);
  and (_18669_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  or (_09000_, _18669_, _18668_);
  and (_18670_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_18671_, _10259_, _23768_);
  or (_09002_, _18671_, _18670_);
  and (_18672_, _18650_, _26170_);
  and (_18673_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_09010_, _18673_, _18672_);
  and (_18674_, _18650_, _23768_);
  and (_18675_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_09012_, _18675_, _18674_);
  and (_18676_, _26421_, _26355_);
  and (_18677_, _18676_, _26242_);
  not (_18678_, _18676_);
  and (_18679_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_09015_, _18679_, _18677_);
  and (_18680_, _18676_, _23830_);
  and (_18681_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_27293_, _18681_, _18680_);
  and (_18682_, _18676_, _23768_);
  and (_18683_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_09020_, _18683_, _18682_);
  and (_18684_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_18685_, _09450_, _26242_);
  or (_27089_, _18685_, _18684_);
  and (_18686_, _26355_, _26150_);
  and (_18687_, _18686_, _25927_);
  not (_18688_, _18686_);
  and (_18689_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_09024_, _18689_, _18687_);
  and (_18690_, _14392_, _26242_);
  and (_18691_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_09027_, _18691_, _18690_);
  and (_18692_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  and (_18693_, _04143_, _26085_);
  or (_09030_, _18693_, _18692_);
  and (_18694_, _26355_, _25932_);
  and (_18695_, _18694_, _26085_);
  not (_18696_, _18694_);
  and (_18697_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_09036_, _18697_, _18695_);
  and (_18698_, _04096_, _26170_);
  and (_18699_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_09038_, _18699_, _18698_);
  and (_18700_, _14558_, _25886_);
  and (_18701_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or (_09039_, _18701_, _18700_);
  and (_18702_, _18694_, _26170_);
  and (_18703_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_09046_, _18703_, _18702_);
  and (_18704_, _26202_, _25938_);
  and (_18705_, _18704_, _26185_);
  not (_18706_, _18704_);
  and (_18707_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_09048_, _18707_, _18705_);
  and (_18708_, _17830_, _25886_);
  and (_18709_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_09051_, _18709_, _18708_);
  and (_18710_, _18704_, _26085_);
  and (_18711_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_09055_, _18711_, _18710_);
  and (_18712_, _10455_, _26170_);
  and (_18713_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_26973_, _18713_, _18712_);
  and (_18714_, _18704_, _23830_);
  and (_18715_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_09058_, _18715_, _18714_);
  and (_18716_, _18704_, _25886_);
  and (_18717_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_09060_, _18717_, _18716_);
  and (_18718_, _17840_, _26242_);
  and (_18719_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_09063_, _18719_, _18718_);
  nand (_18720_, _02406_, _25279_);
  or (_18721_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_18722_, _18721_, _23049_);
  and (_09065_, _18722_, _18720_);
  and (_18723_, _18628_, _26085_);
  and (_18724_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_09071_, _18724_, _18723_);
  and (_18725_, _18628_, _25927_);
  and (_18726_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_09073_, _18726_, _18725_);
  and (_18727_, _18632_, _26185_);
  and (_18728_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_09075_, _18728_, _18727_);
  and (_18729_, _18676_, _26170_);
  and (_18730_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_09081_, _18730_, _18729_);
  and (_18731_, _18686_, _26242_);
  and (_18732_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_09083_, _18732_, _18731_);
  and (_18733_, _18686_, _23830_);
  and (_18734_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_09086_, _18734_, _18733_);
  and (_18735_, _18638_, _23768_);
  and (_18736_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_09088_, _18736_, _18735_);
  nand (_18737_, _02406_, _23761_);
  or (_18738_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_18739_, _18738_, _23049_);
  and (_09091_, _18739_, _18737_);
  and (_18740_, _17834_, _26185_);
  and (_18741_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_09093_, _18741_, _18740_);
  and (_18742_, _17840_, _23768_);
  and (_18743_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_09096_, _18743_, _18742_);
  and (_18744_, _17846_, _23768_);
  and (_18745_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_27301_, _18745_, _18744_);
  and (_18746_, _05799_, _26242_);
  and (_18747_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_09099_, _18747_, _18746_);
  and (_18748_, _26542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  and (_18749_, _26541_, _26185_);
  or (_09101_, _18749_, _18748_);
  and (_18750_, _14388_, _23830_);
  and (_18751_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_09105_, _18751_, _18750_);
  and (_18752_, _14388_, _25886_);
  and (_18753_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or (_09108_, _18753_, _18752_);
  and (_18754_, _14388_, _26170_);
  and (_18755_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_09109_, _18755_, _18754_);
  and (_18756_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_18757_, _10259_, _26170_);
  or (_09145_, _18757_, _18756_);
  and (_18758_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_18759_, _09304_, _23768_);
  or (_09147_, _18759_, _18758_);
  and (_18760_, _10455_, _26085_);
  and (_18761_, _10457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_09157_, _18761_, _18760_);
  and (_18762_, _10260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_18763_, _10259_, _25886_);
  or (_27093_, _18763_, _18762_);
  and (_18764_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  and (_18765_, _02576_, _26242_);
  or (_27079_, _18765_, _18764_);
  and (_18766_, _04812_, _23830_);
  and (_18767_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or (_27107_, _18767_, _18766_);
  and (_18768_, _09128_, _26242_);
  and (_18769_, _09130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or (_09183_, _18769_, _18768_);
  and (_18770_, _17822_, _23768_);
  and (_18771_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or (_09185_, _18771_, _18770_);
  and (_18772_, _26224_, _23848_);
  and (_18773_, _18772_, _26170_);
  not (_18774_, _18772_);
  and (_18775_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_09210_, _18775_, _18773_);
  and (_18776_, _09122_, _23768_);
  and (_18777_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_09219_, _18777_, _18776_);
  and (_18778_, _18772_, _23830_);
  and (_18779_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_09238_, _18779_, _18778_);
  and (_18780_, _18772_, _25886_);
  and (_18781_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_09303_, _18781_, _18780_);
  and (_18782_, _09122_, _25886_);
  and (_18783_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_09329_, _18783_, _18782_);
  and (_18784_, _09122_, _26085_);
  and (_18785_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_09359_, _18785_, _18784_);
  and (_18786_, _09122_, _26242_);
  and (_18787_, _09124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_27159_, _18787_, _18786_);
  and (_18788_, _01871_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nand (_18789_, _25059_, _25095_);
  or (_18790_, _15196_, _03526_);
  or (_18791_, _18790_, _15205_);
  or (_18792_, _18791_, _18789_);
  and (_18793_, _18792_, _22836_);
  not (_18794_, _24145_);
  or (_18795_, _18794_, _25101_);
  or (_18796_, _15384_, _01901_);
  or (_18797_, _18796_, _18795_);
  and (_18798_, _23052_, _23032_);
  or (_18799_, _09032_, _24154_);
  or (_18800_, _18799_, _18798_);
  or (_18801_, _18800_, _01889_);
  or (_18802_, _18801_, _09031_);
  or (_18803_, _18802_, _18797_);
  or (_18804_, _18803_, _18793_);
  and (_18805_, _18804_, _01913_);
  or (_26899_[0], _18805_, _18788_);
  and (_18806_, _00115_, _26085_);
  and (_18807_, _00117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_09426_, _18807_, _18806_);
  and (_18808_, _10724_, _26185_);
  and (_18809_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_09429_, _18809_, _18808_);
  and (_18810_, _10463_, _25886_);
  and (_18811_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_09430_, _18811_, _18810_);
  and (_18812_, _10463_, _23768_);
  and (_18813_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_09433_, _18813_, _18812_);
  and (_18814_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  and (_18815_, _06369_, _25886_);
  or (_09443_, _18815_, _18814_);
  and (_18816_, _10724_, _26170_);
  and (_18817_, _10726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_09445_, _18817_, _18816_);
  and (_18818_, _10463_, _23830_);
  and (_18819_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_09447_, _18819_, _18818_);
  and (_18820_, _09756_, _25886_);
  and (_18821_, _09758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_09458_, _18821_, _18820_);
  and (_18822_, _10463_, _26085_);
  and (_18823_, _10465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_27001_, _18823_, _18822_);
  and (_18824_, _23840_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_18825_, _18824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_26926_[7], _18825_, _23049_);
  and (_18826_, _26615_, _26185_);
  and (_18827_, _26617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_27272_, _18827_, _18826_);
  or (_18828_, _25080_, _23031_);
  or (_18829_, _18828_, _15291_);
  or (_18830_, _18829_, _15279_);
  and (_18831_, _18830_, _22739_);
  and (_18832_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_18833_, _18832_, _15301_);
  or (_18834_, _18833_, _18831_);
  and (_26900_[0], _18834_, _23049_);
  and (_18835_, _18704_, _26242_);
  and (_18836_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_09530_, _18836_, _18835_);
  and (_18837_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18838_, _25096_, _22973_);
  or (_18839_, _18838_, _23021_);
  or (_18840_, _18839_, _15288_);
  or (_18841_, _18840_, _08641_);
  and (_18842_, _18841_, _22739_);
  or (_18843_, _18842_, _18837_);
  or (_18844_, _18843_, _15300_);
  and (_26900_[1], _18844_, _23049_);
  and (_18845_, _17846_, _25927_);
  and (_18846_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_09582_, _18846_, _18845_);
  or (_18847_, _14971_, _00773_);
  or (_18848_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18849_, _18848_, _25128_);
  and (_18850_, _18849_, _18847_);
  and (_18852_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18853_, _14977_, _26136_);
  nand (_18854_, _18853_, _23729_);
  or (_18855_, _18853_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18856_, _18855_, _25618_);
  and (_18857_, _18856_, _18854_);
  or (_18858_, _18857_, _18852_);
  or (_18859_, _18858_, _18850_);
  and (_09585_, _18859_, _23049_);
  and (_18860_, _10475_, _23768_);
  and (_18861_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_09590_, _18861_, _18860_);
  and (_18862_, _00049_, _23830_);
  and (_18863_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_09591_, _18863_, _18862_);
  and (_18864_, _26375_, _26202_);
  and (_18865_, _18864_, _26085_);
  not (_18866_, _18864_);
  and (_18867_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_09602_, _18867_, _18865_);
  and (_18868_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  and (_18869_, _00089_, _25886_);
  or (_09604_, _18869_, _18868_);
  and (_18870_, _18864_, _26170_);
  and (_18871_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_27321_, _18871_, _18870_);
  and (_18872_, _23008_, _22972_);
  and (_18873_, _18872_, _23052_);
  or (_18874_, _18873_, _23053_);
  or (_18875_, _18874_, _15382_);
  or (_18876_, _09032_, _24155_);
  or (_18877_, _18876_, _18875_);
  or (_18878_, _08650_, _23054_);
  and (_18879_, _25585_, _01873_);
  or (_18880_, _18879_, _18878_);
  and (_18881_, _23052_, _25071_);
  or (_18882_, _15205_, _15199_);
  or (_18883_, _18882_, _18881_);
  or (_18884_, _18883_, _22996_);
  or (_18885_, _18884_, _18880_);
  or (_18886_, _18885_, _18877_);
  and (_18887_, _23052_, _22940_);
  or (_18888_, _15286_, _01883_);
  or (_18889_, _18888_, _18887_);
  or (_18890_, _15281_, _15389_);
  or (_18891_, _18890_, _22985_);
  or (_18892_, _18891_, _18889_);
  or (_18893_, _18892_, _15369_);
  and (_18894_, _15271_, _23008_);
  and (_18895_, _23027_, _22994_);
  and (_18896_, _15196_, _22973_);
  or (_18897_, _18896_, _18895_);
  or (_18898_, _18897_, _18894_);
  or (_18899_, _18898_, _08641_);
  or (_18900_, _18899_, _18893_);
  or (_18901_, _18900_, _18886_);
  and (_18902_, _18901_, _22739_);
  and (_18903_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_18904_, _15209_, _08654_);
  or (_18905_, _18904_, _18903_);
  or (_18906_, _18905_, _18902_);
  and (_26901_[0], _18906_, _23049_);
  and (_18907_, _18864_, _23768_);
  and (_18908_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_09607_, _18908_, _18907_);
  and (_18909_, _26375_, _23220_);
  and (_18910_, _18909_, _26242_);
  not (_18911_, _18909_);
  and (_18912_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_09609_, _18912_, _18910_);
  and (_18913_, _24164_, _23008_);
  or (_18914_, _18913_, _25080_);
  and (_18915_, _23008_, _23000_);
  or (_18916_, _18915_, _15253_);
  nor (_18917_, _18916_, _18914_);
  nand (_18918_, _18917_, _22986_);
  and (_18919_, _18789_, _22835_);
  or (_18920_, _18919_, _15369_);
  or (_18921_, _18920_, _18918_);
  or (_18922_, _23054_, _23023_);
  or (_18923_, _15272_, _25102_);
  or (_18924_, _18923_, _18922_);
  or (_18925_, _18924_, _18884_);
  or (_18926_, _18925_, _18877_);
  or (_18927_, _18926_, _18921_);
  and (_18928_, _18927_, _22739_);
  and (_18929_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_18930_, _18929_, _18904_);
  or (_18931_, _18930_, _18928_);
  and (_26901_[1], _18931_, _23049_);
  and (_18932_, _26301_, _25886_);
  and (_18933_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_09613_, _18933_, _18932_);
  and (_18934_, _18909_, _26085_);
  and (_18935_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_09615_, _18935_, _18934_);
  or (_18936_, _14971_, _00557_);
  or (_18937_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18938_, _18937_, _25128_);
  and (_18939_, _18938_, _18936_);
  and (_18940_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18941_, _14977_, _25224_);
  nand (_18942_, _18941_, _23729_);
  or (_18943_, _18941_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18944_, _18943_, _25618_);
  and (_18945_, _18944_, _18942_);
  or (_18946_, _18945_, _18940_);
  or (_18947_, _18946_, _18939_);
  and (_09617_, _18947_, _23049_);
  and (_18948_, _18909_, _25927_);
  and (_18949_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_27320_, _18949_, _18948_);
  and (_18950_, _26375_, _26072_);
  and (_18951_, _18950_, _25886_);
  not (_18952_, _18950_);
  and (_18953_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_09626_, _18953_, _18951_);
  and (_18954_, _18950_, _23768_);
  and (_18955_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_09630_, _18955_, _18954_);
  and (_18956_, _26375_, _25932_);
  and (_18957_, _18956_, _23830_);
  not (_18958_, _18956_);
  and (_18959_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_27317_, _18959_, _18957_);
  and (_18960_, _14388_, _25927_);
  and (_18961_, _14390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_09636_, _18961_, _18960_);
  and (_18962_, _18956_, _26170_);
  and (_18963_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_09638_, _18963_, _18962_);
  nand (_18964_, _14970_, _00608_);
  or (_18965_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_18966_, _18965_, _25128_);
  and (_18967_, _18966_, _18964_);
  and (_18968_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_18969_, _14977_, _25905_);
  and (_18970_, _18969_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_18971_, _25223_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_18972_, _18971_, _25896_);
  and (_18973_, _18972_, _14977_);
  or (_18974_, _18973_, _18970_);
  and (_18975_, _18974_, _25618_);
  or (_18976_, _18975_, _18968_);
  or (_18977_, _18976_, _18967_);
  and (_09640_, _18977_, _23049_);
  and (_18978_, _04096_, _26085_);
  and (_18979_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_09653_, _18979_, _18978_);
  and (_18980_, _25938_, _23220_);
  and (_18981_, _18980_, _26185_);
  not (_18982_, _18980_);
  and (_18983_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_09655_, _18983_, _18981_);
  and (_18984_, _26375_, _26340_);
  and (_18985_, _18984_, _26085_);
  not (_18986_, _18984_);
  and (_18987_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_09660_, _18987_, _18985_);
  and (_18988_, _18984_, _25886_);
  and (_18989_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_09662_, _18989_, _18988_);
  and (_18990_, _26421_, _26375_);
  and (_18991_, _18990_, _26185_);
  not (_18992_, _18990_);
  and (_18993_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_09671_, _18993_, _18991_);
  and (_18994_, _18990_, _23830_);
  and (_18995_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_27316_, _18995_, _18994_);
  or (_18996_, _14971_, _00659_);
  or (_18997_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_18998_, _18997_, _25128_);
  and (_18999_, _18998_, _18996_);
  and (_19000_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_19001_, _14977_, _26473_);
  nand (_19002_, _19001_, _23729_);
  or (_19003_, _19001_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_19004_, _19003_, _25618_);
  and (_19005_, _19004_, _19002_);
  or (_19006_, _19005_, _19000_);
  or (_19007_, _19006_, _18999_);
  and (_09674_, _19007_, _23049_);
  or (_19008_, _14971_, _00713_);
  or (_19009_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_19010_, _19009_, _25128_);
  and (_19011_, _19010_, _19008_);
  and (_19012_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_19013_, _14977_);
  or (_19014_, _19013_, _26563_);
  and (_19015_, _19014_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_19016_, _23215_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_19017_, _19016_, _26557_);
  and (_19018_, _19017_, _14977_);
  or (_19019_, _19018_, _19015_);
  and (_19020_, _19019_, _25618_);
  or (_19021_, _19020_, _19012_);
  or (_19022_, _19021_, _19011_);
  and (_09677_, _19022_, _23049_);
  and (_19023_, _18990_, _23768_);
  and (_19024_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_09678_, _19024_, _19023_);
  and (_19025_, _26375_, _26150_);
  and (_19026_, _19025_, _26242_);
  not (_19027_, _19025_);
  and (_19028_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_09681_, _19028_, _19026_);
  and (_19029_, _19025_, _26085_);
  and (_19030_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_09683_, _19030_, _19029_);
  and (_09699_, _25419_, _23049_);
  and (_09701_, _26941_, _25215_);
  and (_19031_, _26375_, _26283_);
  and (_19032_, _19031_, _25927_);
  not (_19033_, _19031_);
  and (_19034_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_09703_, _19034_, _19032_);
  and (_19035_, _02519_, _26242_);
  and (_19036_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_09708_, _19036_, _19035_);
  and (_19037_, _04096_, _23830_);
  and (_19038_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_09710_, _19038_, _19037_);
  and (_19039_, _26375_, _23847_);
  and (_19040_, _19039_, _26170_);
  not (_19041_, _19039_);
  and (_19042_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_27309_, _19042_, _19040_);
  and (_19043_, _19039_, _23768_);
  and (_19044_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_09717_, _19044_, _19043_);
  and (_19045_, _26432_, _26242_);
  and (_19046_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_27308_, _19046_, _19045_);
  and (_19047_, _14392_, _23768_);
  and (_19048_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_09727_, _19048_, _19047_);
  and (_19049_, _01871_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_19050_, _24146_, _22949_);
  nor (_19051_, _03987_, _19050_);
  nand (_19052_, _19051_, _02672_);
  or (_19053_, _19052_, _15205_);
  or (_19054_, _03543_, _15389_);
  or (_19055_, _03995_, _03994_);
  nor (_19056_, _19055_, _19054_);
  nand (_19057_, _19056_, _25065_);
  or (_19058_, _15276_, _03993_);
  or (_19059_, _19058_, _19057_);
  or (_19060_, _01873_, _24143_);
  and (_19061_, _19060_, _25584_);
  and (_19062_, _23052_, _23018_);
  or (_19063_, _19062_, _01896_);
  and (_19064_, _15198_, _22972_);
  or (_19065_, _19064_, _19063_);
  or (_19066_, _19065_, _19061_);
  and (_19067_, _24141_, _22949_);
  or (_19068_, _19067_, _25090_);
  and (_19069_, _25584_, _22949_);
  or (_19070_, _15199_, _03988_);
  or (_19071_, _19070_, _19069_);
  or (_19072_, _19071_, _19068_);
  or (_19073_, _19072_, _19066_);
  or (_19074_, _19073_, _19059_);
  or (_19075_, _19074_, _19053_);
  and (_19076_, _19075_, _01913_);
  or (_26902_[0], _19076_, _19049_);
  and (_19077_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_19078_, _09450_, _25927_);
  or (_09738_, _19078_, _19077_);
  and (_19079_, _26432_, _25886_);
  and (_19080_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_09740_, _19080_, _19079_);
  and (_19081_, _26375_, _26224_);
  and (_19082_, _19081_, _23830_);
  not (_19083_, _19081_);
  and (_19084_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_09745_, _19084_, _19082_);
  and (_19085_, _18980_, _26085_);
  and (_19086_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_09747_, _19086_, _19085_);
  and (_19087_, _06370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  and (_19088_, _06369_, _26170_);
  or (_09749_, _19088_, _19087_);
  and (_19089_, _19081_, _26170_);
  and (_19090_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_09751_, _19090_, _19089_);
  and (_19091_, _18864_, _26242_);
  and (_19092_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_09753_, _19092_, _19091_);
  and (_19093_, _00419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  and (_19094_, _00418_, _26242_);
  or (_27064_, _19094_, _19093_);
  and (_19095_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_19096_, _09450_, _23768_);
  or (_09764_, _19096_, _19095_);
  and (_19097_, _18956_, _26185_);
  and (_19098_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_27319_, _19098_, _19097_);
  and (_19099_, _18984_, _26242_);
  and (_19100_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_09767_, _19100_, _19099_);
  or (_19101_, _14971_, _00500_);
  or (_19102_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_19103_, _19102_, _25128_);
  and (_19104_, _19103_, _19101_);
  and (_19105_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_19106_, _14970_, _23729_);
  and (_19107_, _19102_, _25618_);
  and (_19108_, _19107_, _19106_);
  or (_19109_, _19108_, _19105_);
  or (_19110_, _19109_, _19104_);
  and (_09774_, _19110_, _23049_);
  and (_19111_, _14392_, _26170_);
  and (_19112_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_09778_, _19112_, _19111_);
  and (_19113_, _04202_, _26085_);
  and (_19114_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_09779_, _19114_, _19113_);
  and (_19115_, _14392_, _23830_);
  and (_19116_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_09783_, _19116_, _19115_);
  and (_19117_, _19039_, _23830_);
  and (_19118_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_09785_, _19118_, _19117_);
  or (_19119_, _14971_, _00836_);
  or (_19120_, _14970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_19121_, _19120_, _25128_);
  and (_19122_, _19121_, _19119_);
  and (_19123_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_19124_, _14977_, _26524_);
  nand (_19125_, _19124_, _23729_);
  or (_19126_, _19124_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_19127_, _19126_, _25618_);
  and (_19128_, _19127_, _19125_);
  or (_19129_, _19128_, _19123_);
  or (_19130_, _19129_, _19122_);
  and (_09790_, _19130_, _23049_);
  and (_19131_, _01871_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_19132_, _19062_, _19069_);
  or (_19133_, _19132_, _19050_);
  not (_19134_, _25081_);
  or (_19135_, _01885_, _19134_);
  or (_19136_, _19135_, _19133_);
  or (_19137_, _01886_, _22996_);
  or (_19138_, _18896_, _15368_);
  or (_19139_, _19138_, _19137_);
  or (_19140_, _22985_, _22977_);
  or (_19141_, _01899_, _23061_);
  or (_19142_, _19141_, _25061_);
  or (_19143_, _01887_, _01875_);
  or (_19144_, _19143_, _19142_);
  or (_19145_, _19144_, _19140_);
  or (_19146_, _19145_, _19139_);
  or (_19147_, _19146_, _18880_);
  or (_19148_, _19147_, _19136_);
  or (_19149_, _23054_, _23040_);
  nor (_19150_, rst, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_19151_, _19150_, _19149_);
  and (_19152_, _19151_, _19148_);
  or (_26903_[0], _19152_, _19131_);
  and (_19153_, _19025_, _25927_);
  and (_19154_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_27312_, _19154_, _19153_);
  and (_19155_, _19081_, _26185_);
  and (_19156_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_09802_, _19156_, _19155_);
  and (_19157_, _15146_, _26170_);
  and (_19158_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_27277_, _19158_, _19157_);
  and (_19159_, _14392_, _25886_);
  and (_19160_, _14394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_09812_, _19160_, _19159_);
  nand (_09828_, _25665_, _23049_);
  and (_19161_, _18909_, _26170_);
  and (_19162_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_09830_, _19162_, _19161_);
  and (_19163_, _01997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  and (_19164_, _01996_, _26085_);
  or (_09833_, _19164_, _19163_);
  and (_19165_, _09667_, _26085_);
  and (_19166_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_09834_, _19166_, _19165_);
  and (_19167_, _18990_, _25927_);
  and (_19168_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_09843_, _19168_, _19167_);
  nor (_09848_, _25295_, rst);
  and (_19169_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  and (_19170_, _10218_, _26242_);
  or (_09850_, _19170_, _19169_);
  nor (_09878_, _25374_, rst);
  nand (_09880_, _25702_, _23049_);
  or (_19171_, _03526_, _25080_);
  or (_19172_, _19171_, _25079_);
  and (_19173_, _24141_, _24143_);
  or (_19174_, _01875_, _19173_);
  or (_19175_, _19174_, _15205_);
  or (_19176_, _19175_, _19172_);
  or (_19177_, _19176_, _15252_);
  and (_19178_, _03538_, _22972_);
  or (_19179_, _19178_, _15375_);
  and (_19180_, _22992_, _22949_);
  and (_19181_, _24141_, _22948_);
  or (_19182_, _19181_, _18873_);
  or (_19183_, _19182_, _19180_);
  or (_19184_, _19183_, _19179_);
  and (_19185_, _01873_, _24141_);
  or (_19186_, _09032_, _19185_);
  or (_19187_, _25063_, _23021_);
  or (_19188_, _19187_, _19186_);
  or (_19189_, _19070_, _18922_);
  or (_19190_, _19189_, _19188_);
  or (_19191_, _19190_, _19184_);
  or (_19192_, _19191_, _01897_);
  or (_19193_, _19192_, _19177_);
  and (_19194_, _19193_, _19151_);
  and (_19195_, _01871_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_26903_[1], _19195_, _19194_);
  and (_19196_, _22997_, _22949_);
  or (_19197_, _19063_, _19196_);
  or (_19198_, _19182_, _19179_);
  or (_19199_, _19198_, _19197_);
  or (_19200_, _23021_, _22998_);
  or (_19201_, _19200_, _01907_);
  or (_19202_, _03989_, _19171_);
  or (_19203_, _19202_, _19201_);
  not (_19204_, _02672_);
  or (_19205_, _19204_, _01895_);
  or (_19206_, _19205_, _19203_);
  or (_19207_, _19206_, _19199_);
  and (_19208_, _19207_, _22739_);
  and (_19209_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_19210_, _23053_, _22734_);
  or (_19211_, _19210_, _19209_);
  or (_19212_, _19211_, _19208_);
  and (_26903_[2], _19212_, _23049_);
  and (_19213_, _18956_, _26242_);
  and (_19214_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_09902_, _19214_, _19213_);
  and (_19215_, _18984_, _23768_);
  and (_19216_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_09907_, _19216_, _19215_);
  and (_19217_, _19039_, _26085_);
  and (_19218_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_09910_, _19218_, _19217_);
  and (_19219_, _19025_, _26170_);
  and (_19220_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_09912_, _19220_, _19219_);
  and (_19221_, _04825_, _26185_);
  and (_19222_, _04827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or (_09920_, _19222_, _19221_);
  and (_19223_, _14665_, _26185_);
  and (_19224_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_09925_, _19224_, _19223_);
  nand (_09927_, _25719_, _23049_);
  nor (_09929_, _25497_, rst);
  nor (_09930_, _25455_, rst);
  and (_19225_, _19081_, _25927_);
  and (_19226_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_09934_, _19226_, _19225_);
  and (_19227_, _18694_, _25927_);
  and (_19228_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_27296_, _19228_, _19227_);
  and (_19229_, _26284_, _26242_);
  and (_19230_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_09938_, _19230_, _19229_);
  and (_19231_, _18650_, _26242_);
  and (_19232_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_09941_, _19232_, _19231_);
  and (_19233_, _19031_, _26242_);
  and (_19234_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_09947_, _19234_, _19233_);
  and (_19235_, _14665_, _26085_);
  and (_19236_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_09949_, _19236_, _19235_);
  and (_19237_, _26301_, _26242_);
  and (_19238_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_09951_, _19238_, _19237_);
  and (_19239_, _14665_, _23830_);
  and (_19240_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_09953_, _19240_, _19239_);
  and (_19241_, _19081_, _23768_);
  and (_19242_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_09955_, _19242_, _19241_);
  and (_19243_, _18694_, _23768_);
  and (_19244_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_09957_, _19244_, _19243_);
  and (_19245_, _14665_, _25886_);
  and (_19246_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_09959_, _19246_, _19245_);
  and (_19247_, _26176_, _26170_);
  and (_19248_, _26188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_26971_, _19248_, _19247_);
  not (_19249_, _03819_);
  nor (_19250_, _19249_, _01012_);
  and (_19251_, _26473_, _25227_);
  nand (_19252_, _19251_, _00608_);
  or (_19253_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_19254_, _19253_, _19249_);
  and (_19255_, _19254_, _19252_);
  or (_19256_, _19255_, _19250_);
  and (_09969_, _19256_, _23049_);
  and (_19257_, _25894_, _25227_);
  nor (_19258_, _19257_, _03819_);
  or (_19259_, _19258_, _00500_);
  not (_19260_, _19258_);
  or (_19261_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_19262_, _19261_, _23049_);
  and (_09971_, _19262_, _19259_);
  and (_19263_, _18704_, _25927_);
  and (_19264_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_09974_, _19264_, _19263_);
  and (_19265_, _26284_, _26170_);
  and (_19266_, _26286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_09984_, _19266_, _19265_);
  and (_19267_, _09667_, _26170_);
  and (_19268_, _09669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_09985_, _19268_, _19267_);
  and (_19269_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  and (_19270_, _00089_, _26085_);
  or (_09990_, _19270_, _19269_);
  and (_19271_, _19081_, _25886_);
  and (_19272_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_09993_, _19272_, _19271_);
  and (_19273_, _18694_, _25886_);
  and (_19274_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_09995_, _19274_, _19273_);
  and (_19275_, _04096_, _23768_);
  and (_19276_, _04098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_09997_, _19276_, _19275_);
  and (_19277_, _01871_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_19278_, _19185_, _25088_);
  nand (_19279_, _19278_, _25065_);
  or (_19280_, _19279_, _19132_);
  or (_19281_, _09025_, _18794_);
  or (_19282_, _19281_, _19067_);
  or (_19283_, _19282_, _15203_);
  or (_19284_, _19283_, _19280_);
  or (_19285_, _19284_, _19053_);
  and (_19286_, _19285_, _01913_);
  or (_26904_[0], _19286_, _19277_);
  and (_19287_, _19081_, _26085_);
  and (_19288_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_27311_, _19288_, _19287_);
  nor (_19289_, _19249_, _01160_);
  not (_19290_, _19251_);
  or (_19291_, _19290_, _00773_);
  or (_19292_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_19293_, _19292_, _19249_);
  and (_19294_, _19293_, _19291_);
  or (_19295_, _19294_, _19289_);
  and (_10008_, _19295_, _23049_);
  or (_19296_, _19258_, _00659_);
  or (_19297_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_19298_, _19297_, _23049_);
  and (_10009_, _19298_, _19296_);
  and (_19299_, _18704_, _23768_);
  and (_19300_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_10017_, _19300_, _19299_);
  and (_19301_, _18694_, _23830_);
  and (_19302_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_10019_, _19302_, _19301_);
  and (_19303_, _19081_, _26242_);
  and (_19304_, _19083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_10022_, _19304_, _19303_);
  and (_19305_, _18694_, _26185_);
  and (_19306_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_10023_, _19306_, _19305_);
  and (_19307_, _26170_, _26151_);
  and (_19308_, _26153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_10027_, _19308_, _19307_);
  or (_19309_, _19258_, _00713_);
  or (_19310_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_19311_, _19310_, _23049_);
  and (_10035_, _19311_, _19309_);
  and (_19312_, _19025_, _23768_);
  and (_19313_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_10040_, _19313_, _19312_);
  and (_19314_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  and (_19315_, _04148_, _26085_);
  or (_27179_, _19315_, _19314_);
  and (_19317_, _04202_, _26242_);
  and (_19318_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_10045_, _19318_, _19317_);
  and (_19319_, _03819_, _00959_);
  or (_19320_, _19290_, _00557_);
  or (_19321_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_19322_, _19321_, _19249_);
  and (_19323_, _19322_, _19320_);
  or (_19324_, _19323_, _19319_);
  and (_10048_, _19324_, _23049_);
  and (_19325_, _03819_, _00910_);
  or (_19326_, _19290_, _00500_);
  or (_19327_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_19328_, _19327_, _19249_);
  and (_19329_, _19328_, _19326_);
  or (_19330_, _19329_, _19325_);
  and (_10051_, _19330_, _23049_);
  and (_19331_, _18694_, _26242_);
  and (_19332_, _18696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_10054_, _19332_, _19331_);
  and (_19333_, _26432_, _25927_);
  and (_19334_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_10058_, _19334_, _19333_);
  and (_19335_, _26458_, _26242_);
  and (_19336_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_10062_, _19336_, _19335_);
  and (_19337_, _26432_, _26170_);
  and (_19338_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_10068_, _19338_, _19337_);
  and (_19339_, _18686_, _23768_);
  and (_19340_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_10071_, _19340_, _19339_);
  or (_19341_, _19258_, _00836_);
  or (_19342_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_19343_, _19342_, _23049_);
  and (_10074_, _19343_, _19341_);
  and (_19344_, _26432_, _23830_);
  and (_19345_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_10076_, _19345_, _19344_);
  and (_19346_, _18686_, _26170_);
  and (_19347_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_10078_, _19347_, _19346_);
  and (_19348_, _26185_, _23231_);
  and (_19349_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_10081_, _19349_, _19348_);
  or (_19350_, _19258_, _00773_);
  or (_19351_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_19352_, _19351_, _23049_);
  and (_10083_, _19352_, _19350_);
  nand (_19353_, _00071_, _25279_);
  and (_19354_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_19355_, _19354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_19356_, _10307_, _01674_);
  and (_19357_, _19356_, _19355_);
  or (_19358_, _10293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_19359_, _10295_, _02503_);
  and (_19360_, _09310_, _01666_);
  and (_19361_, _19360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_19362_, _19361_, _10293_);
  or (_19363_, _19360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_19364_, _19363_, _01673_);
  and (_19365_, _19364_, _19362_);
  or (_19366_, _19365_, _19359_);
  and (_19367_, _19366_, _19358_);
  or (_19368_, _19367_, _19357_);
  or (_19369_, _19368_, _00071_);
  and (_19370_, _19369_, _00070_);
  and (_19371_, _19370_, _19353_);
  and (_19372_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_19373_, _19372_, _19371_);
  and (_10087_, _19373_, _23049_);
  and (_19374_, _26432_, _26085_);
  and (_19375_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_10095_, _19375_, _19374_);
  and (_19376_, _18686_, _25886_);
  and (_19377_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_10099_, _19377_, _19376_);
  and (_19378_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  and (_19379_, _09103_, _26170_);
  or (_10101_, _19379_, _19378_);
  and (_19381_, _18686_, _26085_);
  and (_19382_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_10105_, _19382_, _19381_);
  and (_19383_, _26432_, _26185_);
  and (_19384_, _26434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_10107_, _19384_, _19383_);
  and (_19385_, _14665_, _26242_);
  and (_19386_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_26999_, _19386_, _19385_);
  and (_19387_, _18772_, _26242_);
  and (_19388_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_10110_, _19388_, _19387_);
  and (_19389_, _18686_, _26185_);
  and (_19390_, _18688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_10114_, _19390_, _19389_);
  and (_19391_, _00049_, _26170_);
  and (_19392_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_10116_, _19392_, _19391_);
  and (_19393_, _15146_, _26242_);
  and (_19394_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_10117_, _19394_, _19393_);
  and (_19395_, _03819_, _01204_);
  or (_19396_, _19290_, _00836_);
  or (_19397_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_19398_, _19397_, _19249_);
  and (_19399_, _19398_, _19396_);
  or (_19400_, _19399_, _19395_);
  and (_10125_, _19400_, _23049_);
  and (_19401_, _00049_, _26185_);
  and (_19402_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_10129_, _19402_, _19401_);
  and (_19403_, _19039_, _25927_);
  and (_19404_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_10131_, _19404_, _19403_);
  or (_19405_, _19258_, _25053_);
  or (_19406_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_19407_, _19406_, _23049_);
  and (_10133_, _19407_, _19405_);
  and (_19408_, _00049_, _26085_);
  and (_19409_, _00051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_10136_, _19409_, _19408_);
  and (_19410_, _03819_, _01109_);
  or (_19411_, _19290_, _00713_);
  or (_19412_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_19413_, _19412_, _19249_);
  and (_19414_, _19413_, _19411_);
  or (_19415_, _19414_, _19410_);
  and (_10141_, _19415_, _23049_);
  nand (_19416_, _19260_, _00608_);
  or (_19417_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_19418_, _19417_, _23049_);
  and (_10142_, _19418_, _19416_);
  and (_19419_, _19039_, _25886_);
  and (_19420_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_10144_, _19420_, _19419_);
  and (_19421_, _18676_, _25927_);
  and (_19422_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_10146_, _19422_, _19421_);
  and (_19423_, _03204_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_19424_, _19423_, _03206_);
  and (_19425_, _19424_, _25630_);
  or (_19426_, _25630_, _25625_);
  nor (_19427_, _19426_, _23729_);
  and (_19428_, _25631_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_19429_, _19428_, _25135_);
  or (_19430_, _19429_, _19427_);
  or (_19431_, _19430_, _19425_);
  nand (_19432_, _25417_, _25135_);
  and (_19433_, _19432_, _23049_);
  and (_10149_, _19433_, _19431_);
  and (_19434_, _01371_, _23768_);
  and (_19435_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_10151_, _19435_, _19434_);
  and (_19436_, _19039_, _26185_);
  and (_19437_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_10153_, _19437_, _19436_);
  and (_19438_, _03819_, _25846_);
  or (_19439_, _19290_, _25053_);
  or (_19440_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_19441_, _19440_, _19249_);
  and (_19442_, _19441_, _19439_);
  or (_19443_, _19442_, _19438_);
  and (_10154_, _19443_, _23049_);
  and (_19444_, _03819_, _01059_);
  or (_19445_, _19290_, _00659_);
  or (_19446_, _19251_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_19447_, _19446_, _19249_);
  and (_19448_, _19447_, _19445_);
  or (_19449_, _19448_, _19444_);
  and (_10161_, _19449_, _23049_);
  or (_19451_, _19258_, _00557_);
  or (_19452_, _19260_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_19453_, _19452_, _23049_);
  and (_10163_, _19453_, _19451_);
  and (_19454_, _01371_, _26242_);
  and (_19455_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_10165_, _19455_, _19454_);
  and (_19456_, _18772_, _26185_);
  and (_19457_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_10168_, _19457_, _19456_);
  and (_19458_, _18676_, _25886_);
  and (_19459_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_10171_, _19459_, _19458_);
  or (_19460_, _02497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_19461_, _10293_, _02503_);
  and (_19462_, _19461_, _19460_);
  or (_19463_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_19464_, _19354_, _01674_);
  and (_19465_, _19464_, _19463_);
  not (_19466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_19467_, _01670_, _01666_);
  nor (_19468_, _19467_, _19466_);
  and (_19469_, _19467_, _19466_);
  or (_19470_, _19469_, _19468_);
  and (_19471_, _19470_, _01673_);
  or (_19472_, _19471_, _19465_);
  or (_19473_, _19472_, _19462_);
  or (_19474_, _19473_, _00071_);
  nand (_19475_, _00071_, _23761_);
  and (_19476_, _19475_, _19474_);
  or (_19477_, _19476_, _00069_);
  nand (_19478_, _00069_, _19466_);
  and (_19479_, _19478_, _23049_);
  and (_10174_, _19479_, _19477_);
  and (_19480_, _04202_, _23768_);
  and (_19481_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_10177_, _19481_, _19480_);
  and (_19482_, _18676_, _26085_);
  and (_19483_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_10179_, _19483_, _19482_);
  and (_19484_, _01604_, _25886_);
  and (_19485_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_10182_, _19485_, _19484_);
  and (_19486_, _14657_, _26242_);
  and (_19487_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_10186_, _19487_, _19486_);
  and (_19488_, _19039_, _26242_);
  and (_19489_, _19041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_10188_, _19489_, _19488_);
  and (_19490_, _01604_, _25927_);
  and (_19491_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_10195_, _19491_, _19490_);
  and (_19492_, _14657_, _26185_);
  and (_19493_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or (_10197_, _19493_, _19492_);
  and (_19494_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_19495_, _23550_, _23238_);
  and (_19496_, _23652_, _23601_);
  or (_19497_, _19496_, _19495_);
  and (_19498_, _19497_, _19494_);
  not (_19499_, _19494_);
  or (_19500_, _19499_, _23711_);
  and (_19501_, _19500_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_19502_, _19501_, _25630_);
  or (_19503_, _19502_, _19498_);
  or (_19504_, _26524_, _00644_);
  nand (_19505_, _19504_, _25630_);
  or (_19506_, _19505_, _00244_);
  and (_19507_, _19506_, _19503_);
  or (_19508_, _19507_, _25135_);
  nand (_19509_, _25135_, _25332_);
  and (_19510_, _19509_, _23049_);
  and (_10199_, _19510_, _19508_);
  and (_19511_, _19031_, _23768_);
  and (_19512_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_27310_, _19512_, _19511_);
  and (_19513_, _18676_, _26185_);
  and (_19514_, _18678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_10211_, _19514_, _19513_);
  and (_19515_, _01604_, _26185_);
  and (_19516_, _01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_10217_, _19516_, _19515_);
  and (_19517_, _19031_, _26170_);
  and (_19518_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_10219_, _19518_, _19517_);
  and (_19519_, _01568_, _26185_);
  and (_19520_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_10223_, _19520_, _19519_);
  and (_19521_, _14657_, _26085_);
  and (_19522_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or (_10224_, _19522_, _19521_);
  and (_19523_, _04139_, _26242_);
  and (_19524_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_10227_, _19524_, _19523_);
  and (_19525_, _01568_, _25886_);
  and (_19526_, _01570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_10228_, _19526_, _19525_);
  and (_19527_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  and (_19528_, _09103_, _25886_);
  or (_10230_, _19528_, _19527_);
  or (_19529_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_19530_, _23656_, _23604_);
  not (_19531_, _23656_);
  and (_19532_, _23659_, _19531_);
  or (_19533_, _19532_, _19530_);
  and (_19534_, _19533_, _23601_);
  nand (_19535_, _23590_, _23291_);
  and (_19536_, _23592_, _23238_);
  and (_19537_, _19536_, _19535_);
  and (_19538_, _23354_, _23607_);
  and (_19539_, _19538_, _24666_);
  and (_19540_, _19539_, _25778_);
  nand (_19541_, _19540_, _23752_);
  nand (_19542_, _19541_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_19543_, _19542_, _19537_);
  nor (_19544_, _19543_, _19534_);
  nand (_19545_, _19544_, _00804_);
  or (_19546_, _00530_, _00483_);
  or (_19547_, _19546_, _00575_);
  or (_19548_, _19547_, _00638_);
  or (_19549_, _00743_, _00688_);
  or (_19550_, _19549_, _19548_);
  and (_19551_, _19550_, _24794_);
  nor (_19552_, _19551_, _19545_);
  nand (_19553_, _19552_, _24993_);
  and (_19554_, _19553_, _19529_);
  or (_19555_, _19554_, _25630_);
  and (_19556_, _25895_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_19557_, _19556_, _25896_);
  nand (_19558_, _19557_, _25630_);
  and (_19559_, _19558_, _19555_);
  or (_19560_, _19559_, _25135_);
  or (_19561_, _25136_, _25258_);
  and (_19562_, _19561_, _23049_);
  and (_10232_, _19562_, _19560_);
  and (_19563_, _19031_, _25886_);
  and (_19564_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_10234_, _19564_, _19563_);
  and (_19565_, _02512_, _23830_);
  and (_19566_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_10239_, _19566_, _19565_);
  and (_19567_, _18650_, _25927_);
  and (_19568_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_27294_, _19568_, _19567_);
  and (_19569_, _19031_, _23830_);
  and (_19570_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_10247_, _19570_, _19569_);
  and (_19571_, _18650_, _25886_);
  and (_19572_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_10249_, _19572_, _19571_);
  and (_19573_, _26473_, _25630_);
  nand (_19574_, _19573_, _23729_);
  or (_19575_, _19573_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_19576_, _19575_, _25136_);
  and (_19577_, _19576_, _19574_);
  or (_19578_, _19577_, _25161_);
  and (_10253_, _19578_, _23049_);
  and (_19579_, _25630_, _26136_);
  nand (_19580_, _19579_, _23729_);
  or (_19581_, _19579_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_19582_, _19581_, _25136_);
  and (_19583_, _19582_, _19580_);
  nor (_19584_, _25136_, _25362_);
  or (_19585_, _19584_, _19583_);
  and (_10261_, _19585_, _23049_);
  and (_19586_, _19031_, _26085_);
  and (_19587_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_10263_, _19587_, _19586_);
  and (_19588_, _18650_, _23830_);
  and (_19589_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_10269_, _19589_, _19588_);
  and (_19590_, _14665_, _23768_);
  and (_19591_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_10277_, _19591_, _19590_);
  and (_19592_, _19031_, _26185_);
  and (_19593_, _19033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_10280_, _19593_, _19592_);
  and (_19594_, _18650_, _26085_);
  and (_19595_, _18652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_27295_, _19595_, _19594_);
  and (_19596_, _26301_, _26170_);
  and (_19597_, _26303_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_10292_, _19597_, _19596_);
  and (_19598_, _19025_, _25886_);
  and (_19599_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_10294_, _19599_, _19598_);
  and (_19600_, _10475_, _25886_);
  and (_19601_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_10300_, _19601_, _19600_);
  and (_19602_, _14665_, _25927_);
  and (_19603_, _14667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_10302_, _19603_, _19602_);
  and (_19604_, _04202_, _26170_);
  and (_19605_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_10310_, _19605_, _19604_);
  and (_19606_, _18638_, _25927_);
  and (_19607_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_10317_, _19607_, _19606_);
  and (_19608_, _10475_, _25927_);
  and (_19609_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_10319_, _19609_, _19608_);
  and (_19610_, _18772_, _26085_);
  and (_19611_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_10322_, _19611_, _19610_);
  and (_19612_, _26341_, _23768_);
  and (_19613_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_10323_, _19613_, _19612_);
  and (_19614_, _19025_, _23830_);
  and (_19615_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_27313_, _19615_, _19614_);
  and (_19616_, _18638_, _26170_);
  and (_19617_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_10332_, _19617_, _19616_);
  and (_10334_, _03216_, _23049_);
  and (_19618_, _10475_, _26185_);
  and (_19619_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_10339_, _19619_, _19618_);
  and (_19620_, _04202_, _25927_);
  and (_19621_, _04204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_10341_, _19621_, _19620_);
  and (_19622_, _18638_, _23830_);
  and (_19623_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_10343_, _19623_, _19622_);
  and (_19624_, _26341_, _26185_);
  and (_19625_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_10345_, _19625_, _19624_);
  and (_19626_, _19025_, _26185_);
  and (_19627_, _19027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_10346_, _19627_, _19626_);
  and (_19628_, _26341_, _25886_);
  and (_19629_, _26345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_10349_, _19629_, _19628_);
  and (_19630_, _25630_, _26130_);
  nand (_19631_, _19630_, _23729_);
  or (_19632_, _19630_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_19633_, _19632_, _25136_);
  and (_19634_, _19633_, _19631_);
  or (_19635_, _19634_, _25138_);
  and (_10350_, _19635_, _23049_);
  and (_19636_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_19637_, _09450_, _23830_);
  or (_10353_, _19637_, _19636_);
  and (_19638_, _18638_, _26085_);
  and (_19639_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_10356_, _19639_, _19638_);
  and (_19640_, _18990_, _26170_);
  and (_19641_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_10359_, _19641_, _19640_);
  and (_19642_, _14657_, _25927_);
  and (_19643_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_10362_, _19643_, _19642_);
  and (_19644_, _25630_, _25224_);
  nand (_19645_, _19644_, _23729_);
  or (_19646_, _19644_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_19647_, _19646_, _25136_);
  and (_19648_, _19647_, _19645_);
  nor (_19649_, _25136_, _25279_);
  or (_19650_, _19649_, _19648_);
  and (_10364_, _19650_, _23049_);
  and (_19651_, _18638_, _26185_);
  and (_19652_, _18640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_10367_, _19652_, _19651_);
  and (_19653_, _26072_, _25938_);
  and (_19654_, _19653_, _26242_);
  not (_19655_, _19653_);
  and (_19656_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_10373_, _19656_, _19654_);
  and (_19657_, _18990_, _25886_);
  and (_19658_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_10374_, _19658_, _19657_);
  and (_19659_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  and (_19660_, _09103_, _26085_);
  or (_10376_, _19660_, _19659_);
  and (_19661_, _19653_, _23830_);
  and (_19662_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_10379_, _19662_, _19661_);
  and (_19663_, _09104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  and (_19664_, _09103_, _26242_);
  or (_10381_, _19664_, _19663_);
  and (_19665_, _18632_, _25927_);
  and (_19666_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_10407_, _19666_, _19665_);
  and (_19667_, _18990_, _26085_);
  and (_19668_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_10413_, _19668_, _19667_);
  and (_19669_, _14657_, _23768_);
  and (_19670_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or (_10421_, _19670_, _19669_);
  and (_19671_, _18990_, _26242_);
  and (_19672_, _18992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_10444_, _19672_, _19671_);
  and (_19673_, _18632_, _26170_);
  and (_19674_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_27297_, _19674_, _19673_);
  nor (_10449_, _03260_, rst);
  and (_19675_, _18704_, _26170_);
  and (_19676_, _18706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_10467_, _19676_, _19675_);
  and (_19677_, _14398_, _26242_);
  and (_19678_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_10470_, _19678_, _19677_);
  and (_19679_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_19680_, _09087_, _25927_);
  or (_10484_, _19680_, _19679_);
  and (_19681_, _18980_, _26242_);
  and (_19682_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_10490_, _19682_, _19681_);
  and (_19683_, _18984_, _25927_);
  and (_19684_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_10491_, _19684_, _19683_);
  and (_10496_, _03201_, _23049_);
  and (_10498_, _03234_, _23049_);
  and (_19685_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_19686_, _09087_, _25886_);
  or (_10500_, _19686_, _19685_);
  and (_19687_, _17822_, _25927_);
  and (_19688_, _17824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or (_10512_, _19688_, _19687_);
  and (_10519_, _03187_, _23049_);
  and (_10520_, _03246_, _23049_);
  and (_19689_, _18632_, _25886_);
  and (_19690_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_10523_, _19690_, _19689_);
  and (_19691_, _18632_, _26085_);
  and (_19692_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_10526_, _19692_, _19691_);
  and (_19693_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_19694_, _09450_, _25886_);
  or (_10527_, _19694_, _19693_);
  and (_10536_, _03174_, _23049_);
  and (_10537_, _03270_, _23049_);
  and (_19695_, _18984_, _26170_);
  and (_19696_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_10546_, _19696_, _19695_);
  and (_19697_, _04139_, _25886_);
  and (_19698_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or (_27186_, _19698_, _19697_);
  and (_19699_, _18632_, _26242_);
  and (_19700_, _18634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_10555_, _19700_, _19699_);
  and (_19701_, _16208_, _26185_);
  and (_19702_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_10557_, _19702_, _19701_);
  and (_19703_, _14731_, _26242_);
  and (_19704_, _14733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_27250_, _19704_, _19703_);
  and (_19705_, _18984_, _23830_);
  and (_19706_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_10560_, _19706_, _19705_);
  and (_19707_, _18980_, _26170_);
  and (_19709_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_10563_, _19709_, _19707_);
  and (_19710_, _18984_, _26185_);
  and (_19711_, _18986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_10572_, _19711_, _19710_);
  and (_19712_, _18628_, _23768_);
  and (_19713_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_10574_, _19713_, _19712_);
  and (_19714_, _09451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_19715_, _09450_, _26170_);
  or (_10576_, _19715_, _19714_);
  and (_19716_, _18980_, _25927_);
  and (_19717_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_10580_, _19717_, _19716_);
  and (_19718_, _18956_, _23768_);
  and (_19719_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_10587_, _19719_, _19718_);
  and (_19720_, _18980_, _23768_);
  and (_19721_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_10590_, _19721_, _19720_);
  and (_19722_, _05551_, _26185_);
  and (_19723_, _05553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_10593_, _19723_, _19722_);
  and (_19724_, _18628_, _26170_);
  and (_19725_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_10601_, _19725_, _19724_);
  and (_19726_, _18628_, _23830_);
  and (_19727_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_10604_, _19727_, _19726_);
  and (_19728_, _18956_, _25927_);
  and (_19730_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_10606_, _19730_, _19728_);
  and (_19731_, _18628_, _26185_);
  and (_19732_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_10611_, _19732_, _19731_);
  and (_19733_, _18956_, _25886_);
  and (_19734_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_10620_, _19734_, _19733_);
  and (_19735_, _18956_, _26085_);
  and (_19736_, _18958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_27318_, _19736_, _19735_);
  and (_19737_, _26329_, _26085_);
  and (_19738_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_10626_, _19738_, _19737_);
  and (_19739_, _18628_, _26242_);
  and (_19740_, _18630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_10628_, _19740_, _19739_);
  and (_19741_, _26329_, _25886_);
  and (_19742_, _26332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_10631_, _19742_, _19741_);
  and (_19743_, _17846_, _26170_);
  and (_19744_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_10636_, _19744_, _19743_);
  and (_19745_, _18950_, _25927_);
  and (_19746_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_10639_, _19746_, _19745_);
  and (_19747_, _16208_, _25886_);
  and (_19748_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_10642_, _19748_, _19747_);
  and (_19749_, _17846_, _25886_);
  and (_19751_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_10648_, _19751_, _19749_);
  nor (_26893_[2], _23063_, rst);
  and (_19752_, _14991_, _26242_);
  and (_19753_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_10654_, _19753_, _19752_);
  and (_19754_, _18772_, _25927_);
  and (_19755_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_10656_, _19755_, _19754_);
  and (_19756_, _18950_, _26170_);
  and (_19757_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_10658_, _19757_, _19756_);
  and (_19758_, _17846_, _26085_);
  and (_19759_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_10659_, _19759_, _19758_);
  and (_19760_, _16208_, _26085_);
  and (_19761_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_27265_, _19761_, _19760_);
  and (_19762_, _00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  and (_19763_, _00089_, _23830_);
  or (_10665_, _19763_, _19762_);
  and (_19764_, _18950_, _23830_);
  and (_19765_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_10669_, _19765_, _19764_);
  and (_19766_, _17846_, _26242_);
  and (_19767_, _17848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_10671_, _19767_, _19766_);
  and (_19768_, _26294_, _26242_);
  and (_19769_, _26296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_10674_, _19769_, _19768_);
  and (_19770_, _01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_19771_, _01608_, _25927_);
  or (_10678_, _19771_, _19770_);
  and (_19772_, _15146_, _25927_);
  and (_19773_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_10679_, _19773_, _19772_);
  and (_19774_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  and (_19775_, _04148_, _23768_);
  or (_10684_, _19775_, _19774_);
  and (_19776_, _14657_, _25886_);
  and (_19777_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_10687_, _19777_, _19776_);
  and (_19778_, _17840_, _25927_);
  and (_19779_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_10692_, _19779_, _19778_);
  and (_19780_, _04139_, _26170_);
  and (_19781_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or (_10694_, _19781_, _19780_);
  and (_19782_, _18950_, _26085_);
  and (_19783_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_10696_, _19783_, _19782_);
  or (_19785_, _22968_, _00137_);
  or (_19786_, _22738_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_19787_, _19786_, _23049_);
  and (_26896_[4], _19787_, _19785_);
  and (_19788_, _14906_, _23830_);
  and (_19789_, _14908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_10701_, _19789_, _19788_);
  and (_19790_, _09053_, _26085_);
  and (_19791_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_10708_, _19791_, _19790_);
  and (_19792_, _18950_, _26185_);
  and (_19793_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_10709_, _19793_, _19792_);
  and (_19794_, _17840_, _26170_);
  and (_19795_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_10712_, _19795_, _19794_);
  and (_19796_, _14657_, _26170_);
  and (_19797_, _14659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or (_10713_, _19797_, _19796_);
  and (_19798_, _09053_, _26170_);
  and (_19799_, _09056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_10716_, _19799_, _19798_);
  and (_19800_, _05755_, _23830_);
  and (_19801_, _05758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_10718_, _19801_, _19800_);
  and (_19802_, _25886_, _23231_);
  and (_19803_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_27232_, _19803_, _19802_);
  and (_19804_, _18950_, _26242_);
  and (_19805_, _18952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_10720_, _19805_, _19804_);
  and (_19806_, _17840_, _23830_);
  and (_19807_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_10723_, _19807_, _19806_);
  and (_19808_, _18980_, _23830_);
  and (_19809_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_10727_, _19809_, _19808_);
  and (_19810_, _17840_, _26185_);
  and (_19811_, _17842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_10729_, _19811_, _19810_);
  and (_19812_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  and (_19813_, _10218_, _26170_);
  or (_10730_, _19813_, _19812_);
  and (_19814_, _03115_, _25886_);
  and (_19815_, _03117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_10733_, _19815_, _19814_);
  and (_19816_, _18909_, _23768_);
  and (_19817_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_10735_, _19817_, _19816_);
  and (_19818_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  and (_19819_, _10218_, _25927_);
  or (_10737_, _19819_, _19818_);
  and (_19820_, _18909_, _25886_);
  and (_19821_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_10741_, _19821_, _19820_);
  and (_19822_, _17834_, _23768_);
  and (_19823_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_10744_, _19823_, _19822_);
  and (_19824_, _18980_, _25886_);
  and (_19826_, _18982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_10747_, _19826_, _19824_);
  nor (_19827_, _00404_, _03204_);
  nand (_19828_, _19827_, _23729_);
  or (_19829_, _19827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_19830_, _19829_, _25618_);
  and (_19831_, _19830_, _19828_);
  nand (_19832_, _00410_, _25417_);
  or (_19833_, _00410_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_19834_, _19833_, _25128_);
  and (_19835_, _19834_, _19832_);
  and (_19836_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_19837_, _19836_, rst);
  or (_19838_, _19837_, _19835_);
  or (_10749_, _19838_, _19831_);
  and (_19839_, _18909_, _23830_);
  and (_19840_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_10753_, _19840_, _19839_);
  and (_19841_, _17834_, _25927_);
  and (_19842_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_10755_, _19842_, _19841_);
  nand (_19843_, _24809_, _24794_);
  or (_19844_, _24794_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_19845_, _19844_, _23049_);
  and (_10757_, _19845_, _19843_);
  and (_19846_, _17834_, _25886_);
  and (_19847_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_10758_, _19847_, _19846_);
  and (_19848_, _18909_, _26185_);
  and (_19849_, _18911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_10764_, _19849_, _19848_);
  and (_19850_, _19653_, _23768_);
  and (_19851_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_10771_, _19851_, _19850_);
  and (_19852_, _26351_, _26085_);
  and (_19853_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_10773_, _19853_, _19852_);
  and (_19854_, _17834_, _23830_);
  and (_19855_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_10774_, _19855_, _19854_);
  and (_19856_, _17834_, _26242_);
  and (_19857_, _17836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_10778_, _19857_, _19856_);
  and (_19858_, _18864_, _25927_);
  and (_19859_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_10781_, _19859_, _19858_);
  and (_19860_, _18864_, _25886_);
  and (_19861_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_10792_, _19861_, _19860_);
  and (_19862_, _15050_, _23830_);
  and (_19863_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_10796_, _19863_, _19862_);
  and (_19864_, _15050_, _26185_);
  and (_19865_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_10799_, _19865_, _19864_);
  and (_19866_, _18864_, _23830_);
  and (_19867_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_10801_, _19867_, _19866_);
  and (_19868_, _17830_, _23768_);
  and (_19869_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_10803_, _19869_, _19868_);
  and (_19870_, _15146_, _25886_);
  and (_19871_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_10805_, _19871_, _19870_);
  and (_19872_, _18864_, _26185_);
  and (_19873_, _18866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_10809_, _19873_, _19872_);
  and (_19874_, _14398_, _25886_);
  and (_19875_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or (_10811_, _19875_, _19874_);
  and (_19876_, _17830_, _26170_);
  and (_19877_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_10813_, _19877_, _19876_);
  nand (_19878_, _02406_, _25417_);
  or (_19879_, _02406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_19880_, _19879_, _23049_);
  and (_10817_, _19880_, _19878_);
  nor (_19881_, _01574_, _03204_);
  nand (_19882_, _19881_, _23729_);
  or (_19883_, _19881_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_19884_, _19883_, _25618_);
  and (_19885_, _19884_, _19882_);
  nand (_19886_, _01578_, _25417_);
  or (_19887_, _01578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_19888_, _19887_, _25128_);
  and (_19889_, _19888_, _19886_);
  and (_19890_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_19891_, _19890_, rst);
  or (_19892_, _19891_, _19889_);
  or (_10819_, _19892_, _19885_);
  and (_19893_, _00016_, _25886_);
  and (_19894_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_10821_, _19894_, _19893_);
  and (_19895_, _00016_, _23768_);
  and (_19896_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_10824_, _19896_, _19895_);
  and (_19897_, _15081_, _25927_);
  and (_19898_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_10829_, _19898_, _19897_);
  and (_19899_, _15081_, _26170_);
  and (_19900_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_10831_, _19900_, _19899_);
  and (_19901_, _15081_, _23830_);
  and (_19902_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_10843_, _19902_, _19901_);
  and (_19903_, _14398_, _26170_);
  and (_19904_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_10845_, _19904_, _19903_);
  and (_19905_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_19906_, _09087_, _26085_);
  or (_10847_, _19906_, _19905_);
  and (_19907_, _04139_, _26085_);
  and (_19908_, _04141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or (_10854_, _19908_, _19907_);
  and (_19909_, _09089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_19910_, _09087_, _26185_);
  or (_10866_, _19910_, _19909_);
  and (_19911_, _14629_, _23768_);
  and (_19912_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_10871_, _19912_, _19911_);
  and (_19913_, _15081_, _26085_);
  and (_19914_, _15084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_10874_, _19914_, _19913_);
  and (_19915_, _26170_, _23849_);
  and (_19916_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_27263_, _19916_, _19915_);
  and (_19917_, _26446_, _25886_);
  and (_19918_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_10880_, _19918_, _19917_);
  and (_19919_, _25536_, _01826_);
  nand (_19920_, _19919_, _23729_);
  or (_19921_, _19919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19922_, _19921_, _25618_);
  and (_19923_, _19922_, _19920_);
  nand (_19924_, _01834_, _25417_);
  or (_19925_, _01834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_19926_, _19925_, _25128_);
  and (_19927_, _19926_, _19924_);
  and (_19928_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_19929_, _19928_, rst);
  or (_19930_, _19929_, _19927_);
  or (_10889_, _19930_, _19923_);
  and (_19931_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_19932_, _09047_, _23768_);
  or (_10892_, _19932_, _19931_);
  and (_19933_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_19934_, _09047_, _26170_);
  or (_10894_, _19934_, _19933_);
  and (_19935_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_19936_, _09047_, _23830_);
  or (_27161_, _19936_, _19935_);
  and (_19937_, _26446_, _23830_);
  and (_19938_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_10900_, _19938_, _19937_);
  and (_19939_, _26446_, _26085_);
  and (_19940_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_10903_, _19940_, _19939_);
  and (_19941_, _26446_, _26242_);
  and (_19942_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_10908_, _19942_, _19941_);
  and (_19943_, _15064_, _25927_);
  and (_19944_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_10915_, _19944_, _19943_);
  and (_19945_, _09049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_19946_, _09047_, _26085_);
  or (_10917_, _19946_, _19945_);
  and (_19947_, _18772_, _23768_);
  and (_19948_, _18774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_10920_, _19948_, _19947_);
  and (_19949_, _00251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_19950_, _03204_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_19951_, _19950_, _03206_);
  and (_19952_, _19951_, _00249_);
  or (_19953_, _19952_, _19949_);
  and (_19954_, _19953_, _25618_);
  nand (_19955_, _00257_, _25417_);
  or (_19956_, _00257_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_19957_, _19956_, _25128_);
  and (_19958_, _19957_, _19955_);
  and (_19959_, _25751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_19960_, _19959_, rst);
  or (_19961_, _19960_, _19958_);
  or (_10922_, _19961_, _19954_);
  and (_19962_, _15064_, _26170_);
  and (_19963_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_26949_, _19963_, _19962_);
  and (_19964_, _14398_, _26085_);
  and (_19965_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_10928_, _19965_, _19964_);
  and (_19966_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_19967_, _04105_, _25927_);
  or (_10931_, _19967_, _19966_);
  and (_19968_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  and (_19969_, _04148_, _26170_);
  or (_10934_, _19969_, _19968_);
  and (_19970_, _16208_, _26242_);
  and (_19971_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_10941_, _19971_, _19970_);
  and (_19972_, _14398_, _23830_);
  and (_19973_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or (_26997_, _19973_, _19972_);
  and (_19974_, _15064_, _23830_);
  and (_19975_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_10945_, _19975_, _19974_);
  and (_19976_, _09418_, _26170_);
  and (_19977_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_27109_, _19977_, _19976_);
  and (_19978_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_19979_, _04105_, _23768_);
  or (_10955_, _19979_, _19978_);
  and (_19980_, _09418_, _25927_);
  and (_19981_, _09420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_10957_, _19981_, _19980_);
  and (_19982_, _26085_, _23849_);
  and (_19983_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_10973_, _19983_, _19982_);
  and (_19984_, _01371_, _23830_);
  and (_19985_, _01373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_10976_, _19985_, _19984_);
  and (_19986_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  and (_19987_, _10218_, _23768_);
  or (_10979_, _19987_, _19986_);
  and (_19988_, _14404_, _26085_);
  and (_19989_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_26996_, _19989_, _19988_);
  and (_19990_, _26370_, _26085_);
  and (_19991_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_10982_, _19991_, _19990_);
  and (_19992_, _26356_, _26085_);
  and (_19993_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_10984_, _19993_, _19992_);
  and (_19994_, _26376_, _26170_);
  and (_19995_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_10989_, _19995_, _19994_);
  and (_19996_, _26442_, _26242_);
  and (_19997_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_10992_, _19997_, _19996_);
  and (_19998_, _25891_, _25131_);
  nand (_19999_, _19998_, _23729_);
  or (_20000_, _19998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_20001_, _20000_, _25910_);
  and (_20002_, _20001_, _19999_);
  and (_20003_, _25903_, _25283_);
  or (_20004_, _20003_, _20002_);
  and (_10997_, _20004_, _23049_);
  and (_20005_, _26442_, _26085_);
  and (_20006_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_27322_, _20006_, _20005_);
  and (_20007_, _15064_, _26085_);
  and (_20008_, _15066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_11002_, _20008_, _20007_);
  and (_20009_, _26366_, _26185_);
  and (_20010_, _26368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_11004_, _20010_, _20009_);
  and (_20011_, _26376_, _25927_);
  and (_20012_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_11006_, _20012_, _20011_);
  and (_20013_, _26376_, _25886_);
  and (_20014_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_11009_, _20014_, _20013_);
  and (_20015_, _26442_, _26185_);
  and (_20016_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_11011_, _20016_, _20015_);
  and (_20017_, _15054_, _25927_);
  and (_20018_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_11013_, _20018_, _20017_);
  and (_20019_, _26356_, _25927_);
  and (_20020_, _26359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_11015_, _20020_, _20019_);
  and (_20021_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  and (_20022_, _04148_, _25927_);
  or (_27178_, _20022_, _20021_);
  and (_20023_, _26428_, _25927_);
  and (_20024_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_27323_, _20024_, _20023_);
  and (_20025_, _16208_, _23768_);
  and (_20026_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_11024_, _20026_, _20025_);
  and (_20027_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_20028_, _26096_, _14829_);
  and (_20029_, _20028_, _26120_);
  and (_20030_, _26117_, _26104_);
  nor (_20031_, _20030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_20032_, _20031_, _05618_);
  or (_20033_, _20032_, _26093_);
  or (_20034_, _20033_, _20029_);
  nand (_20035_, _26093_, _14829_);
  and (_20036_, _20035_, _05563_);
  and (_20037_, _20036_, _20034_);
  or (_20038_, _20037_, _20027_);
  nor (_20039_, _26142_, _25332_);
  or (_20040_, _20039_, _20038_);
  and (_11027_, _20040_, _23049_);
  and (_20041_, _26428_, _25886_);
  and (_20042_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_11029_, _20042_, _20041_);
  and (_20043_, _15054_, _26170_);
  and (_20044_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_26950_, _20044_, _20043_);
  and (_20045_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_20046_, _04105_, _26085_);
  or (_27177_, _20046_, _20045_);
  and (_20047_, _26596_, _26242_);
  and (_20048_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_11033_, _20048_, _20047_);
  and (_20049_, _26458_, _26185_);
  and (_20050_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_11035_, _20050_, _20049_);
  nor (_20051_, _26096_, _14822_);
  and (_20052_, _20051_, _26120_);
  not (_20053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand (_20054_, _26116_, _26104_);
  and (_20055_, _20054_, _20053_);
  nor (_20056_, _20055_, _20030_);
  or (_20057_, _20056_, _26093_);
  or (_20058_, _20057_, _20052_);
  nand (_20059_, _26093_, _14822_);
  and (_20060_, _20059_, _05563_);
  and (_20061_, _20060_, _20058_);
  and (_20062_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_20063_, _20062_, _20061_);
  nor (_20064_, _26142_, _25362_);
  or (_20065_, _20064_, _20063_);
  and (_11037_, _20065_, _23049_);
  and (_20066_, _26376_, _26185_);
  and (_20067_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_11039_, _20067_, _20066_);
  nor (_20068_, _23215_, _23153_);
  and (_20069_, _20068_, _25182_);
  and (_20070_, _20069_, _25900_);
  and (_20071_, _20070_, _25128_);
  not (_20072_, _20071_);
  and (_20073_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_20074_, _20073_, _26120_);
  and (_20075_, _26115_, _26104_);
  or (_20076_, _20075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_20077_, _20076_, _20054_);
  or (_20078_, _20077_, _26093_);
  or (_20079_, _20078_, _20074_);
  nor (_20080_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_20081_, _20080_, _26132_);
  and (_20082_, _20081_, _20079_);
  and (_20083_, _20068_, _25130_);
  and (_20084_, _20083_, _25900_);
  and (_20085_, _20084_, _25128_);
  and (_20086_, _20085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_20087_, _20086_, _20082_);
  and (_20088_, _20087_, _20072_);
  nor (_20089_, _20072_, _23824_);
  or (_20090_, _20089_, _20088_);
  and (_11041_, _20090_, _23049_);
  and (_20091_, _26370_, _25927_);
  and (_20092_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_11046_, _20092_, _20091_);
  and (_20093_, _26370_, _25886_);
  and (_20094_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_11048_, _20094_, _20093_);
  and (_20095_, _15054_, _25886_);
  and (_20096_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_26951_, _20096_, _20095_);
  or (_20097_, _15280_, _01875_);
  or (_20098_, _20097_, _15254_);
  and (_20099_, _20098_, _22739_);
  and (_20100_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_20101_, _20100_, _15299_);
  or (_20102_, _20101_, _20099_);
  and (_26898_[1], _20102_, _23049_);
  and (_20103_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_20104_, _04105_, _23830_);
  or (_11052_, _20104_, _20103_);
  and (_20105_, _26370_, _23768_);
  and (_20106_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_11055_, _20106_, _20105_);
  and (_20107_, _26376_, _26085_);
  and (_20108_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_11057_, _20108_, _20107_);
  and (_20109_, _04106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_20110_, _04105_, _25886_);
  or (_11061_, _20110_, _20109_);
  and (_20111_, _26596_, _25886_);
  and (_20112_, _26598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_11063_, _20112_, _20111_);
  and (_20113_, _26370_, _26170_);
  and (_20114_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_11066_, _20114_, _20113_);
  and (_20115_, _14398_, _23768_);
  and (_20116_, _14400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_11068_, _20116_, _20115_);
  and (_20117_, _26376_, _26242_);
  and (_20118_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_27307_, _20118_, _20117_);
  and (_20119_, _26458_, _26085_);
  and (_20120_, _26460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_27292_, _20120_, _20119_);
  and (_20121_, _15054_, _26085_);
  and (_20122_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_11073_, _20122_, _20121_);
  and (_20123_, _15054_, _26242_);
  and (_20124_, _15056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_26952_, _20124_, _20123_);
  and (_20125_, _14404_, _26242_);
  and (_20126_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_11078_, _20126_, _20125_);
  and (_20127_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_20128_, _20127_, _26120_);
  and (_20129_, _26113_, _26104_);
  or (_20130_, _20129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_20131_, _20130_, _09373_);
  or (_20132_, _20131_, _26093_);
  or (_20133_, _20132_, _20128_);
  nor (_20134_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_20135_, _20134_, _26132_);
  and (_20136_, _20135_, _20133_);
  and (_20137_, _20085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_20138_, _20137_, _20136_);
  and (_20139_, _20138_, _20072_);
  and (_20140_, _20071_, _25258_);
  or (_20141_, _20140_, _20139_);
  and (_11081_, _20141_, _23049_);
  and (_20142_, _26097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_20143_, _20142_, _26120_);
  and (_20144_, _26112_, _26104_);
  nor (_20145_, _20144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_20146_, _20145_, _20129_);
  or (_20147_, _20146_, _26093_);
  or (_20148_, _20147_, _20143_);
  nor (_20149_, _26095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_20150_, _20149_, _09072_);
  and (_20151_, _20150_, _20148_);
  and (_20152_, _26132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_20153_, _26142_, _25279_);
  or (_20154_, _20153_, _20152_);
  or (_20155_, _20154_, _20151_);
  and (_11083_, _20155_, _23049_);
  and (_20156_, _26242_, _23849_);
  and (_20157_, _23851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_11086_, _20157_, _20156_);
  and (_20158_, _26446_, _23768_);
  and (_20159_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_11090_, _20159_, _20158_);
  and (_20160_, _26428_, _26242_);
  and (_20161_, _26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_11092_, _20161_, _20160_);
  and (_20162_, _26446_, _26170_);
  and (_20163_, _26448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_11094_, _20163_, _20162_);
  and (_20164_, _15050_, _23768_);
  and (_20165_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_11096_, _20165_, _20164_);
  and (_20166_, _26085_, _23231_);
  and (_20167_, _23770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_11098_, _20167_, _20166_);
  nor (_20168_, _26133_, _25362_);
  nor (_20169_, _26096_, _09685_);
  nand (_20170_, _20169_, _26120_);
  and (_20171_, _26108_, _26104_);
  nor (_20172_, _20171_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_20173_, _20172_, _09353_);
  and (_20174_, _20173_, _26095_);
  nand (_20175_, _20174_, _20170_);
  and (_20176_, _26093_, _09685_);
  nor (_20177_, _20176_, _09072_);
  and (_20178_, _20177_, _20175_);
  and (_20179_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_20180_, _20179_, _20178_);
  or (_20181_, _20180_, _20168_);
  and (_11100_, _20181_, _23049_);
  and (_20182_, _26783_, _26170_);
  and (_20183_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_27282_, _20183_, _20182_);
  and (_20184_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_20185_, _09304_, _25886_);
  or (_27080_, _20185_, _20184_);
  nor (_20186_, _26133_, _23824_);
  nor (_20187_, _26096_, _14920_);
  nand (_20188_, _20187_, _26120_);
  and (_20189_, _26107_, _26104_);
  nor (_20190_, _20189_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_20191_, _20190_, _20171_);
  and (_20192_, _20191_, _26095_);
  nand (_20193_, _20192_, _20188_);
  and (_20194_, _26093_, _14920_);
  nor (_20195_, _20194_, _09072_);
  and (_20196_, _20195_, _20193_);
  and (_20197_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_20198_, _20197_, _20196_);
  or (_20199_, _20198_, _20186_);
  and (_11104_, _20199_, _23049_);
  and (_20200_, _00038_, _26242_);
  and (_20201_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_27287_, _20201_, _20200_);
  nor (_20202_, _26096_, _14930_);
  nand (_20203_, _20202_, _26120_);
  not (_20204_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_20205_, _26124_, _20204_);
  or (_20206_, _20205_, _20189_);
  and (_20207_, _20206_, _26095_);
  nand (_20208_, _20207_, _20203_);
  and (_20209_, _26093_, _14930_);
  nor (_20210_, _20209_, _09072_);
  and (_20211_, _20210_, _20208_);
  and (_20212_, _26138_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_20213_, _26133_, _25160_);
  or (_20214_, _20213_, _20212_);
  or (_20215_, _20214_, _20211_);
  and (_11108_, _20215_, _23049_);
  and (_20216_, _00038_, _25927_);
  and (_20217_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_27285_, _20217_, _20216_);
  and (_20218_, _15050_, _26170_);
  and (_20219_, _15052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_26953_, _20219_, _20218_);
  and (_20220_, _17830_, _26085_);
  and (_20221_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_27305_, _20221_, _20220_);
  and (_20222_, _26376_, _23768_);
  and (_20223_, _26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_11115_, _20223_, _20222_);
  and (_20224_, _17830_, _26242_);
  and (_20225_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_27306_, _20225_, _20224_);
  and (_20226_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  and (_20227_, _04143_, _23768_);
  or (_11121_, _20227_, _20226_);
  and (_20228_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_20229_, _04113_, _26170_);
  or (_27175_, _20229_, _20228_);
  and (_20230_, _26442_, _23768_);
  and (_20231_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_11124_, _20231_, _20230_);
  and (_20232_, _26442_, _26170_);
  and (_20233_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_11126_, _20233_, _20232_);
  and (_20234_, _26442_, _25886_);
  and (_20235_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_11128_, _20235_, _20234_);
  and (_20236_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_20237_, _04113_, _25886_);
  or (_11134_, _20237_, _20236_);
  and (_20238_, _00038_, _23830_);
  and (_20239_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_11137_, _20239_, _20238_);
  and (_20240_, _25891_, _26136_);
  nand (_20241_, _20240_, _23729_);
  or (_20242_, _20240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_20243_, _20242_, _25910_);
  and (_20244_, _20243_, _20241_);
  nor (_20245_, _25910_, _25362_);
  or (_20246_, _20245_, _20244_);
  and (_11139_, _20246_, _23049_);
  and (_20247_, _23215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_20248_, _20247_, _26557_);
  and (_20249_, _20248_, _25891_);
  not (_20250_, _25891_);
  or (_20251_, _26563_, _20250_);
  and (_20252_, _20251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_20253_, _20252_, _25903_);
  or (_20254_, _20253_, _20249_);
  nand (_20255_, _25903_, _23824_);
  and (_20256_, _20255_, _23049_);
  and (_11141_, _20256_, _20254_);
  nand (_20257_, _00071_, _25332_);
  or (_20258_, _09313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_20259_, _20258_, _09316_);
  and (_20260_, _00083_, _00072_);
  or (_20261_, _20260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_20262_, _20261_, _09318_);
  and (_20263_, _02497_, _00083_);
  or (_20264_, _20263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_20265_, _09321_, _02503_);
  and (_20266_, _20265_, _20264_);
  or (_20267_, _20266_, _20262_);
  or (_20268_, _20267_, _20259_);
  or (_20269_, _20268_, _00071_);
  and (_20270_, _20269_, _00070_);
  and (_20271_, _20270_, _20257_);
  and (_20272_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_20273_, _20272_, _20271_);
  and (_11145_, _20273_, _23049_);
  and (_20274_, _15044_, _23768_);
  and (_20275_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_26957_, _20275_, _20274_);
  and (_20276_, _26473_, _25891_);
  nand (_20277_, _20276_, _23729_);
  or (_20278_, _20276_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_20279_, _20278_, _25910_);
  and (_20280_, _20279_, _20277_);
  nor (_20281_, _25910_, _25160_);
  or (_20282_, _20281_, _20280_);
  and (_11152_, _20282_, _23049_);
  and (_20283_, _17830_, _23830_);
  and (_20284_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_27304_, _20284_, _20283_);
  and (_20285_, _00016_, _26242_);
  and (_20286_, _00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_27281_, _20286_, _20285_);
  and (_20287_, _26442_, _25927_);
  and (_20288_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_11157_, _20288_, _20287_);
  and (_20289_, _17830_, _26185_);
  and (_20290_, _17832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_11159_, _20290_, _20289_);
  and (_20291_, _00038_, _23768_);
  and (_20292_, _00041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_11161_, _20292_, _20291_);
  nand (_20293_, _00071_, _25362_);
  not (_20294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_20295_, _09311_, _00081_);
  and (_20296_, _20295_, _09309_);
  and (_20297_, _20296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_20298_, _20297_, _20294_);
  and (_20299_, _20297_, _20294_);
  or (_20300_, _20299_, _20298_);
  and (_20301_, _20300_, _01673_);
  and (_20302_, _00082_, _00072_);
  or (_20303_, _20302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_20304_, _20260_, _01674_);
  and (_20305_, _20304_, _20303_);
  and (_20306_, _02497_, _00082_);
  or (_20307_, _20306_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_20308_, _20263_, _02503_);
  and (_20309_, _20308_, _20307_);
  or (_20310_, _20309_, _20305_);
  or (_20311_, _20310_, _20301_);
  or (_20312_, _20311_, _00071_);
  and (_20313_, _20312_, _00070_);
  and (_20314_, _20313_, _20293_);
  and (_20315_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_20316_, _20315_, _20314_);
  and (_11163_, _20316_, _23049_);
  nand (_20317_, _00071_, _23824_);
  or (_20318_, _20296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_20319_, _20297_);
  and (_20320_, _20319_, _01673_);
  and (_20321_, _20320_, _20318_);
  and (_20322_, _00081_, _00072_);
  or (_20323_, _20322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_20324_, _20302_, _01674_);
  and (_20325_, _20324_, _20323_);
  not (_20326_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_20327_, _02497_, _00081_);
  nor (_20328_, _20327_, _20326_);
  and (_20329_, _20327_, _20326_);
  or (_20330_, _20329_, _20328_);
  and (_20331_, _20330_, _01664_);
  or (_20332_, _20331_, _20325_);
  or (_20333_, _20332_, _20321_);
  or (_20334_, _20333_, _00071_);
  and (_20335_, _20334_, _00070_);
  and (_20336_, _20335_, _20317_);
  and (_20337_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_20338_, _20337_, _20336_);
  and (_11165_, _20338_, _23049_);
  and (_20339_, _26783_, _26085_);
  and (_20340_, _26785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_11167_, _20340_, _20339_);
  and (_20341_, _14408_, _26242_);
  and (_20342_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_26995_, _20342_, _20341_);
  and (_20343_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_20344_, _09304_, _26170_);
  or (_11174_, _20344_, _20343_);
  and (_20345_, _15044_, _25927_);
  and (_20346_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_26958_, _20346_, _20345_);
  and (_20347_, _10299_, _01666_);
  or (_20348_, _20347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_20349_, _20347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_20350_, _20349_, _01673_);
  and (_20351_, _20350_, _20348_);
  and (_20352_, _00080_, _00072_);
  or (_20353_, _20352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_20354_, _20322_, _01674_);
  and (_20355_, _20354_, _20353_);
  and (_20356_, _02497_, _00080_);
  or (_20357_, _20356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_20358_, _20327_, _02503_);
  and (_20359_, _20358_, _20357_);
  or (_20360_, _20359_, _20355_);
  or (_20361_, _20360_, _20351_);
  or (_20362_, _20361_, _00071_);
  nand (_20363_, _00071_, _25160_);
  and (_20364_, _20363_, _20362_);
  or (_20365_, _20364_, _00069_);
  or (_20366_, _00070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_20367_, _20366_, _23049_);
  and (_11183_, _20367_, _20365_);
  and (_20368_, _15044_, _25886_);
  and (_20369_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_11186_, _20369_, _20368_);
  and (_20370_, _15044_, _26085_);
  and (_20371_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_11190_, _20371_, _20370_);
  and (_20372_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_20373_, _25091_, _22739_);
  or (_20374_, _20373_, _20372_);
  or (_20375_, _20374_, _15299_);
  and (_26900_[2], _20375_, _23049_);
  and (_20376_, _01367_, _23830_);
  and (_20377_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_11198_, _20377_, _20376_);
  and (_20378_, _01367_, _23768_);
  and (_20379_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_11203_, _20379_, _20378_);
  and (_20380_, _10475_, _26170_);
  and (_20381_, _10477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_11209_, _20381_, _20380_);
  and (_20382_, _00428_, _26085_);
  and (_20383_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_11211_, _20383_, _20382_);
  and (_20384_, _00428_, _26170_);
  and (_20385_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_27223_, _20385_, _20384_);
  and (_20386_, _15044_, _26242_);
  and (_20387_, _15046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_11215_, _20387_, _20386_);
  and (_20388_, _00400_, _26242_);
  and (_20389_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_27222_, _20389_, _20388_);
  and (_20390_, _00400_, _25886_);
  and (_20391_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_27220_, _20391_, _20390_);
  and (_20392_, _15029_, _23768_);
  and (_20393_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_11223_, _20393_, _20392_);
  and (_20394_, _15029_, _26170_);
  and (_20395_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_11225_, _20395_, _20394_);
  and (_20396_, _00292_, _25886_);
  and (_20397_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_11229_, _20397_, _20396_);
  and (_20398_, _04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  and (_20399_, _04148_, _26242_);
  or (_11232_, _20399_, _20398_);
  and (_20400_, _15029_, _25886_);
  and (_20401_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_11234_, _20401_, _20400_);
  and (_20402_, _00266_, _23830_);
  and (_20403_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_11236_, _20403_, _20402_);
  and (_20404_, _15029_, _26085_);
  and (_20405_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_11238_, _20405_, _20404_);
  and (_20406_, _00185_, _25886_);
  and (_20407_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_11240_, _20407_, _20406_);
  and (_20408_, _00185_, _25927_);
  and (_20409_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_27183_, _20409_, _20408_);
  and (_20410_, _15029_, _26185_);
  and (_20411_, _15032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_11244_, _20411_, _20410_);
  and (_20412_, _00171_, _23830_);
  and (_20413_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_11246_, _20413_, _20412_);
  and (_20414_, _00171_, _26170_);
  and (_20415_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_11248_, _20415_, _20414_);
  and (_20416_, _19653_, _25886_);
  and (_20417_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_11251_, _20417_, _20416_);
  and (_20418_, _14404_, _26170_);
  and (_20419_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_11256_, _20419_, _20418_);
  and (_20420_, _00155_, _26185_);
  and (_20421_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_11258_, _20421_, _20420_);
  and (_20422_, _00155_, _26170_);
  and (_20423_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_11260_, _20423_, _20422_);
  and (_20424_, _15017_, _23768_);
  and (_20425_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_26960_, _20425_, _20424_);
  and (_20426_, _00133_, _26242_);
  and (_20427_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_11265_, _20427_, _20426_);
  and (_20428_, _00133_, _25886_);
  and (_20429_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_27116_, _20429_, _20428_);
  and (_20430_, _14404_, _25927_);
  and (_20431_, _14406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_11269_, _20431_, _20430_);
  and (_20432_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_20433_, _04113_, _26185_);
  or (_11271_, _20433_, _20432_);
  and (_20434_, _00119_, _26242_);
  and (_20435_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_11274_, _20435_, _20434_);
  and (_20436_, _02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  and (_20437_, _02019_, _25927_);
  or (_11276_, _20437_, _20436_);
  and (_20438_, _00119_, _25886_);
  and (_20439_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_11278_, _20439_, _20438_);
  and (_20440_, _00119_, _25927_);
  and (_20441_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_11280_, _20441_, _20440_);
  and (_20442_, _09305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_20443_, _09304_, _25927_);
  or (_11282_, _20443_, _20442_);
  and (_20444_, _00105_, _26085_);
  and (_20445_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_11284_, _20445_, _20444_);
  and (_20446_, _00105_, _26170_);
  and (_20447_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_27152_, _20447_, _20446_);
  and (_20448_, _01367_, _26185_);
  and (_20449_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_27229_, _20449_, _20448_);
  and (_20450_, _01367_, _26170_);
  and (_20451_, _01369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_11289_, _20451_, _20450_);
  and (_20452_, _00428_, _26242_);
  and (_20453_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_11291_, _20453_, _20452_);
  and (_20454_, _15017_, _25927_);
  and (_20455_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_11293_, _20455_, _20454_);
  and (_20456_, _15017_, _23830_);
  and (_20457_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_11295_, _20457_, _20456_);
  and (_20458_, _00400_, _23768_);
  and (_20459_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_11297_, _20459_, _20458_);
  and (_20460_, _00292_, _23768_);
  and (_20461_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_11299_, _20461_, _20460_);
  and (_20462_, _00266_, _25927_);
  and (_20463_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_11301_, _20463_, _20462_);
  and (_20464_, _00185_, _26085_);
  and (_20465_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_11303_, _20465_, _20464_);
  and (_20466_, _15017_, _26085_);
  and (_20467_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_26961_, _20467_, _20466_);
  and (_20468_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_20469_, _04113_, _26085_);
  or (_27176_, _20469_, _20468_);
  and (_20470_, _00171_, _26185_);
  and (_20471_, _00173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_11309_, _20471_, _20470_);
  and (_20472_, _02102_, _26085_);
  and (_20473_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_11313_, _20473_, _20472_);
  and (_20474_, _15017_, _26242_);
  and (_20475_, _15019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_11316_, _20475_, _20474_);
  and (_20476_, _00133_, _23768_);
  and (_20477_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_11318_, _20477_, _20476_);
  and (_20478_, _00119_, _26085_);
  and (_20479_, _00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_11323_, _20479_, _20478_);
  and (_20480_, _00105_, _26242_);
  and (_20481_, _00107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_11326_, _20481_, _20480_);
  and (_20482_, _26073_, _25927_);
  and (_20483_, _26075_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_11328_, _20483_, _20482_);
  and (_20484_, _14408_, _25886_);
  and (_20485_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_11330_, _20485_, _20484_);
  and (_20486_, _00428_, _25886_);
  and (_20487_, _00430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_27224_, _20487_, _20486_);
  and (_20488_, _00400_, _23830_);
  and (_20489_, _00402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_27221_, _20489_, _20488_);
  and (_20490_, _00292_, _23830_);
  and (_20491_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_11337_, _20491_, _20490_);
  and (_20492_, _00266_, _26085_);
  and (_20493_, _00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_11339_, _20493_, _20492_);
  and (_20494_, _00155_, _25886_);
  and (_20495_, _00157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_11344_, _20495_, _20494_);
  and (_20496_, _00133_, _23830_);
  and (_20497_, _00135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_11346_, _20497_, _20496_);
  and (_20498_, _15009_, _23768_);
  and (_20499_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_11349_, _20499_, _20498_);
  and (_20500_, _15009_, _23830_);
  and (_20501_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_11351_, _20501_, _20500_);
  and (_20502_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  and (_20503_, _04143_, _26170_);
  or (_11353_, _20503_, _20502_);
  and (_20504_, _00185_, _26185_);
  and (_20505_, _00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_11356_, _20505_, _20504_);
  and (_20506_, _14408_, _26170_);
  and (_20507_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_11360_, _20507_, _20506_);
  and (_20508_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  and (_20509_, _06617_, _23830_);
  or (_11362_, _20509_, _20508_);
  and (_20510_, _00292_, _26085_);
  and (_20511_, _00294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_11365_, _20511_, _20510_);
  and (_20512_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  and (_20513_, _06617_, _26185_);
  or (_27173_, _20513_, _20512_);
  and (_20514_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  and (_20515_, _02576_, _23830_);
  or (_27077_, _20515_, _20514_);
  and (_20516_, _15009_, _26085_);
  and (_20517_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_26962_, _20517_, _20516_);
  and (_20518_, _15009_, _26242_);
  and (_20519_, _15011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_11398_, _20519_, _20518_);
  and (_20520_, _02519_, _25927_);
  and (_20521_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_11403_, _20521_, _20520_);
  and (_20522_, _02026_, _26085_);
  and (_20523_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_11418_, _20523_, _20522_);
  and (_20524_, _02480_, _23768_);
  and (_20525_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_11423_, _20525_, _20524_);
  and (_20526_, _04812_, _26170_);
  and (_20527_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_11429_, _20527_, _20526_);
  and (_20528_, _19653_, _26170_);
  and (_20529_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_11432_, _20529_, _20528_);
  and (_20530_, _02570_, _26170_);
  and (_20531_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_11446_, _20531_, _20530_);
  and (_20532_, _02609_, _26185_);
  and (_20533_, _02611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_11448_, _20533_, _20532_);
  and (_20534_, _19653_, _25927_);
  and (_20535_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_11451_, _20535_, _20534_);
  and (_20536_, _02102_, _26242_);
  and (_20537_, _02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_26982_, _20537_, _20536_);
  and (_20538_, _14999_, _23768_);
  and (_20539_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_11455_, _20539_, _20538_);
  and (_20540_, _05799_, _25927_);
  and (_20541_, _05801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_26976_, _20541_, _20540_);
  and (_20542_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  and (_20543_, _06617_, _26085_);
  or (_11459_, _20543_, _20542_);
  and (_20544_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _01425_);
  and (_20545_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_20546_, _20545_, _20544_);
  and (_26931_[7], _20546_, _23049_);
  and (_20547_, _04812_, _25927_);
  and (_20548_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or (_11466_, _20548_, _20547_);
  and (_20549_, _14408_, _26085_);
  and (_20550_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_11479_, _20550_, _20549_);
  and (_20551_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  and (_20552_, _10218_, _26085_);
  or (_11481_, _20552_, _20551_);
  and (_20553_, _16208_, _26170_);
  and (_20554_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_11491_, _20554_, _20553_);
  and (_20555_, _22928_, _22879_);
  and (_20556_, _20555_, _22964_);
  and (_20557_, _22737_, _22743_);
  and (_20558_, _20557_, _01913_);
  and (_20559_, _20558_, _22823_);
  not (_20560_, _22852_);
  and (_20561_, _22905_, _20560_);
  and (_20562_, _20561_, _20559_);
  and (_20563_, _22800_, _22773_);
  and (_20564_, _20563_, _20562_);
  and (_26930_, _20564_, _20556_);
  and (_20565_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  and (_20566_, _10218_, _23830_);
  or (_11503_, _20566_, _20565_);
  and (_20567_, _19653_, _26085_);
  and (_20568_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_11520_, _20568_, _20567_);
  and (_20569_, _10220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  and (_20570_, _10218_, _25886_);
  or (_11523_, _20570_, _20569_);
  and (_20571_, _14408_, _23830_);
  and (_20572_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_11534_, _20572_, _20571_);
  and (_20573_, _14999_, _25886_);
  and (_20574_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_11536_, _20574_, _20573_);
  and (_11550_, _00900_, _23049_);
  and (_11552_, _00948_, _23049_);
  and (_20575_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  and (_20576_, _06617_, _26242_);
  or (_11554_, _20576_, _20575_);
  and (_11556_, _01086_, _23049_);
  and (_11558_, _01137_, _23049_);
  and (_11561_, _25840_, _23049_);
  and (_11563_, _00483_, _23049_);
  and (_11565_, _00638_, _23049_);
  and (_11567_, _00688_, _23049_);
  and (_20577_, _04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_20578_, _04113_, _23768_);
  or (_27174_, _20578_, _20577_);
  and (_20579_, _26308_, _23830_);
  and (_20580_, _26311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_27270_, _20580_, _20579_);
  and (_20581_, _04145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  and (_20582_, _04143_, _25927_);
  or (_27180_, _20582_, _20581_);
  and (_11572_, _00998_, _23049_);
  and (_11574_, _01199_, _23049_);
  and (_11576_, _00530_, _23049_);
  and (_11578_, _00743_, _23049_);
  and (_11581_, _01041_, _23049_);
  and (_11585_, _00575_, _23049_);
  and (_20583_, _14999_, _23830_);
  and (_20584_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_26964_, _20584_, _20583_);
  and (_20585_, _02590_, _23830_);
  and (_20586_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_27252_, _20586_, _20585_);
  and (_20587_, _14999_, _26085_);
  and (_20588_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_26965_, _20588_, _20587_);
  and (_20589_, _02800_, _26185_);
  and (_20590_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_27119_, _20590_, _20589_);
  or (_20591_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_26946_, _20591_, _02893_);
  nor (_20592_, _24794_, _24804_);
  and (_20593_, _24794_, _24804_);
  or (_20594_, _20593_, _20592_);
  and (_11628_, _20594_, _23049_);
  and (_20595_, _15146_, _26085_);
  and (_20596_, _15148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_27279_, _20596_, _20595_);
  and (_20597_, _02577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  and (_20598_, _02576_, _26085_);
  or (_27078_, _20598_, _20597_);
  and (_20599_, _14639_, _26085_);
  and (_20600_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_26991_, _20600_, _20599_);
  and (_20601_, _15231_, _23830_);
  and (_20602_, _15233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_27239_, _20602_, _20601_);
  and (_20603_, _14639_, _23830_);
  and (_20604_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_26990_, _20604_, _20603_);
  and (_20605_, _14639_, _25886_);
  and (_20606_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_26989_, _20606_, _20605_);
  and (_20607_, _02026_, _26185_);
  and (_20608_, _02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_27300_, _20608_, _20607_);
  and (_20609_, _14999_, _26185_);
  and (_20610_, _15001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_26966_, _20610_, _20609_);
  and (_20611_, _14991_, _23768_);
  and (_20612_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_26967_, _20612_, _20611_);
  and (_20613_, _02590_, _26085_);
  and (_20614_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_27253_, _20614_, _20613_);
  and (_20615_, _16208_, _25927_);
  and (_20616_, _16210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_27264_, _20616_, _20615_);
  and (_20617_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  and (_20618_, _04243_, _26242_);
  or (_27170_, _20618_, _20617_);
  and (_20619_, _14408_, _23768_);
  and (_20620_, _14410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_26994_, _20620_, _20619_);
  and (_20621_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  and (_20622_, _06617_, _23768_);
  or (_27171_, _20622_, _20621_);
  and (_20623_, _14639_, _26242_);
  and (_20624_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or (_26993_, _20624_, _20623_);
  and (_20625_, _14639_, _26185_);
  and (_20626_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or (_26992_, _20626_, _20625_);
  and (_20627_, _19653_, _26185_);
  and (_20628_, _19655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_27248_, _20628_, _20627_);
  and (_20629_, _02329_, _23768_);
  and (_20630_, _02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_27275_, _20630_, _20629_);
  and (_20631_, _25943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_20632_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_20633_, _25943_, _20632_);
  or (_20634_, _20633_, _20631_);
  and (_26915_[15], _20634_, _23049_);
  and (_20635_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20636_, _20635_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20637_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_20638_, _20637_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_20639_, _20638_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_20640_, _20639_, _20636_);
  and (_20641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_20642_, _20641_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_20643_, _20642_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20644_, _20643_, _20640_);
  and (_20645_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20646_, _20645_, _20644_);
  and (_20647_, _20646_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20648_, _20646_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20649_, _20648_, _20647_);
  nor (_20650_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20651_, _20650_);
  and (_20652_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26017_);
  and (_20653_, _26021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_20654_, _20653_, _20652_);
  and (_20655_, _20654_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20657_, _20656_, _20655_);
  not (_20658_, _20657_);
  and (_20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20660_, _20659_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_20661_, _20660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20662_, _20636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20663_, _20662_, _20661_);
  nor (_20664_, _20663_, _05411_);
  and (_20665_, _20663_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_20666_, _20665_, _20664_);
  nor (_20667_, _20666_, _20658_);
  nor (_20668_, _20663_, _04941_);
  and (_20669_, _20663_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_20670_, _20669_, _20668_);
  nor (_20671_, _20670_, _20657_);
  nor (_20672_, _20671_, _20667_);
  nor (_20673_, _20672_, _20651_);
  and (_20674_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26013_);
  not (_20675_, _20674_);
  nor (_20676_, _20663_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_20677_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_20678_, _20663_, _20677_);
  or (_20679_, _20678_, _20657_);
  or (_20680_, _20679_, _20676_);
  and (_20681_, _20663_, _04968_);
  nor (_20682_, _20663_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_20683_, _20682_, _20681_);
  or (_20684_, _20683_, _20658_);
  and (_20685_, _20684_, _20680_);
  nor (_20686_, _20685_, _20675_);
  nor (_20687_, _20686_, _20673_);
  not (_20688_, _20659_);
  not (_20689_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_20690_, _20663_, _20689_);
  nor (_20691_, _20663_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_20692_, _20691_, _20657_);
  or (_20693_, _20692_, _20690_);
  nor (_20694_, _20663_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_20695_, _20663_);
  or (_20696_, _20695_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_20697_, _20696_, _20657_);
  or (_20698_, _20697_, _20694_);
  and (_20699_, _20698_, _20693_);
  nor (_20700_, _20699_, _20688_);
  and (_20701_, _26017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20702_, _20701_);
  nor (_20703_, _20663_, _05474_);
  and (_20704_, _20663_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_20705_, _20704_, _20703_);
  nor (_20706_, _20705_, _20658_);
  not (_20707_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_20708_, _20663_, _20707_);
  and (_20709_, _20663_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_20710_, _20709_, _20708_);
  nor (_20711_, _20710_, _20657_);
  nor (_20712_, _20711_, _20706_);
  nor (_20713_, _20712_, _20702_);
  nor (_20714_, _20713_, _20700_);
  and (_20715_, _20714_, _20687_);
  and (_20716_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_20717_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_20718_, _20717_, _20716_);
  and (_20719_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_20720_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_20721_, _20720_, _20719_);
  and (_20722_, _20721_, _20718_);
  and (_20723_, _20722_, _20658_);
  and (_20724_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_20725_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_20726_, _20725_, _20724_);
  and (_20727_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_20728_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_20729_, _20728_, _20727_);
  and (_20730_, _20729_, _20726_);
  and (_20731_, _20730_, _20657_);
  or (_20732_, _20731_, _20663_);
  nor (_20733_, _20732_, _20723_);
  and (_20734_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_20735_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_20736_, _20735_, _20734_);
  and (_20737_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_20738_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_20739_, _20738_, _20737_);
  and (_20740_, _20739_, _20736_);
  nor (_20741_, _20740_, _20657_);
  and (_20742_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_20743_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_20744_, _20743_, _20742_);
  and (_20745_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_20746_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_20747_, _20746_, _20745_);
  and (_20748_, _20747_, _20744_);
  nor (_20749_, _20748_, _20658_);
  or (_20750_, _20749_, _20741_);
  and (_20751_, _20750_, _20663_);
  nor (_20752_, _20751_, _20733_);
  nor (_20753_, _20752_, _20715_);
  and (_20754_, _20753_, _20649_);
  and (_20755_, _20644_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_20756_, _20755_, _26063_);
  nor (_20757_, _20755_, _26063_);
  nor (_20758_, _20757_, _20756_);
  not (_20759_, _20758_);
  and (_20760_, _20759_, _20753_);
  nor (_20761_, _20644_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20762_, _20761_, _20755_);
  and (_20763_, _20762_, _20753_);
  nor (_20764_, _20759_, _20753_);
  nor (_20765_, _20764_, _20760_);
  and (_20766_, _20642_, _20640_);
  nor (_20767_, _20766_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_20768_, _20766_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20769_, _20768_, _20767_);
  and (_20770_, _20769_, _20753_);
  nor (_20771_, _20769_, _20753_);
  and (_20772_, _20640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_20773_, _20772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20774_, _20773_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20775_, _20774_, _20766_);
  and (_20776_, _20775_, _20753_);
  nor (_20777_, _20775_, _20753_);
  nor (_20778_, _20777_, _20776_);
  nor (_20779_, _20772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20780_, _20779_, _20773_);
  and (_20781_, _20780_, _20753_);
  nor (_20782_, _20780_, _20753_);
  nor (_20783_, _20640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20784_, _20783_, _20772_);
  and (_20785_, _20784_, _20753_);
  and (_20786_, _20638_, _20636_);
  nor (_20787_, _20786_, _26040_);
  and (_20788_, _20786_, _26040_);
  nor (_20789_, _20788_, _20787_);
  not (_20790_, _20789_);
  and (_20791_, _20790_, _20753_);
  nor (_20792_, _20790_, _20753_);
  and (_20793_, _20637_, _20636_);
  nor (_20794_, _20793_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20795_, _20794_, _20786_);
  and (_20796_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_20797_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_20798_, _20797_, _20796_);
  and (_20799_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_20800_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_20801_, _20800_, _20799_);
  and (_20802_, _20801_, _20798_);
  and (_20803_, _20802_, _20658_);
  and (_20804_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_20805_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_20806_, _20805_, _20804_);
  and (_20807_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_20808_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_20809_, _20808_, _20807_);
  and (_20810_, _20809_, _20806_);
  and (_20811_, _20810_, _20657_);
  or (_20812_, _20811_, _20663_);
  nor (_20813_, _20812_, _20803_);
  and (_20814_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_20815_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_20816_, _20815_, _20814_);
  and (_20817_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_20818_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_20819_, _20818_, _20817_);
  and (_20820_, _20819_, _20816_);
  and (_20821_, _20820_, _20658_);
  and (_20822_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_20823_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20824_, _20823_, _20822_);
  and (_20825_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_20826_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_20827_, _20826_, _20825_);
  and (_20828_, _20827_, _20824_);
  and (_20829_, _20828_, _20657_);
  nor (_20830_, _20829_, _20821_);
  and (_20831_, _20830_, _20663_);
  nor (_20832_, _20831_, _20813_);
  nor (_20833_, _20832_, _20715_);
  and (_20834_, _20833_, _20795_);
  nor (_20835_, _20833_, _20795_);
  nor (_20836_, _20835_, _20834_);
  not (_20837_, _20836_);
  and (_20838_, _20636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20839_, _20838_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_20840_, _20839_, _20793_);
  and (_20841_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_20842_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_20843_, _20842_, _20841_);
  and (_20844_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_20845_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_20846_, _20845_, _20844_);
  and (_20847_, _20846_, _20843_);
  and (_20848_, _20847_, _20658_);
  and (_20849_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_20850_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_20851_, _20850_, _20849_);
  and (_20852_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_20853_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_20854_, _20853_, _20852_);
  and (_20855_, _20854_, _20851_);
  and (_20856_, _20855_, _20657_);
  or (_20857_, _20856_, _20663_);
  nor (_20858_, _20857_, _20848_);
  and (_20859_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_20860_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_20861_, _20860_, _20859_);
  and (_20862_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_20863_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_20864_, _20863_, _20862_);
  and (_20865_, _20864_, _20861_);
  nor (_20866_, _20865_, _20657_);
  and (_20867_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_20868_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_20869_, _20868_, _20867_);
  and (_20870_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_20871_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_20872_, _20871_, _20870_);
  and (_20873_, _20872_, _20869_);
  nor (_20874_, _20873_, _20658_);
  or (_20875_, _20874_, _20866_);
  and (_20876_, _20875_, _20663_);
  nor (_20877_, _20876_, _20858_);
  nor (_20878_, _20877_, _20715_);
  and (_20879_, _20878_, _20840_);
  nor (_20880_, _20878_, _20840_);
  nor (_20881_, _20880_, _20879_);
  not (_20882_, _20881_);
  and (_20883_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_20884_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_20885_, _20884_, _20883_);
  and (_20886_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_20887_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_20888_, _20887_, _20886_);
  and (_20889_, _20888_, _20885_);
  and (_20890_, _20889_, _20657_);
  and (_20891_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_20892_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_20893_, _20892_, _20891_);
  and (_20894_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_20895_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_20896_, _20895_, _20894_);
  and (_20897_, _20896_, _20893_);
  and (_20898_, _20897_, _20658_);
  or (_20899_, _20898_, _20663_);
  nor (_20900_, _20899_, _20890_);
  and (_20901_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_20902_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_20903_, _20902_, _20901_);
  and (_20904_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_20905_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_20906_, _20905_, _20904_);
  and (_20907_, _20906_, _20903_);
  nor (_20908_, _20907_, _20657_);
  and (_20909_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_20910_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20911_, _20910_, _20909_);
  and (_20912_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_20913_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20914_, _20913_, _20912_);
  and (_20915_, _20914_, _20911_);
  nor (_20916_, _20915_, _20658_);
  or (_20917_, _20916_, _20908_);
  and (_20918_, _20917_, _20663_);
  nor (_20919_, _20918_, _20900_);
  nor (_20920_, _20919_, _20715_);
  nor (_20921_, _20636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20922_, _20921_, _20838_);
  and (_20923_, _20922_, _20920_);
  nor (_20924_, _20635_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20925_, _20924_, _20636_);
  and (_20926_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_20927_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_20928_, _20927_, _20926_);
  and (_20929_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_20930_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_20931_, _20930_, _20929_);
  and (_20932_, _20931_, _20928_);
  and (_20933_, _20932_, _20658_);
  and (_20934_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_20935_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_20936_, _20935_, _20934_);
  and (_20937_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_20938_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_20939_, _20938_, _20937_);
  and (_20940_, _20939_, _20936_);
  and (_20941_, _20940_, _20657_);
  or (_20942_, _20941_, _20663_);
  nor (_20943_, _20942_, _20933_);
  and (_20944_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_20945_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_20946_, _20945_, _20944_);
  and (_20947_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_20948_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_20949_, _20948_, _20947_);
  and (_20950_, _20949_, _20946_);
  and (_20951_, _20950_, _20658_);
  and (_20952_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_20953_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20954_, _20953_, _20952_);
  and (_20955_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_20956_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20957_, _20956_, _20955_);
  and (_20958_, _20957_, _20954_);
  and (_20959_, _20958_, _20657_);
  nor (_20960_, _20959_, _20951_);
  and (_20961_, _20960_, _20663_);
  nor (_20962_, _20961_, _20943_);
  nor (_20963_, _20962_, _20715_);
  and (_20964_, _20963_, _20925_);
  nor (_20965_, _20963_, _20925_);
  nor (_20966_, _20965_, _20964_);
  not (_20967_, _20966_);
  not (_20968_, _20654_);
  and (_20969_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_20970_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_20971_, _20970_, _20969_);
  and (_20972_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_20973_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_20974_, _20973_, _20972_);
  and (_20975_, _20974_, _20971_);
  and (_20976_, _20975_, _20658_);
  and (_20977_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_20978_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_20979_, _20978_, _20977_);
  and (_20980_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_20981_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_20982_, _20981_, _20980_);
  and (_20983_, _20982_, _20979_);
  and (_20984_, _20983_, _20657_);
  or (_20985_, _20984_, _20663_);
  nor (_20986_, _20985_, _20976_);
  and (_20987_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_20988_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_20989_, _20988_, _20987_);
  and (_20990_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_20991_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_20992_, _20991_, _20990_);
  and (_20993_, _20992_, _20989_);
  nor (_20994_, _20993_, _20657_);
  and (_20995_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_20996_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_20997_, _20996_, _20995_);
  and (_20998_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_20999_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_21000_, _20999_, _20998_);
  and (_21001_, _21000_, _20997_);
  nor (_21002_, _21001_, _20658_);
  or (_21003_, _21002_, _20994_);
  and (_21004_, _21003_, _20663_);
  nor (_21005_, _21004_, _20986_);
  nor (_21006_, _21005_, _20715_);
  and (_21007_, _21006_, _20968_);
  and (_21008_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_21009_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_21010_, _21009_, _21008_);
  and (_21011_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_21012_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_21013_, _21012_, _21011_);
  and (_21014_, _21013_, _21010_);
  and (_21015_, _21014_, _20658_);
  and (_21016_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_21017_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_21018_, _21017_, _21016_);
  and (_21019_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_21020_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_21021_, _21020_, _21019_);
  and (_21022_, _21021_, _21018_);
  and (_21023_, _21022_, _20657_);
  or (_21024_, _21023_, _20663_);
  nor (_21025_, _21024_, _21015_);
  and (_21026_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21027_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_21028_, _21027_, _21026_);
  and (_21029_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_21030_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_21031_, _21030_, _21029_);
  and (_21032_, _21031_, _21028_);
  nor (_21033_, _21032_, _20657_);
  and (_21034_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_21035_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_21036_, _21035_, _21034_);
  and (_21037_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21038_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_21039_, _21038_, _21037_);
  and (_21040_, _21039_, _21036_);
  nor (_21041_, _21040_, _20658_);
  or (_21042_, _21041_, _21033_);
  and (_21043_, _21042_, _20663_);
  nor (_21044_, _21043_, _21025_);
  nor (_21045_, _21044_, _20715_);
  and (_21046_, _21045_, _26017_);
  and (_21047_, _20674_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_21048_, _20659_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_21049_, _21048_, _21047_);
  and (_21050_, _20701_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_21051_, _20650_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_21052_, _21051_, _21050_);
  and (_21053_, _21052_, _21049_);
  and (_21054_, _21053_, _20658_);
  and (_21055_, _20674_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_21056_, _20650_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_21057_, _21056_, _21055_);
  and (_21058_, _20701_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_21059_, _20659_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _21057_);
  and (_21062_, _21061_, _20657_);
  or (_21063_, _21062_, _20663_);
  nor (_21064_, _21063_, _21054_);
  and (_21065_, _20674_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_21066_, _20659_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_21067_, _21066_, _21065_);
  and (_21068_, _20701_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_21069_, _20650_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_21070_, _21069_, _21068_);
  and (_21071_, _21070_, _21067_);
  nor (_21072_, _21071_, _20657_);
  and (_21073_, _20701_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_21074_, _20659_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_21075_, _21074_, _21073_);
  and (_21076_, _20674_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_21077_, _20650_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_21078_, _21077_, _21076_);
  and (_21079_, _21078_, _21075_);
  nor (_21080_, _21079_, _20658_);
  or (_21081_, _21080_, _21072_);
  and (_21082_, _21081_, _20663_);
  nor (_21083_, _21082_, _21064_);
  nor (_21084_, _21083_, _20715_);
  and (_21085_, _21084_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21086_, _21045_, _26017_);
  nor (_21087_, _21086_, _21046_);
  and (_21088_, _21087_, _21085_);
  nor (_21089_, _21088_, _21046_);
  nor (_21090_, _21006_, _20968_);
  nor (_21091_, _21090_, _21007_);
  not (_21092_, _21091_);
  nor (_21093_, _21092_, _21089_);
  nor (_21094_, _21093_, _21007_);
  nor (_21095_, _21094_, _20967_);
  nor (_21096_, _21095_, _20964_);
  nor (_21097_, _20922_, _20920_);
  nor (_21098_, _21097_, _20923_);
  not (_21099_, _21098_);
  nor (_21100_, _21099_, _21096_);
  nor (_21101_, _21100_, _20923_);
  nor (_21102_, _21101_, _20882_);
  nor (_21103_, _21102_, _20879_);
  nor (_21104_, _21103_, _20837_);
  nor (_21105_, _21104_, _20834_);
  nor (_21106_, _21105_, _20792_);
  or (_21107_, _21106_, _20791_);
  nor (_21108_, _20784_, _20753_);
  nor (_21109_, _21108_, _20785_);
  and (_21110_, _21109_, _21107_);
  nor (_21111_, _21110_, _20785_);
  nor (_21112_, _21111_, _20782_);
  or (_21113_, _21112_, _20781_);
  and (_21114_, _21113_, _20778_);
  nor (_21115_, _21114_, _20776_);
  nor (_21116_, _21115_, _20771_);
  nor (_21117_, _21116_, _20770_);
  nor (_21118_, _20762_, _20753_);
  nor (_21119_, _21118_, _20763_);
  not (_21120_, _21119_);
  nor (_21121_, _21120_, _21117_);
  and (_21122_, _21121_, _20765_);
  or (_21123_, _21122_, _20763_);
  nor (_21124_, _21123_, _20760_);
  nor (_21125_, _20753_, _20649_);
  nor (_21126_, _21125_, _20754_);
  not (_21127_, _21126_);
  nor (_21128_, _21127_, _21124_);
  nor (_21129_, _21128_, _20754_);
  nor (_21130_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_21131_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_21132_, _21131_, _21130_);
  not (_21133_, _21132_);
  and (_21134_, _21133_, _20647_);
  nor (_21135_, _21133_, _20647_);
  nor (_21136_, _21135_, _21134_);
  not (_21137_, _21136_);
  and (_21138_, _21137_, _20753_);
  nor (_21139_, _21137_, _20753_);
  nor (_21140_, _21139_, _21138_);
  not (_21141_, _21140_);
  nand (_21142_, _21141_, _21129_);
  or (_21143_, _21141_, _21129_);
  and (_21144_, _21143_, _21142_);
  and (_21145_, _21127_, _21124_);
  nor (_21146_, _21145_, _21128_);
  and (_21147_, _21146_, _26009_);
  nor (_21148_, _21146_, _26009_);
  nor (_21149_, _21121_, _20763_);
  nor (_21150_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_21151_, _20758_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_21152_, _21151_, _21150_);
  nand (_21153_, _21152_, _20753_);
  or (_21154_, _21152_, _20753_);
  and (_21155_, _21154_, _21153_);
  not (_21156_, _21155_);
  nand (_21157_, _21156_, _21149_);
  or (_21158_, _21156_, _21149_);
  and (_21159_, _21158_, _21157_);
  and (_21160_, _21120_, _21117_);
  nor (_21161_, _21160_, _21121_);
  nor (_21162_, _21161_, _26001_);
  and (_21163_, _21161_, _26001_);
  nor (_21164_, _20769_, _25996_);
  and (_21165_, _20769_, _25996_);
  or (_21166_, _21165_, _21164_);
  nand (_21167_, _21166_, _20753_);
  or (_21168_, _21166_, _20753_);
  and (_21169_, _21168_, _21167_);
  not (_21170_, _21169_);
  nand (_21171_, _21170_, _21115_);
  or (_21172_, _21170_, _21115_);
  and (_21173_, _21172_, _21171_);
  nor (_21174_, _21113_, _20778_);
  nor (_21175_, _21174_, _21114_);
  nor (_21176_, _21175_, _25990_);
  and (_21177_, _21175_, _25990_);
  nor (_21178_, _21109_, _21107_);
  nor (_21179_, _21178_, _21110_);
  nand (_21180_, _21179_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_21181_, _21179_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_21182_, _21181_, _21180_);
  not (_21183_, _20753_);
  nor (_21184_, _20780_, _25985_);
  and (_21185_, _20780_, _25985_);
  or (_21186_, _21185_, _21184_);
  nand (_21187_, _21186_, _21183_);
  or (_21188_, _21186_, _21183_);
  and (_21189_, _21188_, _21187_);
  or (_21190_, _21189_, _21111_);
  nand (_21191_, _21189_, _21111_);
  and (_21192_, _21191_, _21190_);
  nor (_21193_, _20791_, _20792_);
  nor (_21194_, _21193_, _21105_);
  and (_21195_, _21193_, _21105_);
  or (_21196_, _21195_, _21194_);
  nor (_21197_, _21196_, _25976_);
  and (_21198_, _21196_, _25976_);
  and (_21199_, _21103_, _20837_);
  nor (_21200_, _21199_, _21104_);
  and (_21201_, _21200_, _25971_);
  nor (_21202_, _21200_, _25971_);
  and (_21203_, _21101_, _20882_);
  nor (_21204_, _21203_, _21102_);
  nor (_21205_, _21204_, _25966_);
  and (_21206_, _21204_, _25966_);
  and (_21207_, _21099_, _21096_);
  nor (_21208_, _21207_, _21100_);
  nor (_21209_, _21208_, _25962_);
  and (_21210_, _21094_, _20967_);
  nor (_21211_, _21210_, _21095_);
  nor (_21212_, _21211_, _25958_);
  and (_21213_, _21211_, _25958_);
  and (_21214_, _21092_, _21089_);
  nor (_21215_, _21214_, _21093_);
  and (_21216_, _21215_, _25953_);
  and (_21217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21218_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21219_, _21218_, _21217_);
  and (_21220_, _21219_, _21084_);
  nor (_21221_, _21219_, _21084_);
  or (_21222_, _21221_, _21220_);
  nor (_21223_, _21087_, _21085_);
  nor (_21224_, _21223_, _21088_);
  nor (_21225_, _21224_, _25949_);
  and (_21226_, _21224_, _25949_);
  or (_21227_, _21226_, _21225_);
  or (_21228_, _21227_, _21222_);
  nor (_21229_, _21215_, _25953_);
  or (_21230_, _21229_, _21228_);
  or (_21231_, _21230_, _21216_);
  or (_21232_, _21231_, _21213_);
  or (_21233_, _21232_, _21212_);
  and (_21234_, _21208_, _25962_);
  or (_21235_, _21234_, _21233_);
  or (_21236_, _21235_, _21209_);
  or (_21237_, _21236_, _21206_);
  or (_21238_, _21237_, _21205_);
  or (_21239_, _21238_, _21202_);
  or (_21240_, _21239_, _21201_);
  or (_21241_, _21240_, _21198_);
  or (_21242_, _21241_, _21197_);
  or (_21243_, _21242_, _21192_);
  or (_21244_, _21243_, _21182_);
  or (_21245_, _21244_, _21177_);
  or (_21246_, _21245_, _21176_);
  or (_21247_, _21246_, _21173_);
  or (_21248_, _21247_, _21163_);
  or (_21249_, _21248_, _21162_);
  or (_21250_, _21249_, _21159_);
  or (_21251_, _21250_, _21148_);
  or (_21252_, _21251_, _21147_);
  or (_21253_, _21252_, _21144_);
  or (_21254_, \oc8051_symbolic_cxrom1.regvalid [1], _25958_);
  and (_21255_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21256_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21257_, _21256_, _21255_);
  and (_21258_, _21257_, _21254_);
  or (_21259_, \oc8051_symbolic_cxrom1.regvalid [13], _25958_);
  or (_21260_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21261_, _21260_, _21259_);
  and (_21262_, _25953_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21263_, _21262_, _21261_);
  or (_21264_, _21263_, _21258_);
  nor (_21265_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21266_, _21265_, _25953_);
  nor (_21267_, _21266_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21268_, _21266_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21269_, _21268_, _21267_);
  and (_21270_, _21269_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_21271_, _21265_, _25953_);
  nor (_21272_, _21271_, _21266_);
  or (_21273_, _05532_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21274_, _21273_, _21272_);
  or (_21275_, _21274_, _21270_);
  and (_21276_, _21275_, _25949_);
  nand (_21277_, _21269_, _20677_);
  or (_21278_, _21269_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_21279_, _21278_, _21277_);
  or (_21280_, _21272_, _21279_);
  and (_21281_, _21280_, _21276_);
  or (_21282_, _21281_, _21264_);
  and (_21283_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21284_, \oc8051_symbolic_cxrom1.regvalid [0], _25958_);
  or (_21285_, _21284_, _21283_);
  and (_21286_, _21285_, _25953_);
  and (_21287_, \oc8051_symbolic_cxrom1.regvalid [4], _25958_);
  and (_21288_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21289_, _21288_, _21287_);
  and (_21290_, _21289_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21291_, _21290_, _21286_);
  and (_21292_, _21291_, _25949_);
  and (_21293_, _21255_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21294_, _21293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21295_, _21293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21296_, _21295_, _21294_);
  or (_21297_, _21296_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_21299_, _21298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_21300_, _21299_, _21293_);
  and (_21301_, _21300_, _21259_);
  and (_21302_, _21301_, _21297_);
  or (_21303_, _21296_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_21304_, _21300_);
  nand (_21305_, _21296_, _05592_);
  and (_21306_, _21305_, _21304_);
  and (_21307_, _21306_, _21303_);
  or (_21308_, _21307_, _21302_);
  and (_21309_, _21308_, _21292_);
  or (_21310_, _21296_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_21311_, \oc8051_symbolic_cxrom1.regvalid [15], _25958_);
  and (_21312_, _21311_, _21300_);
  and (_21313_, _21312_, _21310_);
  or (_21314_, _21296_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_21315_, _21296_, _20677_);
  and (_21316_, _21315_, _21304_);
  and (_21317_, _21316_, _21314_);
  or (_21318_, _21317_, _21313_);
  and (_21319_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21320_, \oc8051_symbolic_cxrom1.regvalid [6], _25958_);
  or (_21321_, _21320_, _25953_);
  or (_21322_, _21321_, _21319_);
  or (_21323_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21324_, \oc8051_symbolic_cxrom1.regvalid [10], _25958_);
  and (_21325_, _21324_, _21323_);
  or (_21326_, _21325_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21327_, _21326_, _21322_);
  and (_21328_, _21327_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21329_, _21289_, _21262_);
  or (_21330_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21331_, \oc8051_symbolic_cxrom1.regvalid [0], _25958_);
  and (_21332_, _21331_, _21255_);
  and (_21333_, _21332_, _21330_);
  or (_21334_, _21333_, _21329_);
  and (_21335_, _21334_, _21328_);
  and (_21336_, _21335_, _21318_);
  or (_21337_, _21336_, _21309_);
  or (_21338_, _21334_, _21327_);
  and (_21339_, _21338_, _25945_);
  and (_21340_, _21339_, _21337_);
  and (_21341_, _21340_, _21282_);
  or (_21342_, \oc8051_symbolic_cxrom1.regvalid [2], _25949_);
  or (_21343_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_21344_, _21343_, _21342_);
  or (_21345_, _21344_, _21269_);
  or (_21346_, \oc8051_symbolic_cxrom1.regvalid [10], _25949_);
  or (_21347_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_21348_, _21347_, _21346_);
  and (_21349_, _21348_, _21269_);
  nor (_21350_, _21349_, _21272_);
  and (_21351_, _21350_, _21345_);
  and (_21352_, _21269_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_21353_, _21287_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_21354_, _21353_, _21352_);
  and (_21355_, _21269_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_21356_, _21320_, _25949_);
  or (_21357_, _21356_, _21355_);
  and (_21358_, _21357_, _21272_);
  and (_21359_, _21358_, _21354_);
  or (_21360_, _21359_, _21351_);
  or (_21361_, _21296_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_21362_, \oc8051_symbolic_cxrom1.regvalid [14], _25958_);
  and (_21363_, _21362_, _21361_);
  or (_21364_, _21363_, _21304_);
  nand (_21365_, _21296_, _05656_);
  or (_21366_, _21296_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_21367_, _21366_, _21365_);
  or (_21368_, _21367_, _21300_);
  and (_21369_, _21368_, _21364_);
  or (_21370_, _21369_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_21371_, _21296_, _20689_);
  or (_21372_, _21296_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_21373_, _21372_, _21304_);
  and (_21374_, _21373_, _21371_);
  or (_21375_, _21296_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_21376_, \oc8051_symbolic_cxrom1.regvalid [12], _25958_);
  and (_21377_, _21376_, _21300_);
  and (_21378_, _21377_, _21375_);
  or (_21379_, _21378_, _25949_);
  or (_21380_, _21379_, _21374_);
  or (_21381_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21382_, _21381_, _21311_);
  or (_21383_, _21382_, _25953_);
  or (_21384_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21385_, \oc8051_symbolic_cxrom1.regvalid [11], _25958_);
  and (_21386_, _21385_, _21384_);
  or (_21387_, _21386_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21388_, _21387_, _21383_);
  and (_21389_, _21388_, _21298_);
  and (_21390_, _25949_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_21391_, _21261_, _25953_);
  or (_21392_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21393_, \oc8051_symbolic_cxrom1.regvalid [9], _25958_);
  and (_21394_, _21393_, _21392_);
  or (_21395_, _21394_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21396_, _21395_, _21391_);
  and (_21397_, _21396_, _21390_);
  or (_21398_, _21397_, _21389_);
  and (_21399_, _21388_, _25949_);
  or (_21400_, _21399_, _21264_);
  and (_21401_, _21400_, _21398_);
  and (_21402_, _21401_, _21380_);
  and (_21403_, _21402_, _21370_);
  and (_21404_, _21403_, _21360_);
  or (_21405_, _21404_, _21341_);
  nor (_21406_, _20650_, _26021_);
  and (_21407_, _20656_, _26017_);
  nor (_21408_, _21407_, _21406_);
  not (_21409_, _21408_);
  and (_21410_, _21406_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21411_, _21406_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21412_, _21411_, _21410_);
  and (_21413_, _21412_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21414_, _21412_, _04961_);
  or (_21415_, _21414_, _21413_);
  and (_21416_, _21415_, _21409_);
  nand (_21417_, _21412_, _04968_);
  nor (_21418_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21419_, _21418_);
  and (_21420_, _21419_, _21408_);
  and (_21421_, _21420_, _21417_);
  or (_21422_, _21421_, _21416_);
  and (_21423_, _21422_, _20650_);
  or (_21424_, _21412_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_21425_, _21412_, _20689_);
  and (_21426_, _21425_, _21409_);
  and (_21427_, _21426_, _21424_);
  or (_21428_, _21412_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_21429_, \oc8051_symbolic_cxrom1.regvalid [12], _26025_);
  nor (_21430_, _21429_, _21409_);
  and (_21431_, _21430_, _21428_);
  or (_21432_, _21431_, _21427_);
  and (_21433_, _21432_, _20701_);
  or (_21434_, _21433_, _21423_);
  and (_21435_, _21412_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_21436_, _21412_, _20707_);
  or (_21437_, _21436_, _21435_);
  and (_21438_, _21437_, _21409_);
  or (_21439_, _21412_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_21440_, _04993_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_21441_, _21440_);
  and (_21442_, _21441_, _21408_);
  and (_21443_, _21442_, _21439_);
  or (_21444_, _21443_, _21438_);
  and (_21445_, _21444_, _20659_);
  and (_21446_, _21412_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_21447_, _21412_, _04941_);
  or (_21448_, _21447_, _21446_);
  and (_21449_, _21448_, _21409_);
  or (_21450_, _21412_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_21451_, _04950_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21452_, _21451_, _21409_);
  and (_21453_, _21452_, _21450_);
  or (_21454_, _21453_, _21449_);
  and (_21455_, _21454_, _20674_);
  or (_21456_, _21455_, _21445_);
  or (_21457_, _21456_, _21434_);
  or (_21458_, \oc8051_symbolic_cxrom1.regvalid [0], _26025_);
  or (_21459_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_21460_, _21459_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_21461_, _21460_, _21458_);
  and (_21462_, _21461_, _20674_);
  and (_21463_, _04968_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21464_, _21463_, _26021_);
  and (_21465_, _21464_, _21419_);
  and (_21466_, _20677_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21467_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21468_, _21467_, _21466_);
  and (_21469_, _21468_, _26021_);
  nor (_21470_, _21469_, _21465_);
  nor (_21471_, _21470_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21472_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21473_, _21472_, _21451_);
  and (_21474_, _21473_, _20653_);
  or (_21475_, _21474_, _21471_);
  and (_21476_, _21475_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21477_, _21476_, _21462_);
  and (_21478_, _04941_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21479_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21480_, _21479_, _21478_);
  and (_21481_, _21480_, _20660_);
  nor (_21482_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21483_, _21482_, _26021_);
  and (_21484_, _21483_, _21441_);
  and (_21485_, _05656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21486_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21487_, _21486_, _21485_);
  and (_21488_, _21487_, _26021_);
  nor (_21489_, _21488_, _21484_);
  nor (_21490_, _21489_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21491_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21492_, _21491_, _21429_);
  and (_21493_, _21492_, _20653_);
  or (_21494_, _21493_, _21490_);
  and (_21495_, _21494_, _26013_);
  nor (_21496_, _21495_, _21481_);
  and (_21497_, _21496_, _21477_);
  nor (_21498_, _21489_, _26017_);
  nor (_21499_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21500_, _20689_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21501_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21502_, _21501_, _21500_);
  and (_21503_, _21502_, _21499_);
  and (_21504_, _21492_, _20652_);
  or (_21505_, _21504_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_21506_, _21505_, _21503_);
  nor (_21507_, _21506_, _21498_);
  nor (_21508_, _21470_, _26017_);
  and (_21509_, _05592_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21510_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21511_, _21510_, _21509_);
  and (_21512_, _21511_, _21499_);
  and (_21513_, _21473_, _20652_);
  or (_21514_, _21513_, _26013_);
  or (_21515_, _21514_, _21512_);
  nor (_21516_, _21515_, _21508_);
  nor (_21517_, _21516_, _21507_);
  not (_21518_, _25943_);
  nor (_21519_, _21518_, first_instr);
  nand (_21520_, _21519_, _21517_);
  or (_21521_, _21520_, _21497_);
  nor (_21522_, _21521_, _20715_);
  and (_21523_, _21522_, _21457_);
  and (_21524_, _21523_, _21405_);
  nor (_21525_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21526_, _07872_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21527_, _21526_, _21525_);
  and (_21528_, _21527_, _20635_);
  nor (_21529_, _21528_, _26025_);
  nor (_21530_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21531_, _07116_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21532_, _21531_, _21530_);
  and (_21533_, _21532_, _21499_);
  not (_21534_, _21533_);
  nor (_21535_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21536_, _07388_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21537_, _21536_, _21535_);
  and (_21538_, _21537_, _20653_);
  nor (_21539_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21540_, _07654_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21541_, _21540_, _21539_);
  and (_21542_, _21541_, _20652_);
  nor (_21543_, _21542_, _21538_);
  and (_21544_, _21543_, _21534_);
  and (_21545_, _21544_, _21529_);
  nor (_21546_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21547_, _06822_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21548_, _21547_, _21546_);
  and (_21549_, _21548_, _20635_);
  nor (_21550_, _21549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21551_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21552_, _06009_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21553_, _21552_, _21551_);
  and (_21554_, _21553_, _21499_);
  not (_21555_, _21554_);
  nor (_21556_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21557_, _06255_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21558_, _21557_, _21556_);
  and (_21559_, _21558_, _20653_);
  nor (_21560_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21561_, _06532_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21562_, _21561_, _21560_);
  and (_21563_, _21562_, _20652_);
  nor (_21564_, _21563_, _21559_);
  and (_21565_, _21564_, _21555_);
  and (_21566_, _21565_, _21550_);
  nor (_21567_, _21566_, _21545_);
  and (_21568_, _21567_, _21517_);
  nor (_21569_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21570_, _06269_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21571_, _21570_, _21569_);
  and (_21572_, _21571_, _20653_);
  nor (_21573_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21574_, _06554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21575_, _21574_, _21573_);
  and (_21576_, _21575_, _20652_);
  nor (_21577_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21578_, _06020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21579_, _21578_, _21577_);
  and (_21580_, _21579_, _21499_);
  nor (_21581_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21582_, _06840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21583_, _21582_, _21581_);
  and (_21584_, _21583_, _20635_);
  or (_21585_, _21584_, _21580_);
  or (_21586_, _21585_, _21576_);
  or (_21587_, _21586_, _21572_);
  and (_21588_, _21587_, _26025_);
  nor (_21589_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21590_, _07413_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21591_, _21590_, _21589_);
  and (_21592_, _21591_, _20653_);
  nor (_21593_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21594_, _07668_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21595_, _21594_, _21593_);
  and (_21596_, _21595_, _20652_);
  nor (_21597_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21598_, _07126_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21599_, _21598_, _21597_);
  and (_21600_, _21599_, _21499_);
  nor (_21601_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21602_, _07885_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21603_, _21602_, _21601_);
  and (_21604_, _21603_, _20635_);
  or (_21605_, _21604_, _21600_);
  or (_21606_, _21605_, _21596_);
  or (_21607_, _21606_, _21592_);
  and (_21608_, _21607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21609_, _21608_, _21588_);
  and (_21610_, _21609_, _21517_);
  nor (_21611_, _21610_, _21568_);
  nor (_21612_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21613_, _06299_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21614_, _21613_, _21612_);
  and (_21615_, _21614_, _20653_);
  nor (_21616_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21617_, _06590_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21618_, _21617_, _21616_);
  and (_21619_, _21618_, _20652_);
  nor (_21620_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21621_, _06048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21622_, _21621_, _21620_);
  and (_21623_, _21622_, _21499_);
  nor (_21624_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21625_, _06869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21626_, _21625_, _21624_);
  and (_21627_, _21626_, _20635_);
  or (_21628_, _21627_, _21623_);
  or (_21629_, _21628_, _21619_);
  or (_21630_, _21629_, _21615_);
  and (_21631_, _21630_, _26025_);
  nor (_21632_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21633_, _07444_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21634_, _21633_, _21632_);
  and (_21635_, _21634_, _20653_);
  nor (_21636_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21637_, _07693_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21638_, _21637_, _21636_);
  and (_21639_, _21638_, _20652_);
  nor (_21640_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21641_, _07158_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21642_, _21641_, _21640_);
  and (_21643_, _21642_, _21499_);
  nor (_21644_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21645_, _07916_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21646_, _21645_, _21644_);
  and (_21647_, _21646_, _20635_);
  or (_21648_, _21647_, _21643_);
  or (_21649_, _21648_, _21639_);
  or (_21650_, _21649_, _21635_);
  and (_21651_, _21650_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21652_, _21651_, _21631_);
  and (_21653_, _21652_, _21517_);
  nor (_21654_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21655_, _06281_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21656_, _21655_, _21654_);
  and (_21657_, _21656_, _20653_);
  nor (_21658_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21659_, _06572_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21661_, _21659_, _21658_);
  and (_21662_, _21661_, _20652_);
  nor (_21663_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21664_, _06036_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21665_, _21664_, _21663_);
  and (_21666_, _21665_, _21499_);
  nor (_21667_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21668_, _06857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21669_, _21668_, _21667_);
  and (_21670_, _21669_, _20635_);
  or (_21671_, _21670_, _21666_);
  or (_21672_, _21671_, _21662_);
  or (_21673_, _21672_, _21657_);
  and (_21674_, _21673_, _26025_);
  nor (_21675_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21676_, _07430_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21677_, _21676_, _21675_);
  and (_21678_, _21677_, _20653_);
  nor (_21679_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21680_, _07681_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21681_, _21680_, _21679_);
  and (_21682_, _21681_, _20652_);
  nor (_21683_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21684_, _07143_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21685_, _21684_, _21683_);
  and (_21686_, _21685_, _21499_);
  nor (_21687_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21688_, _07898_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21689_, _21688_, _21687_);
  and (_21690_, _21689_, _20635_);
  or (_21691_, _21690_, _21686_);
  or (_21692_, _21691_, _21682_);
  or (_21693_, _21692_, _21678_);
  and (_21694_, _21693_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21695_, _21694_, _21674_);
  and (_21696_, _21695_, _21517_);
  nor (_21697_, _21696_, _21653_);
  and (_21698_, _21697_, _21611_);
  nor (_21699_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21700_, _06078_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21701_, _21700_, _21699_);
  and (_21702_, _21701_, _21499_);
  nor (_21703_, _21702_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21704_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21705_, _06621_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21706_, _21705_, _21704_);
  and (_21707_, _21706_, _20652_);
  not (_21708_, _21707_);
  nor (_21709_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21710_, _06325_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21711_, _21710_, _21709_);
  and (_21712_, _21711_, _20653_);
  nor (_21713_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21714_, _06903_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21715_, _21714_, _21713_);
  and (_21716_, _21715_, _20635_);
  nor (_21717_, _21716_, _21712_);
  and (_21718_, _21717_, _21708_);
  and (_21719_, _21718_, _21703_);
  nor (_21720_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21721_, _07188_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21722_, _21721_, _21720_);
  and (_21723_, _21722_, _21499_);
  nor (_21724_, _21723_, _26025_);
  nor (_21725_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21726_, _07719_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21727_, _21726_, _21725_);
  and (_21728_, _21727_, _20652_);
  not (_21729_, _21728_);
  nor (_21730_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21731_, _07475_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21732_, _21731_, _21730_);
  and (_21733_, _21732_, _20653_);
  nor (_21734_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21735_, _07950_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21736_, _21735_, _21734_);
  and (_21737_, _21736_, _20635_);
  nor (_21738_, _21737_, _21733_);
  and (_21739_, _21738_, _21729_);
  and (_21740_, _21739_, _21724_);
  nor (_21741_, _21740_, _21719_);
  and (_21742_, _21741_, _21517_);
  nor (_21743_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21744_, _07931_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21745_, _21744_, _21743_);
  and (_21746_, _21745_, _20635_);
  nor (_21747_, _21746_, _26025_);
  nor (_21748_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21749_, _07172_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21750_, _21749_, _21748_);
  and (_21751_, _21750_, _21499_);
  not (_21752_, _21751_);
  nor (_21753_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21754_, _07457_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21755_, _21754_, _21753_);
  and (_21756_, _21755_, _20653_);
  nor (_21757_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21758_, _07705_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21759_, _21758_, _21757_);
  and (_21760_, _21759_, _20652_);
  nor (_21761_, _21760_, _21756_);
  and (_21762_, _21761_, _21752_);
  and (_21763_, _21762_, _21747_);
  nor (_21764_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21765_, _06885_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21766_, _21765_, _21764_);
  and (_21767_, _21766_, _20635_);
  nor (_21768_, _21767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21769_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21770_, _06063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21771_, _21770_, _21769_);
  and (_21772_, _21771_, _21499_);
  not (_21773_, _21772_);
  nor (_21774_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21775_, _06312_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21776_, _21775_, _21774_);
  and (_21777_, _21776_, _20653_);
  nor (_21778_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21779_, _06606_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21780_, _21779_, _21778_);
  and (_21781_, _21780_, _20652_);
  nor (_21782_, _21781_, _21777_);
  and (_21783_, _21782_, _21773_);
  and (_21784_, _21783_, _21768_);
  nor (_21785_, _21784_, _21763_);
  and (_21786_, _21785_, _21517_);
  nor (_21787_, _21786_, _21742_);
  not (_21788_, _21517_);
  nor (_21789_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21790_, _05006_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21791_, _21790_, _21789_);
  nand (_21792_, _21791_, _20635_);
  and (_21793_, _21792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_21794_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21795_, _05023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21796_, _21795_, _21794_);
  nand (_21797_, _21796_, _21499_);
  nor (_21798_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21799_, _05011_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21800_, _21799_, _21798_);
  nand (_21801_, _21800_, _20653_);
  nor (_21802_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21803_, _05018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21804_, _21803_, _21802_);
  nand (_21805_, _21804_, _20652_);
  and (_21806_, _21805_, _21801_);
  and (_21807_, _21806_, _21797_);
  and (_21808_, _21807_, _21793_);
  nor (_21809_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21810_, _05045_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21811_, _21810_, _21809_);
  nand (_21812_, _21811_, _20635_);
  and (_21813_, _21812_, _26025_);
  nor (_21814_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21815_, _05036_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21816_, _21815_, _21814_);
  nand (_21817_, _21816_, _21499_);
  nor (_21818_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21819_, _05051_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21820_, _21819_, _21818_);
  nand (_21821_, _21820_, _20653_);
  nor (_21822_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21823_, _05031_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21824_, _21823_, _21822_);
  nand (_21825_, _21824_, _20652_);
  and (_21826_, _21825_, _21821_);
  and (_21827_, _21826_, _21817_);
  and (_21828_, _21827_, _21813_);
  or (_21829_, _21828_, _21808_);
  nor (_21830_, _21829_, _21788_);
  nor (_21831_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21832_, _06338_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21833_, _21832_, _21831_);
  and (_21834_, _21833_, _20653_);
  nor (_21835_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21836_, _06636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21837_, _21836_, _21835_);
  and (_21838_, _21837_, _20652_);
  nor (_21839_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21840_, _06091_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21841_, _21840_, _21839_);
  and (_21842_, _21841_, _21499_);
  nor (_21843_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21844_, _06918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21845_, _21844_, _21843_);
  and (_21846_, _21845_, _20635_);
  or (_21847_, _21846_, _21842_);
  or (_21848_, _21847_, _21838_);
  or (_21849_, _21848_, _21834_);
  and (_21850_, _21849_, _26025_);
  nor (_21851_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21852_, _07492_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21853_, _21852_, _21851_);
  and (_21854_, _21853_, _20653_);
  nor (_21855_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21856_, _07734_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21857_, _21856_, _21855_);
  and (_21858_, _21857_, _20652_);
  nor (_21859_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21860_, _07204_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21861_, _21860_, _21859_);
  and (_21862_, _21861_, _21499_);
  nor (_21863_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21864_, _07963_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_21865_, _21864_, _21863_);
  and (_21866_, _21865_, _20635_);
  or (_21867_, _21866_, _21862_);
  or (_21868_, _21867_, _21858_);
  or (_21869_, _21868_, _21854_);
  and (_21870_, _21869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_21871_, _21870_, _21850_);
  and (_21872_, _21871_, _21517_);
  not (_21873_, _21872_);
  and (_21874_, _21873_, _21830_);
  and (_21875_, _21874_, _21787_);
  and (_21876_, _21875_, _21698_);
  and (_21877_, _21876_, _21524_);
  and (_21878_, _21877_, _21253_);
  not (_21879_, _21830_);
  and (_21880_, _21696_, _21610_);
  and (_21881_, _21880_, _21786_);
  and (_21882_, _21881_, _21742_);
  not (_21883_, _21568_);
  and (_21884_, _21697_, _21883_);
  and (_21885_, _21884_, _21610_);
  not (_21886_, _21567_);
  nor (_21887_, _21652_, _21609_);
  and (_21888_, _21887_, _21696_);
  and (_21889_, _21888_, _21886_);
  and (_21890_, _21652_, _21742_);
  and (_21891_, _21890_, _21786_);
  or (_21892_, _21891_, _21889_);
  or (_21893_, _21892_, _21885_);
  or (_21894_, _21893_, _21882_);
  and (_21895_, _21894_, _21872_);
  not (_21896_, _21742_);
  nor (_21897_, _21871_, _21896_);
  and (_21898_, _21897_, _21888_);
  and (_21899_, _21888_, _21568_);
  and (_21900_, _21899_, _21896_);
  or (_21901_, _21900_, _21898_);
  or (_21902_, _21901_, _21895_);
  and (_21903_, _21902_, _21879_);
  and (_21904_, _21884_, _21741_);
  not (_21905_, _21741_);
  and (_21906_, _21786_, _21905_);
  and (_21907_, _21906_, _21888_);
  not (_21908_, _21785_);
  and (_21909_, _21653_, _21908_);
  not (_21910_, _21786_);
  and (_21911_, _21880_, _21910_);
  or (_21912_, _21911_, _21909_);
  or (_21913_, _21912_, _21907_);
  or (_21914_, _21913_, _21904_);
  and (_21915_, _21914_, _21874_);
  and (_21916_, _21872_, _21908_);
  and (_21917_, _21916_, _21899_);
  and (_21918_, _21885_, _21896_);
  and (_21919_, _21872_, _21905_);
  and (_21920_, _21919_, _21884_);
  and (_21921_, _21872_, _21741_);
  and (_21922_, _21921_, _21899_);
  or (_21923_, _21922_, _21920_);
  or (_21924_, _21923_, _21918_);
  and (_21925_, _21924_, _21830_);
  or (_21926_, _21925_, _21917_);
  or (_21927_, _21926_, _21915_);
  or (_21928_, _21927_, _21903_);
  nor (_21929_, _20762_, _26001_);
  and (_21930_, _20762_, _26001_);
  or (_21931_, _21930_, _21929_);
  or (_21932_, _21931_, _21152_);
  and (_21933_, _20649_, _26009_);
  nor (_21934_, _20649_, _26009_);
  or (_21935_, _21934_, _21933_);
  or (_21936_, _21935_, _21137_);
  or (_21937_, _21936_, _21932_);
  nor (_21938_, _20795_, _25971_);
  and (_21939_, _20795_, _25971_);
  or (_21940_, _21939_, _21938_);
  and (_21941_, _20784_, _25981_);
  or (_21942_, _21941_, _21940_);
  nor (_21943_, _20840_, _25966_);
  and (_21944_, _20789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_21945_, _21944_, _21943_);
  and (_21946_, _20840_, _25966_);
  nor (_21947_, _20789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_21948_, _21947_, _21946_);
  or (_21949_, _21948_, _21945_);
  and (_21950_, _20925_, _25958_);
  nor (_21951_, _20925_, _25958_);
  or (_21952_, _21951_, _21950_);
  nor (_21953_, _20654_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21954_, _20654_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21955_, _21954_, _21953_);
  and (_21956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_21957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_21958_, _21957_, _21956_);
  nand (_21959_, _21958_, _21219_);
  or (_21960_, _21959_, _21955_);
  or (_21961_, _21960_, _21952_);
  and (_21962_, _20922_, _25962_);
  nor (_21963_, _20922_, _25962_);
  or (_21964_, _21963_, _21962_);
  or (_21965_, _21964_, _21961_);
  nor (_21966_, _20784_, _25981_);
  or (_21967_, _21966_, _21965_);
  or (_21968_, _21967_, _21949_);
  or (_21969_, _21968_, _21942_);
  nor (_21970_, _20775_, _25990_);
  and (_21971_, _20775_, _25990_);
  or (_21972_, _21971_, _21970_);
  or (_21973_, _21186_, _21166_);
  or (_21974_, _21973_, _21972_);
  or (_21975_, _21974_, _21969_);
  or (_21976_, _21975_, _21937_);
  and (_21977_, _21976_, _21928_);
  nor (_21978_, _21872_, _21830_);
  and (_21979_, _21787_, _21611_);
  and (_21980_, _21696_, _21886_);
  and (_21982_, _21980_, _21896_);
  or (_21983_, _21982_, _21979_);
  and (_21984_, _21983_, _21978_);
  and (_21985_, _21609_, _21568_);
  nor (_21986_, _21879_, _21652_);
  and (_21987_, _21986_, _21985_);
  or (_21988_, _21987_, _21911_);
  and (_21989_, _21988_, _21872_);
  and (_21990_, _21873_, _21653_);
  or (_21991_, _21906_, _21829_);
  and (_21992_, _21991_, _21990_);
  and (_21993_, _21909_, _21872_);
  and (_21994_, _21978_, _21880_);
  or (_21995_, _21994_, _21993_);
  or (_21996_, _21995_, _21992_);
  or (_21997_, _21996_, _21989_);
  or (_21998_, _21997_, _21984_);
  and (_21999_, _21985_, _21697_);
  and (_22000_, _21889_, _21787_);
  or (_22001_, _22000_, _21999_);
  and (_22002_, _22001_, _21873_);
  and (_22003_, _21898_, _21910_);
  not (_22004_, _21652_);
  and (_22005_, _21696_, _22004_);
  or (_22006_, _22005_, _21742_);
  or (_22007_, _21652_, _21886_);
  and (_22008_, _22007_, _21872_);
  and (_22009_, _22008_, _22006_);
  or (_22010_, _22009_, _22003_);
  and (_22011_, _22010_, _21830_);
  nand (_22012_, _21829_, _21905_);
  nand (_22013_, _22012_, _21653_);
  and (_22014_, _21881_, _21896_);
  or (_22015_, _22014_, _21653_);
  and (_22016_, _22015_, _22013_);
  or (_22017_, _22016_, _22011_);
  or (_22018_, _22017_, _22002_);
  or (_22019_, _22018_, _21998_);
  and (_22020_, _20769_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26013_);
  nor (_22022_, _22021_, _22020_);
  and (_22023_, _22022_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22024_, _20786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22026_, _22025_, _22024_);
  nor (_22027_, _22026_, _20794_);
  and (_22028_, _22027_, _25971_);
  or (_22029_, _22028_, _22023_);
  and (_22030_, _20662_, _20639_);
  nor (_22031_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_22032_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_22033_, _22032_, _22031_);
  and (_22034_, _22033_, _22030_);
  nor (_22035_, _22033_, _22030_);
  or (_22036_, _22035_, _22034_);
  or (_22037_, _20758_, _26013_);
  or (_22038_, _26063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22039_, _22038_, _22037_);
  and (_22040_, _22039_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22041_, _22022_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_22042_, _22041_, _22040_);
  or (_22043_, _22042_, _22036_);
  or (_22044_, _22043_, _22029_);
  and (_22045_, _22030_, _20643_);
  and (_22046_, _22045_, _20645_);
  and (_22047_, _22046_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_22048_, _22047_, _20632_);
  nor (_22049_, _22047_, _20632_);
  nor (_22050_, _22049_, _22048_);
  and (_22051_, _22050_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_22052_, _22030_, _20641_);
  and (_22053_, _22052_, _26052_);
  nor (_22054_, _22052_, _26052_);
  or (_22055_, _22054_, _22053_);
  and (_22056_, _22055_, _25990_);
  or (_22057_, _22056_, _22051_);
  nor (_22058_, _22050_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_22059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_22060_, _22045_, _22059_);
  nor (_22061_, _22045_, _22059_);
  or (_22062_, _22061_, _22060_);
  and (_22063_, _22062_, _26001_);
  nor (_22064_, _22062_, _26001_);
  or (_22065_, _22064_, _22063_);
  or (_22066_, _22065_, _22058_);
  or (_22067_, _22066_, _22057_);
  nor (_22068_, _22039_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22069_, _22046_, _26068_);
  nor (_22070_, _22046_, _26068_);
  or (_22071_, _22070_, _22069_);
  and (_22072_, _22071_, _26009_);
  nor (_22073_, _22071_, _26009_);
  or (_22074_, _22073_, _22072_);
  or (_22075_, _22074_, _22068_);
  or (_22076_, _26048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22077_, _20780_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22078_, _22077_, _22076_);
  nor (_22079_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22080_, _22078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_22081_, _22024_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22082_, _22081_, _22030_);
  and (_22083_, _22082_, _25976_);
  or (_22084_, _22083_, _22080_);
  or (_22085_, _22084_, _22079_);
  nor (_22086_, _22055_, _25990_);
  nor (_22087_, _20663_, _25958_);
  and (_22088_, _20663_, _25958_);
  or (_22089_, _22088_, _22087_);
  nor (_22090_, _22082_, _25976_);
  nor (_22091_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_22092_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_22093_, _22092_, _22091_);
  nand (_22094_, _22093_, _20662_);
  or (_22095_, _22093_, _20662_);
  and (_22096_, _22095_, _22094_);
  or (_22097_, _22096_, _22090_);
  nor (_22098_, _20657_, _25953_);
  and (_22099_, _20657_, _25953_);
  or (_22100_, _22099_, _22098_);
  or (_22101_, _26032_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_22102_, _20840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22103_, _22102_, _22101_);
  and (_22104_, _22103_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22105_, _21958_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_22106_, _21958_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_22107_, _22106_, _22105_);
  or (_22108_, _22107_, _21219_);
  or (_22109_, _22108_, _22104_);
  or (_22110_, _22109_, _22100_);
  nor (_22111_, _22103_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_22112_, _22027_, _25971_);
  or (_22113_, _22112_, _22111_);
  or (_22114_, _22113_, _22110_);
  or (_22115_, _22114_, _22097_);
  or (_22116_, _22115_, _22089_);
  or (_22117_, _22116_, _22086_);
  or (_22118_, _22117_, _22085_);
  or (_22119_, _22118_, _22075_);
  or (_22120_, _22119_, _22067_);
  or (_22121_, _22120_, _22044_);
  and (_22122_, _22121_, _22019_);
  and (_22123_, _21906_, _21698_);
  and (_22124_, _21900_, _21908_);
  or (_22125_, _22124_, _22123_);
  and (_22126_, _22125_, _21874_);
  and (_22127_, _21922_, _21786_);
  or (_22128_, _21919_, _21916_);
  and (_22129_, _22128_, _21999_);
  or (_22130_, _22129_, _22127_);
  and (_22131_, _22130_, _21879_);
  or (_22132_, _22131_, _22126_);
  and (_22133_, _21410_, _20639_);
  and (_22134_, _22133_, _20643_);
  and (_22135_, _22134_, _20645_);
  and (_22136_, _22135_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_22137_, _22136_, _20632_);
  nor (_22138_, _22136_, _20632_);
  nor (_22139_, _22138_, _22137_);
  nor (_22140_, _22139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_22141_, _22133_, _20641_);
  and (_22142_, _22141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22143_, _22141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_22144_, _22143_, _22142_);
  and (_22145_, _22144_, _25990_);
  or (_22146_, _22145_, _22140_);
  and (_22147_, _22134_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_22148_, _22147_, _26063_);
  and (_22149_, _22147_, _26063_);
  nor (_22150_, _22149_, _22148_);
  and (_22151_, _22150_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22152_, _21410_, _20638_);
  and (_22153_, _21410_, _20637_);
  nor (_22154_, _22153_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_22155_, _22154_, _22152_);
  and (_22156_, _22155_, _25971_);
  and (_22157_, _22142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22158_, _22142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_22159_, _22158_, _22157_);
  nor (_22160_, _22159_, _25996_);
  and (_22161_, _22133_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22162_, _22133_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_22163_, _22162_, _22161_);
  nor (_22164_, _22163_, _25981_);
  and (_22165_, _22163_, _25981_);
  or (_22166_, _22165_, _22164_);
  or (_22167_, _22166_, _22160_);
  or (_22168_, _22167_, _22156_);
  or (_22169_, _22168_, _22151_);
  and (_22170_, _22159_, _25996_);
  nor (_22171_, _22161_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22172_, _22171_, _22141_);
  and (_22173_, _22172_, _25985_);
  nor (_22174_, _22172_, _25985_);
  or (_22175_, _22174_, _22173_);
  nor (_22176_, _22144_, _25990_);
  nor (_22177_, _22152_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22178_, _22177_, _22133_);
  and (_22179_, _22178_, _25976_);
  or (_22180_, _22179_, _22176_);
  or (_22181_, _22180_, _22175_);
  or (_22182_, _22093_, _21410_);
  nand (_22183_, _22093_, _21410_);
  and (_22184_, _22183_, _22182_);
  and (_22185_, _21410_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_22186_, _22185_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_22187_, _22186_, _22153_);
  nor (_22188_, _22187_, _25966_);
  or (_22189_, _21408_, _25953_);
  nand (_22190_, _22189_, _22107_);
  and (_22191_, _21408_, _25953_);
  or (_22192_, _22191_, _21219_);
  or (_22193_, _22192_, _22190_);
  or (_22194_, _22193_, _22188_);
  nor (_22195_, _22155_, _25971_);
  and (_22196_, _22187_, _25966_);
  or (_22197_, _22196_, _22195_);
  nor (_22198_, _22178_, _25976_);
  or (_22199_, _21412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22200_, _21412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22201_, _22200_, _22199_);
  or (_22202_, _22201_, _22198_);
  or (_22203_, _22202_, _22197_);
  or (_22204_, _22203_, _22194_);
  or (_22205_, _22204_, _22184_);
  or (_22206_, _22205_, _22181_);
  or (_22207_, _22206_, _22170_);
  or (_22208_, _22207_, _22169_);
  or (_22209_, _22208_, _22146_);
  nor (_22210_, _22150_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_22211_, _22135_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_22212_, _22211_, _22136_);
  and (_22213_, _22212_, _26009_);
  nor (_22214_, _22212_, _26009_);
  or (_22215_, _22214_, _22213_);
  or (_22216_, _22215_, _22210_);
  and (_22217_, _22134_, _22059_);
  nor (_22218_, _22134_, _22059_);
  or (_22219_, _22218_, _22217_);
  nand (_22220_, _22219_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_22221_, _22219_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_22222_, _22221_, _22220_);
  and (_22223_, _22139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_22224_, _22223_, _22222_);
  or (_22225_, _22224_, _22216_);
  or (_22226_, _22225_, _22209_);
  and (_22227_, _22226_, _22132_);
  or (_22228_, _22227_, _22122_);
  or (_22229_, _22228_, _21977_);
  and (_22230_, _22229_, _21524_);
  not (_22231_, _21497_);
  and (_22233_, _21634_, _21499_);
  and (_22234_, _21646_, _20652_);
  and (_22235_, _21642_, _20635_);
  and (_22236_, _21638_, _20653_);
  or (_22237_, _22236_, _22235_);
  or (_22238_, _22237_, _22234_);
  or (_22239_, _22238_, _22233_);
  and (_22240_, _22239_, _20925_);
  not (_22241_, _20925_);
  and (_22242_, _21614_, _21499_);
  and (_22243_, _21626_, _20652_);
  and (_22244_, _21622_, _20635_);
  and (_22245_, _21618_, _20653_);
  or (_22246_, _22245_, _22244_);
  or (_22247_, _22246_, _22243_);
  or (_22248_, _22247_, _22242_);
  and (_22249_, _22248_, _22241_);
  or (_22250_, _22249_, _22240_);
  and (_22251_, _22250_, _22231_);
  nand (_22252_, _22251_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_22254_, _22251_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22255_, _22254_, _22252_);
  and (_22256_, _21677_, _21499_);
  and (_22257_, _21689_, _20652_);
  and (_22258_, _21685_, _20635_);
  and (_22259_, _21681_, _20653_);
  or (_22260_, _22259_, _22258_);
  or (_22261_, _22260_, _22257_);
  or (_22262_, _22261_, _22256_);
  and (_22263_, _22262_, _20925_);
  and (_22264_, _21656_, _21499_);
  and (_22265_, _21669_, _20652_);
  and (_22266_, _21665_, _20635_);
  and (_22267_, _21661_, _20653_);
  or (_22268_, _22267_, _22266_);
  or (_22269_, _22268_, _22265_);
  or (_22270_, _22269_, _22264_);
  and (_22271_, _22270_, _22241_);
  or (_22272_, _22271_, _22263_);
  and (_22273_, _22272_, _22231_);
  and (_22274_, _22273_, _25953_);
  nor (_22275_, _22273_, _25953_);
  or (_22276_, _22275_, _22274_);
  or (_22277_, _22276_, _22255_);
  and (_22278_, _21562_, _20653_);
  and (_22279_, _21548_, _20652_);
  and (_22280_, _21553_, _20635_);
  or (_22281_, _22280_, _22279_);
  or (_22282_, _22281_, _22278_);
  and (_22283_, _21558_, _21499_);
  or (_22284_, _22283_, _20925_);
  or (_22285_, _22284_, _22282_);
  and (_22286_, _21541_, _20653_);
  or (_22287_, _22286_, _22241_);
  and (_22288_, _21532_, _20635_);
  and (_22289_, _21537_, _21499_);
  and (_22290_, _21527_, _20652_);
  or (_22291_, _22290_, _22289_);
  or (_22292_, _22291_, _22288_);
  or (_22293_, _22292_, _22287_);
  nand (_22294_, _22293_, _22285_);
  nor (_22295_, _22294_, _21497_);
  and (_22296_, _22295_, _25945_);
  nor (_22297_, _22295_, _25945_);
  or (_22298_, _22297_, _22296_);
  and (_22299_, _21591_, _21499_);
  and (_22300_, _21603_, _20652_);
  and (_22301_, _21599_, _20635_);
  and (_22302_, _21595_, _20653_);
  or (_22303_, _22302_, _22301_);
  or (_22304_, _22303_, _22300_);
  or (_22305_, _22304_, _22299_);
  and (_22306_, _22305_, _20925_);
  and (_22307_, _21571_, _21499_);
  and (_22308_, _21583_, _20652_);
  and (_22309_, _21575_, _20653_);
  and (_22310_, _21579_, _20635_);
  or (_22311_, _22310_, _22309_);
  or (_22312_, _22311_, _22308_);
  or (_22313_, _22312_, _22307_);
  and (_22314_, _22313_, _22241_);
  or (_22315_, _22314_, _22306_);
  and (_22316_, _22315_, _22231_);
  and (_22317_, _22316_, _25949_);
  nor (_22318_, _22316_, _25949_);
  or (_22319_, _22318_, _22317_);
  or (_22320_, _22319_, _22298_);
  or (_22321_, _22320_, _22277_);
  and (_22322_, _21837_, _20653_);
  nor (_22323_, _22322_, _20925_);
  and (_22324_, _21841_, _20635_);
  and (_22325_, _21833_, _21499_);
  nor (_22326_, _22325_, _22324_);
  and (_22327_, _21845_, _20652_);
  not (_22328_, _22327_);
  and (_22329_, _22328_, _22326_);
  and (_22330_, _22329_, _22323_);
  and (_22331_, _21865_, _20652_);
  and (_22332_, _21857_, _20653_);
  and (_22333_, _21861_, _20635_);
  or (_22334_, _22333_, _22332_);
  nor (_22335_, _22334_, _22331_);
  and (_22336_, _21853_, _21499_);
  nor (_22337_, _22336_, _22241_);
  and (_22338_, _22337_, _22335_);
  nor (_22339_, _22338_, _22330_);
  and (_22340_, _22339_, _22231_);
  nand (_22341_, _22340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_22342_, _22340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_22343_, _22342_, _22341_);
  and (_22344_, _21791_, _20652_);
  and (_22345_, _21804_, _20653_);
  nor (_22346_, _22345_, _22344_);
  and (_22347_, _21796_, _20635_);
  and (_22348_, _21800_, _21499_);
  nor (_22349_, _22348_, _22347_);
  and (_22350_, _22349_, _22346_);
  and (_22351_, _22350_, _20925_);
  and (_22352_, _21816_, _20635_);
  not (_22353_, _22352_);
  and (_22354_, _21811_, _20652_);
  and (_22355_, _21824_, _20653_);
  nor (_22356_, _22355_, _22354_);
  and (_22357_, _22356_, _22353_);
  and (_22358_, _21820_, _21499_);
  nor (_22359_, _22358_, _20925_);
  and (_22360_, _22359_, _22357_);
  nor (_22361_, _22360_, _22351_);
  and (_22362_, _22361_, _22231_);
  nor (_22363_, _22362_, _25976_);
  and (_22364_, _22362_, _25976_);
  or (_22365_, _22364_, _22363_);
  or (_22366_, _22365_, _22343_);
  and (_22367_, _21706_, _20653_);
  or (_22368_, _22367_, _20925_);
  and (_22369_, _21701_, _20635_);
  and (_22370_, _21711_, _21499_);
  and (_22371_, _21715_, _20652_);
  or (_22372_, _22371_, _22370_);
  or (_22373_, _22372_, _22369_);
  or (_22374_, _22373_, _22368_);
  and (_22375_, _21727_, _20653_);
  or (_22376_, _22375_, _22241_);
  and (_22377_, _21722_, _20635_);
  and (_22378_, _21732_, _21499_);
  and (_22379_, _21736_, _20652_);
  or (_22380_, _22379_, _22378_);
  or (_22381_, _22380_, _22377_);
  or (_22382_, _22381_, _22376_);
  nand (_22383_, _22382_, _22374_);
  nor (_22384_, _22383_, _21497_);
  nand (_22385_, _22384_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_22386_, _22384_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22387_, _22386_, _22385_);
  and (_22388_, _21780_, _20653_);
  nor (_22389_, _22388_, _20925_);
  and (_22390_, _21771_, _20635_);
  not (_22391_, _22390_);
  and (_22392_, _21776_, _21499_);
  and (_22393_, _21766_, _20652_);
  nor (_22394_, _22393_, _22392_);
  and (_22395_, _22394_, _22391_);
  and (_22396_, _22395_, _22389_);
  and (_22397_, _21745_, _20652_);
  and (_22398_, _21759_, _20653_);
  and (_22399_, _21750_, _20635_);
  or (_22400_, _22399_, _22398_);
  nor (_22401_, _22400_, _22397_);
  and (_22402_, _21755_, _21499_);
  nor (_22403_, _22402_, _22241_);
  and (_22404_, _22403_, _22401_);
  nor (_22405_, _22404_, _22396_);
  and (_22406_, _22405_, _22231_);
  nor (_22407_, _22406_, _25962_);
  and (_22408_, _22406_, _25962_);
  or (_22409_, _22408_, _22407_);
  or (_22410_, _22409_, _22387_);
  or (_22411_, _22410_, _22366_);
  or (_22412_, _22411_, _22321_);
  or (_22413_, _21045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_22414_, _21045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_22415_, _22414_, _22413_);
  nor (_22416_, _21084_, _25981_);
  and (_22417_, _21084_, _25981_);
  or (_22418_, _22417_, _22416_);
  or (_22419_, _22418_, _22415_);
  or (_22420_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_22421_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_22422_, _22421_, _22420_);
  nor (_22423_, _21006_, _25990_);
  and (_22424_, _21006_, _25990_);
  or (_22425_, _22424_, _22423_);
  or (_22426_, _22425_, _22422_);
  or (_22427_, _22426_, _22419_);
  and (_22428_, _20920_, _26001_);
  nor (_22429_, _20920_, _26001_);
  or (_22430_, _22429_, _22428_);
  or (_22431_, _20878_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_22432_, _20878_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_22433_, _22432_, _22431_);
  or (_22434_, _22433_, _22430_);
  nor (_22435_, _20753_, _14355_);
  and (_22436_, _20753_, _14355_);
  or (_22437_, _22436_, _22435_);
  nor (_22438_, _20833_, _26009_);
  and (_22439_, _20833_, _26009_);
  or (_22440_, _22439_, _22438_);
  or (_22441_, _22440_, _22437_);
  or (_22442_, _22441_, _22434_);
  or (_22443_, _22442_, _22427_);
  or (_22444_, _22443_, _22412_);
  and (_22445_, _21978_, _21918_);
  and (_22446_, _22445_, _21524_);
  and (_22447_, _22446_, _22444_);
  nor (_22448_, _21742_, _25981_);
  and (_22449_, _21742_, _25981_);
  or (_22450_, _22449_, _22448_);
  and (_22451_, _21872_, _25985_);
  nor (_22452_, _21872_, _25985_);
  or (_22453_, _22452_, _22451_);
  or (_22454_, _22453_, _22450_);
  nor (_22455_, _21830_, _25990_);
  and (_22456_, _21830_, _25990_);
  or (_22457_, _22456_, _22455_);
  or (_22458_, _22457_, _21166_);
  or (_22459_, _22458_, _22454_);
  or (_22460_, _22459_, _21937_);
  or (_22461_, _21045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_22462_, _21045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_22463_, _22462_, _22461_);
  nor (_22464_, _21084_, _25945_);
  and (_22465_, _21084_, _25945_);
  or (_22466_, _22465_, _22464_);
  or (_22467_, _22466_, _22463_);
  or (_22468_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_22469_, _20963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_22470_, _22469_, _22468_);
  and (_22471_, _21006_, _25953_);
  nor (_22472_, _21006_, _25953_);
  or (_22473_, _22472_, _22471_);
  or (_22474_, _22473_, _22470_);
  or (_22475_, _22474_, _22467_);
  or (_22476_, _20878_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22477_, _20878_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_22478_, _22477_, _22476_);
  nor (_22479_, _20920_, _25962_);
  and (_22480_, _20920_, _25962_);
  or (_22481_, _22480_, _22479_);
  or (_22482_, _22481_, _22478_);
  nor (_22483_, _20753_, _25976_);
  and (_22484_, _20753_, _25976_);
  or (_22485_, _22484_, _22483_);
  and (_22486_, _20833_, _25971_);
  nor (_22487_, _20833_, _25971_);
  or (_22488_, _22487_, _22486_);
  or (_22489_, _22488_, _22485_);
  or (_22490_, _22489_, _22482_);
  or (_22491_, _22490_, _22475_);
  or (_22492_, _22491_, _22460_);
  nor (_22493_, _21609_, _21883_);
  and (_22494_, _22493_, _21697_);
  and (_22495_, _22494_, _21524_);
  and (_22496_, _22495_, _22492_);
  or (_22497_, _22496_, _22447_);
  or (_22498_, _22497_, _22230_);
  or (property_invalid, _22498_, _21878_);
  and (_22499_, _14558_, _26242_);
  and (_22500_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_12031_, _22500_, _22499_);
  and (_22501_, _21518_, first_instr);
  or (_00000_, _22501_, rst);
  nor (_26929_[0], _24481_, rst);
  and (_22502_, _14558_, _26185_);
  and (_22503_, _14560_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_12054_, _22503_, _22502_);
  nor (_26928_[0], _24498_, rst);
  and (_22504_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_22505_, _26261_, _25886_);
  or (_12072_, _22505_, _22504_);
  nor (_26928_[6], _24262_, rst);
  and (_26892_[6], _22934_, _23049_);
  or (_22506_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_12098_, _22506_, _02890_);
  and (_22507_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  and (_22508_, _06617_, _26170_);
  or (_12104_, _22508_, _22507_);
  and (_22509_, _06618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  and (_22510_, _06617_, _25927_);
  or (_27172_, _22510_, _22509_);
  or (_22511_, _02685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_26948_, _22511_, _02900_);
  and (_22512_, _02800_, _26085_);
  and (_22513_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_27118_, _22513_, _22512_);
  and (_22514_, _02800_, _26170_);
  and (_22515_, _02802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_12133_, _22515_, _22514_);
  and (_22516_, _14639_, _25927_);
  and (_22517_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_12135_, _22517_, _22516_);
  and (_22518_, _02780_, _26170_);
  and (_22519_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_12141_, _22519_, _22518_);
  and (_22520_, _14639_, _23768_);
  and (_22521_, _14641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_12151_, _22521_, _22520_);
  and (_22522_, _02780_, _26085_);
  and (_22523_, _02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_12159_, _22523_, _22522_);
  and (_22524_, _02519_, _26185_);
  and (_22525_, _02521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_12164_, _22525_, _22524_);
  or (_22526_, _00070_, _25258_);
  nor (_22527_, _05695_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_22528_, _22527_, _05696_);
  and (_22529_, _05692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_22530_, _22529_, _22528_);
  nor (_22531_, _22530_, _00071_);
  and (_22532_, _00071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_22533_, _22532_, _22531_);
  or (_22534_, _22533_, _00069_);
  and (_22535_, _22534_, _23049_);
  and (_12166_, _22535_, _22526_);
  and (_22536_, _14991_, _25927_);
  and (_22537_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_26968_, _22537_, _22536_);
  and (_22538_, _02590_, _25886_);
  and (_22539_, _02592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_12172_, _22539_, _22538_);
  nand (_22540_, _00069_, _25279_);
  nor (_22541_, _05694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_22542_, _22541_, _05695_);
  and (_22543_, _01659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_22544_, _22543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_22545_, _01654_, _01667_);
  and (_22546_, _22545_, _22544_);
  and (_22547_, _22546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22548_, _22547_, _22542_);
  nor (_22549_, _22548_, _00071_);
  and (_22550_, _00071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_22551_, _22550_, _22549_);
  or (_22552_, _22551_, _00069_);
  and (_22553_, _22552_, _23049_);
  and (_12174_, _22553_, _22540_);
  and (_22554_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  and (_22555_, _04243_, _25927_);
  or (_12176_, _22555_, _22554_);
  and (_22556_, _14991_, _26170_);
  and (_22557_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_12197_, _22557_, _22556_);
  and (_22558_, _14629_, _26085_);
  and (_22559_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_12199_, _22559_, _22558_);
  and (_22560_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  and (_22561_, _04243_, _23768_);
  or (_12205_, _22561_, _22560_);
  and (_22562_, _14629_, _23830_);
  and (_22563_, _14631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_12208_, _22563_, _22562_);
  and (_22564_, _02570_, _26085_);
  and (_22565_, _02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_12215_, _22565_, _22564_);
  and (_22566_, _02480_, _26242_);
  and (_22567_, _02482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_12221_, _22567_, _22566_);
  and (_22568_, _14991_, _23830_);
  and (_22569_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_12228_, _22569_, _22568_);
  and (_22570_, _26262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_22571_, _26261_, _26170_);
  or (_12230_, _22571_, _22570_);
  and (_22572_, _01966_, _26170_);
  and (_22573_, _01968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_12232_, _22573_, _22572_);
  and (_22574_, _14991_, _26185_);
  and (_22575_, _14993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_12242_, _22575_, _22574_);
  and (_22576_, _00096_, _26085_);
  and (_22577_, _00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_12246_, _22577_, _22576_);
  nor (_22578_, _01654_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_22579_, _15337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22580_, _22579_, _05694_);
  or (_22581_, _22580_, _22578_);
  nor (_22582_, _22581_, _00071_);
  and (_22583_, _00071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_22584_, _22583_, _22582_);
  and (_22585_, _22584_, _00070_);
  and (_22586_, _00069_, _25283_);
  or (_22587_, _22586_, _22585_);
  and (_12248_, _22587_, _23049_);
  and (_22588_, _01564_, _26170_);
  and (_22589_, _01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_12255_, _22589_, _22588_);
  and (_22590_, _04245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  and (_22591_, _04243_, _25886_);
  or (_12261_, _22591_, _22590_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _26875_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _26875_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _26875_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _26875_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _26875_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _26875_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _26875_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _26875_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _26891_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _26874_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _26874_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _26874_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _26874_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _26874_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _26874_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _26874_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _26874_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _26874_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _26874_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _26874_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _26874_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _26874_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _26874_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _26874_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _26882_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _26882_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _26882_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _26882_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _26882_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _26882_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _26882_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _26882_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _26883_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _26883_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _26883_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _26883_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _26883_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _26883_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _26883_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _26883_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _26884_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _26884_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _26884_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _26884_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _26884_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _26884_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _26884_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _26884_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _26885_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _26885_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _26885_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _26885_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _26885_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _26885_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _26885_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _26885_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _26886_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _26886_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _26886_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _26886_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _26886_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _26886_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _26886_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _26886_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _26887_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _26887_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _26887_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _26887_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _26887_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _26887_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _26887_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _26887_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _26888_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _26888_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _26888_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _26888_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _26888_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _26888_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _26888_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _26888_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _26889_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _26889_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _26889_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _26889_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _26889_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _26889_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _26889_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _26889_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _26890_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _26890_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _26890_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _26890_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _26890_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _26890_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _26890_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _26890_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _26876_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _26876_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _26876_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _26876_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _26876_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _26876_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _26876_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _26876_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _26877_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _26877_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _26877_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _26877_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _26877_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _26877_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _26877_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _26877_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _26878_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _26878_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _26878_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _26878_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _26878_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _26878_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _26878_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _26878_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _26879_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _26879_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _26879_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _26879_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _26879_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _26879_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _26879_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _26879_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _26880_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _26880_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _26880_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _26880_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _26880_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _26880_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _26880_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _26880_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _26881_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _26881_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _26881_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _26881_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _26881_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _26881_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _26881_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _26881_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _06284_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _06282_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _06295_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _06291_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _06288_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _05609_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _06331_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _05603_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _06348_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _06351_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _06350_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _06358_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _06375_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _06381_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _06379_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _05606_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11628_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _10757_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11550_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11552_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11572_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11581_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11556_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11558_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11574_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _11561_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11563_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11576_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11585_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11565_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11567_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11578_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26892_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26892_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26892_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26892_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26892_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26892_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26892_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26892_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26928_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26928_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26928_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26928_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26928_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26928_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26928_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26928_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26929_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26929_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26929_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26929_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26929_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26929_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26929_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26929_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26899_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26899_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26900_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26900_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26900_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26901_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26901_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26901_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26902_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26902_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26903_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26903_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26903_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26903_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26904_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26904_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _26905_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26893_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26893_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26893_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26894_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26894_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26894_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _26895_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _26895_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _26896_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _26896_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _26896_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _26896_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _26896_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _26896_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _26896_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _26896_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26897_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26898_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26898_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26944_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26906_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26906_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26906_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26906_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26906_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26906_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26906_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26906_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26907_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26907_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26907_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26907_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26907_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26907_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26907_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26907_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26908_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26908_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26908_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26908_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26908_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26908_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26908_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26908_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26909_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26909_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26909_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26909_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26909_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26909_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26909_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26909_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26910_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26910_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26910_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26910_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26910_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26910_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26910_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26910_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26911_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26911_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26911_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26911_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26911_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26911_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26911_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26911_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26912_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26912_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26912_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26912_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26912_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26912_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26912_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26912_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26913_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26913_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26913_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26913_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26913_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26913_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26913_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26913_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26917_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26917_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26917_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26917_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26917_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26914_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26914_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26914_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26914_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26914_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26914_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26914_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26914_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26914_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26914_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26914_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26914_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26914_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26914_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26914_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26914_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26915_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26915_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26915_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26915_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26915_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26915_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26915_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26915_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26915_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26915_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26915_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26915_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26915_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26915_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26915_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26915_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26935_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26935_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26935_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26935_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26935_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26935_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26935_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26935_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26935_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26935_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26935_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26935_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26935_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26935_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26935_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26935_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26935_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26935_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26935_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26935_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26935_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26935_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26935_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26935_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26935_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26935_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26935_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26935_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26935_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26935_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26935_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26935_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26918_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26918_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26918_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26918_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26918_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26918_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26918_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26918_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26921_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26921_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26921_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26921_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26921_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26921_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26921_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26921_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26921_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26921_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26921_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26921_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26921_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26921_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26921_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26921_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26922_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26922_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26922_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26922_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26922_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26922_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26922_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26922_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26922_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26922_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26922_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26922_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26922_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26922_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26922_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26922_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26926_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26926_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26926_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26926_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26926_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26926_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26926_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26926_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26927_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26927_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26927_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _26930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26931_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26931_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26931_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26931_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26931_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26931_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26931_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26931_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _26932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26934_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26934_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26934_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26934_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26936_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26936_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26936_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26936_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26936_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26936_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26936_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26936_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26936_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26936_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26936_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26936_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26936_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26936_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26936_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26936_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26936_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26936_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26936_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26936_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26936_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26936_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26936_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26936_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26936_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26936_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26936_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26936_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26936_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26936_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26936_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26936_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26940_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26940_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26940_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26940_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26941_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26942_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26943_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26943_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26943_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26943_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26943_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26943_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26943_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26943_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26945_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26945_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26945_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _05371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _05391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _05378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _04229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _05207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _27015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _04501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _05291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _09433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _06079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _06075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _09430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _09447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _27001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _05335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _05339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _05782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _05769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _09445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _05845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _05836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _05821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _09429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _26988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _26969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _22624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _12255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _05894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _05888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _05962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _05952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _05931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _05273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _04225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _04563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _05737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _05730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _27032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _05631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _05622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _22642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _27324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _22637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _22658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _22657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _12246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _16605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _27325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _22604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _11301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _22606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _27203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _11236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _11339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _22608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _27204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _27182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _27183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _27184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _11240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _22599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _11303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _11356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _22602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _22253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _22592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _11248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _22594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _11246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _22595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _11309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _22596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _10017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _09974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _10467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _09060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _09058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _09055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _09048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _09530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _10590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _10580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _10563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _10747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _10727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _09747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _09655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _10490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _10771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _11451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _11432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _11251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _10379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _11520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _27248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _10373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _22671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _23310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _22930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _08777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _22677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _22672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _22674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _08709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _10323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _08739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _00889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _10349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _02627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _02621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _10345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _06192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _09590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _10319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _11209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _10300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _05353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _05347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _10339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _27247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _27245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _26509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _10027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _27246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _25054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _25522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _08675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _08785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _06031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _08684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _03119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _03555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _03458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _02445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _02810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _02758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _05104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _08682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _09984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _04138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _08680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _05785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _05683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _09938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _27242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _07318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _10292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _09613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _06440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _04013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _04935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _09951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _08360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _27237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _08741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _27238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _27239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _27240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _27241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _08582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _11055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _11046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _11066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _11048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _07257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _10982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _07374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _07040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _11124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _11157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _11126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _11128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _09944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _27322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _11011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _10992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _09607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _10781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _27321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _10792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _10801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _09602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _10809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _09753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _10735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _27320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _09830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _10741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _10753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _09615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _10764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _09609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _09630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _10639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _10658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _09626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _10669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _10696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _10709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _10720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _10587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _10606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _09638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _10620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _27317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _27318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _27319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _09902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _09907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _10491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _10546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _09662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _10560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _09660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _10572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _09767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _09678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _09843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _10359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _10374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _27316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _10413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _09671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _10444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _10071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _09024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _10078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _10099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _09086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _10105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _10114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _09083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _10040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _27312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _09912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _10294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _27313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _09683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _10346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _09681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _26960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _11293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _07477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _07906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _11295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _26961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _07472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _11316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _11223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _07497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _11225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _11234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _07919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _11238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _11244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _26959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _26957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _26958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _07504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _11186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _07502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _11190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _07844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _11215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _07581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _10829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _10831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _26956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _10843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _10874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _07554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _07915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _06584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _04772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _04799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _06776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _22650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _10181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _26975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _10674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _07002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _06765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _08987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _06482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _01013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _05504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _26974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _06594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _26972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _26973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _08755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _06504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _09157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _05298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _06754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _27212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _05123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _05114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _02266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _26253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _04813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _04781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _27213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _05233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _05213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _05204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _05386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _05345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _05311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _27211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _05013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _27209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _05459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _05436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _02245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _05579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _02241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _26266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _27210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _27207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _27208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _06008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _25968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _05725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _05713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _05678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _05803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _27205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _06128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _06108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _06549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _06540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _06525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _27206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _05884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _06639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _27199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _06603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _06696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _27200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _27201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _25975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _27202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _26272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _06846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _27198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _06790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _06904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _06891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _06887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _02194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _07237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _02174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _06950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _27197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _07042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _07078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _07063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _07047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _25993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _00198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _07170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _07167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _07151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _07140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _07267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _27196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _27194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _07549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _26043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _07367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _07364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _27195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _07433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _07427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _02150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _07846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _27192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _02145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _26274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _07474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _27193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _07480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _10919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _10787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _11774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _11754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _11683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _27292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _11035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _10062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _08213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _08209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _27190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _08751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _08707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _27191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _07832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _07828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _09997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _27188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _09038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _08935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _09710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _09653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _27189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _00233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _10177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _10341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _10310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _26280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _09779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _02115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _10045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _27185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _00248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _10694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _27186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _02099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _10854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _02094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _10227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _07929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _06900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _01906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _26347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _04109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _27181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _03112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _02889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _11121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _27180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _11353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _26229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _08221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _09030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _08748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _26218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _10684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _27178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _10934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _26226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _01890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _27179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _26223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _11232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _10955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _10931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _02086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _11061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _11052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _27177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _26091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _00240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _27174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _26129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _27175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _11134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _02080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _27176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _11271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _02077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _27171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _27172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _12104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _02048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _11362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _11459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _27173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _11554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _12189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _12346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _12252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _11063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _12750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _12812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _27291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _11033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _12205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _12176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _27169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _12261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _00040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _02039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _26304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _27170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _02027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _08207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _02022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _26307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _01766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _02033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _05349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _26155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _08200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _08099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _08000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _08715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _08626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _08569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _11004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _27288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _27166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _02005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _27167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _09604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _10665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _09990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _02016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _27168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _06398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _11015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _07688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _07632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _07487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _10984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _13216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _27290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _05454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _10678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _01986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _26319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _27165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _02000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _01995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _22715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _27164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _00245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _12230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _12072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _01983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _09436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _03398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _07086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _08910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _08761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _09749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _09443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _27163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _02393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _01974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _04553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _14751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _14716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _27282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _27283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _27284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _11167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _14073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _14032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _11161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _27285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _15180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _27286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _11137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _15758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _15616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _27287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _27275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _07296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _27276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _00098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _08328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _22713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _22718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _25321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _08688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _10679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _27277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _10805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _27278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _27279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _07932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _10117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _24229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _24215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _12133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _27117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _24312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _27118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _27119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _24147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _07022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _25327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _27273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _27274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _06366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _10773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _08691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _22627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _24501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _24563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _12098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _26946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _24371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _26947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _26948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _24463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _27251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _23537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _23508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _12172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _27252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _27253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _23399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _23396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _23778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _27243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _23785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _23924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _27244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _23881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _11448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _23477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _24197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _24190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _12141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _23984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _23981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _12159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _24090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _24082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _22730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _22723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _27299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _22867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _22826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _11418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _27300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _22681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _11423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _22955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _23020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _23014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _23164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _27289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _23141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _12221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _23434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _23431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _11446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _23254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _23241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _12215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _27268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _23330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _22712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _27314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _12232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _22664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _27315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _22669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _22668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _22667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _22593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _11958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _02133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _27162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _26203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _05381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _09101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _01955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _10892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _27160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _10894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _03303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _27161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _10917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _02981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _03426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _03435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _10484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _03061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _10500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _03321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _10847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _10866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _03019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _03083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _03445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _10101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _10230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _03070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _10376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _03064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _10381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _09219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _27157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _03482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _09329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _03111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _09359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _27158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _27159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _03143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _08672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _03350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _08997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _03128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _09000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _03348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _09183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _07392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _07422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _03171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _03451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _07431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _03160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _27156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _03352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _03369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _27153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _07304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _03194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _27154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _07314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _07382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _27155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _03417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _02491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _03979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _03280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _03470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _03506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _07254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _07290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _01510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _03295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _01524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _03420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _27150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _03473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _01945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _02439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _07156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _03224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _07163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _27149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _07177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _07240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _03212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _03454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _03460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _06536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _03236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _06752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _03399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _06992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _07100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _03228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _27146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _03466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _05050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _27147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _03254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _27148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _03244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _05308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _01626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _05577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _27144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _04046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _04864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _03274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _27145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _03271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _27143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _26232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _02697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _00386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _00491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _05464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _00346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _01623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _05426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _05443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _26238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _05523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _05509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _27141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _00343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _27142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _27138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _03857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _27139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _27140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _03850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _05638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _05649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _05620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _27133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _04099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _27134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _27135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _27136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _03866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _27137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _04023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _03894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _04839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _04034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _04867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _27130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _03886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _27131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _03883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _04759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _04788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _03903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _04797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _04039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _27129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _04829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _04036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _04671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _04689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _03923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _27128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _03921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _04711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _04043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _04753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _04593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _27127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _04625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _04639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _03942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _04646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _04665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _03937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _03998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _04253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _03996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _04258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _04124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _04544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _04559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _04578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _04530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _03959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _27126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _04193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _04011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _04168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _04213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _04006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _04435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _03973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _04452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _03972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _04461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _04478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _27125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _04518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _04354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _03980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _04361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _27123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _04371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _04386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _27124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _04419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _02913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _05537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _27120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _04264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _27121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _27122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _04310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _04331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _03134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _03141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _05480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _02765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _02737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _05544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _02924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _26251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _05440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _03285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _03276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _03076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _03072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _03030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _27115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _27114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _26365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _26350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _05413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _26187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _26169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _05446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _26259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _03844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _03826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _27111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _27112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _05617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _26317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _26300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _27113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _03720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _03412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _03373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _03366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _03531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _03525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _03510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _05647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _27108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _10957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _27109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _27110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _03682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _03617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _05645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _03745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _03512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _11466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _11429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _27106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _27107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _00054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _03508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _01325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _27102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _27103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _00954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _27104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _26358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _10743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _09875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _01119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _27100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _27101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _03344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _03081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _03516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _23442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _22978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _08904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _27095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _27096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _27097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _27098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _05805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _05858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _27099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _09002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _27092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _09145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _27093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _27094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _08665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _08661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _08591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _09764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _09738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _10576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _10527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _10353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _27088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _03692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _27089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _10979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _10737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _10730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _11523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _11503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _11481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _27087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _09850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _00755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _04869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _23003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _22673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _27084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _09833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _27085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _27086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _06082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _05539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _03553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _27082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _22649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _27083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _04877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _01107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _09147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _11282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _11174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _27080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _03556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _27081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _03953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _04846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _09955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _09934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _09751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _09745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _27311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _09802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _10022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _27310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _09703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _10219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _10234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _10247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _10263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _10280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _09947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _09717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _10131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _27309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _10144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _09785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _09910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _10153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _10188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _09520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _10058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _09740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _10076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _10095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _10107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _27308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _11115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _11006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _10989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _11009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _07169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _11057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _11039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _27307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _10803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _27303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _10813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _09051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _27304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _27305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _11159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _27306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _10744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _10755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _08881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _10758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _10774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _27302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _09093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _10778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _09096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _10692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _10712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _08889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _10723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _08886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _10729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _09063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _27301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _09582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _10636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _10648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _08898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _10659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _08893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _10671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _10574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _09073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _10601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _27298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _10604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _09071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _10611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _10628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _08922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _10407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _27297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _10523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _08920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _10526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _09075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _10555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _09088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _10317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _10332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _08929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _10343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _10356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _10367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _08925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _09957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _27296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _09046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _09995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _10019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _09036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _10023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _10054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _09012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _27294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _09010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _10249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _10269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _27295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _08941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _09941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _09020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _10146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _09081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _10171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _27293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _10179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _10211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _09015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _03179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _03150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _02516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _03680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _03673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _03585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _10593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _27258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _08308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _08313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _23107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _00058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _10239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _08513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _08507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _08511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _05262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _27254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _05101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _05810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _05828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _27255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _27256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _27257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _22680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _22688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _22725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _10228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _22676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _22625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _10223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _08743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _08735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _07275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _07214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _07011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _08759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _08721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _08713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _27250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _27235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _10195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _01271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _10182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _27236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _22628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _10217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _22675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _09185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _10512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _08853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _08900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _08984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _08992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _08990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _27249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _10151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _27233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _08588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _08781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _10976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _07013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _27234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _10165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _07547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _15240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _10116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _08746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _09591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _10136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _10129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _08389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _23135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _11403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _08609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _08705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _23409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _08195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _12164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _09708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _00877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _08612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _22933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _27232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _22795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _11098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _10081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _22633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _27231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _11328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _13379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _23781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _24246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _24045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _08615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _24702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _11203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _27226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _11289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _27227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _11198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _27228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _27229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _27230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _22615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _22618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _27223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _27224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _22619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _11211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _27225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _11291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _11297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _27218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _27219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _27220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _27221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _22613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _22614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _27222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _11299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _27216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _22609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _11229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _11337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _11365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _22610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _27217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _07519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _07090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _07530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _09458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _05244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _04183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _05250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _05448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _27151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _16927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _27152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _16948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _17068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _11284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _17089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _11326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _11090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _09976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _11094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _10900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _07532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _10908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _04570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _12923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _12791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _03605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _09243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _04586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _11359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _11342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _03602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _07707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _07513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _08527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _08293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _03600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _27056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _05570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _03641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _23927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _23917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _24028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _04365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _03749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _27046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _04380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _27005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _07489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _07499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _07493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _06960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _07535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _07551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _27006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _07397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _27007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _06969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _07465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _06547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _27003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _08201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _08198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _06391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _07602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _07600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _07583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _27004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _08733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _08677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _09039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _06701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _12054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _12031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _09695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _27323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _09768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _11029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _09482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _10505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _10241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _11092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _10824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _06994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _04656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _10821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _08686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _08865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _27280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _27281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _12508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _07939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _15068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _08481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _22607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _04082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _27272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _07936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _01254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _01245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _01147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _07942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _27270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _05137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _05061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _27271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _05415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _06769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _10716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _07272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _07255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _10708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _08694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _27267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _01508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _01434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _27269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _10733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _08693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _08789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _25067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _00792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _02597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _05211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _05054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _05043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _10718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _01385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _01382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _01377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _11024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _27264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _11491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _10642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _08699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _27265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _10557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _10941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _08696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _07319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _07369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _07357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _10701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _08724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _08667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _27266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _10920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _10656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _09210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _09303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _09238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _10322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _10168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _10110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _07949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _06491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _05627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _10631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _15151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _10626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _27261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _08791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _27262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _08844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _27263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _19750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _09853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _10973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _07946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _11086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _19729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _19825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _11260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _11344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _21660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _21981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _11258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _27132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _11318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _18851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _19316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _27116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _11346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _19380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _19708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _11265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _05450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _27067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _05433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _05473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _05486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _09426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _05468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _17400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _17431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _11280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _17452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _11278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _27090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _11323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _27091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _11274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _05707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _05689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _05681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _07187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _05534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _27043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _05521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _05582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _04816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _01259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _27076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _23301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _27077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _27078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _04824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _27079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _27073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _22678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _22679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _08411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _04785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _08310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _08316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _08348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _00062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _27074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _03782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _08557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _27075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _08825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _08400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _08478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _06409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _11276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _04736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _22716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _27071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _04779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _03667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _27072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _03978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _00920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _03503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _27065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _03577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _22600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _12944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _07849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _19784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _27068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _27069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _03785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _08537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _27070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _03298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _04756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _24459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _15256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _07093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _04702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _02939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _04073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _22651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _27066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _27063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _06737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _25527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _03971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _00262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _00865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _03587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _27064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _22601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _22597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _25501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _25480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _27060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _27061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _03727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _27062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _27058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _04636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _00992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _00972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _00887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _26490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _02673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _27059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _04260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _03765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _13620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _13327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _04557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _04549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _12305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _05243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _06565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _06294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _04623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _27057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _03533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _03364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _04739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _25986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _26135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _26101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _03676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _25726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _25765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _25747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _03670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _25690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _25676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _04238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _27053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _25546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _27054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _25229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _24699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _03738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _25929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _25980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _25954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _25823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _25893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _04191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _26064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _16646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _04504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _14602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _14576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _04542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _15165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _15082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _15030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _19450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _04493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _22617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _22611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _03610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _15839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _15637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _16454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _27050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _04450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _22665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _22663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _22662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _04466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _22666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _22670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _03613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _22635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _22634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _27051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _22656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _22654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _04473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _27052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _23314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _03626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _27049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _04442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _23128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _04429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _03743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _22709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _24511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _24602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _04289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _03763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _24368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _04312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _24472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _24488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _03632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _23413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _27047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _27048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _03629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _03794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _23206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _23228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _04336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _24309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _04320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _24111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _27044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _27045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _24187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _24181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _04685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _04729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _05749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _06220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _24648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _04285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _27042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _04270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _05763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _27039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _27040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _04634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _06018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _04650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _05756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _27041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _04574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _27038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _04583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _04596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _05775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _06145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _04599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _05767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _05807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _04521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _06050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _04528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _27036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _05789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _27037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _04565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _04439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _04456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _05817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _04469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _27035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _04486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _06053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _06227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _05851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _04393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _27034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _04423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _05834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _06065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _05979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _27033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _04088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _06241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _04279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _04315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _05881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _04324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _05877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _06183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _04326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _05865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _04358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _05853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _04276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _05890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _06186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _04102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _05986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _04104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _06126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _04110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _04220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _04239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _05921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _06197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _04242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _04266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _04268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _06105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _04178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _04186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _05941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _06205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _04188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _04216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _27028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _07071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _09985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _07416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _07410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _09834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _27029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _27030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _04133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _06116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _27031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _04154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _05956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _06211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _04158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _04171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _04874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _04842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _27026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _27027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _07067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _04021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _04009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _04794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _07050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _27023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _27024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _27025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _07059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _05074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _05062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _06278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _05343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _27021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _27022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _07045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _06522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _05172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _07052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _05231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _05716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _05710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _05685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _07018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _05778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _05760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _05754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _27017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _05484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _05527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _27018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _27019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _05614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _07020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _05364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _27020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _06310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _06635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _05848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _05825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _07007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _05924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _27016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _05916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _06523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _06996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _05990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _05999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _07000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _06094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _06090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _06678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _06671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _06658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _06321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _27014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _06188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _06177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _06998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _27011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _06880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _06870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _06944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _06914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _06981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _27012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _06730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _06723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _06807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _06801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _06795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _27013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _06598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _06596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _07179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _06977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _06543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _27010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _06975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _06966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _07065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _07055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _07269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _27008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _07247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _07359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _07135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _07101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _27009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _08797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _08757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _08753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _27002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _06648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _08188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _07857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _07854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _08933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _09636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _09109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _09108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _09105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _27000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _08701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _06945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _09727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _06935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _09778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _09812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _09783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _06406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _08931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _09027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _10421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _10362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _10713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _10687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _26998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _10224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _10197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _10186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _10277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _10302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _06910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _09959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _09953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _09949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _09925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _26999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _11068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _10845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _10811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _26997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _10928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _06421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _10470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _06893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _11269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _11256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _06426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _06654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _26996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _06897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _11078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _12151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _12135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _06876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _26989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _26990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _26991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _26992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _26993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _26994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _06561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _11360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _11330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _11534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _11479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _06433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _26995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _27214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _02280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _04244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _04328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _27215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _04629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _04589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _04535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _06511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _04293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _04844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _04447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _03362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _04028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _03992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _06742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _26986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _06563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _26987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _06728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _06726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _05959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _06476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _03594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _06858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _03901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _04115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _06856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _06568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _07307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _10871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _08821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _07277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _26984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _12208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _12199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _26985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _08622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _06827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _00075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _06825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _06660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _06851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _09920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _26983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _00845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _26980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _06579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _26981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _11313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _06820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _26982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _06788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _26976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _26977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _26978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _06779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _26979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _09099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _25016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _26970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _26971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _01867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _26396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _26330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _11927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _26967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _26968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _12197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _07429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _12228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _07597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _12242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _10654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _11455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _07458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _26963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _11536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _26964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _26965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _26966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _07438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _11096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _07507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _26953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _07851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _10796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _26954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _10799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _26955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _01003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _01762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _01412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _07952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _23060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _22941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _27259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _27260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _11349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _07469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _07904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _07925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _11351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _26962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _07463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _11398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _07521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _11013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _26950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _26951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _07516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _11073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _07514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _26952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _07913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _10915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _26949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _07896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _10945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _11002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _07524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _07912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _08669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _08770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _27326_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _08768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _08896_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _27327_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27328_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27328_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27328_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27328_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _27329_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _27330_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27331_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27331_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27331_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27331_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27331_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27331_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27331_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27331_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10498_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10449_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10537_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10519_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10496_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _09774_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _09617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _09640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _09674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _09677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _09585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _09790_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _07414_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _10051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _10048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _09969_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _10161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _10141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _10008_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _10125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _10154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09971_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _10163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _10142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _10009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _10035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _10083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _10074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _10133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _06756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _14164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _14273_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _14243_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _14206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _14185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _06762_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _13569_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _05635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _13488_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _05643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _13761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _06001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _13095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _13348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _05987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _06123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _06100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _06068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _12637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _12623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _12608_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _05873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _12128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _11999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _12107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _12084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _12030_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22647_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _12397_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _05868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _11591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _11560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _11532_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _11487_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _11846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _11795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _05997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _22655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _22653_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _22652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _06571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _22661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _22660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _22659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _22626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _06629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _22641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _22640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _22639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _22638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _06582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _22623_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _22622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _22621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _22620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _06632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _00829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _22612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _22616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _06669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _00819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _00892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _00923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _22605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _22603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _10922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10364_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _10149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _09828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _09927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _09880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _09848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _09930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _09929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _09878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _03215_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _00672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _22629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04871_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _23188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _26000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _22598_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _03205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _23172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _23596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _23641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _25995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _22717_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _25315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _24680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _03529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _23033_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12248_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _01225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _08463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _08524_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _22636_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _10174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _10087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _11183_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _11165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _11163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _11145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _03559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _15990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _09091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _09065_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04947_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _22726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _23593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _23638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _23658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _10817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _07057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _07049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _04173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _07327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _07334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _07331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _04144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _07244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _07072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _07284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _07282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _04174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _07203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _07189_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _07198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _07069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _04180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _24066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _11108_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _11104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _11100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _03574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _03595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _11083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _11081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _03589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _11041_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _11037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _11027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _03615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _22232_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _11152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _11141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _11139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _06939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _22884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _22893_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _22890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _22887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01505_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _26328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _26325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _26344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _26342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _02305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01504_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22792_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _26289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _26282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _26288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02381_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _26309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22689_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _26306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22682_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _22692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02378_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22686_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01502_);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
