
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_rom_pc, property_invalid_dec_rom_pc, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IE_gm_next;
  wire [7:0] IP_gm;
  wire [7:0] IP_gm_next;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PCON_gm_next;
  wire [15:0] PC_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SBUF_gm_next;
  wire [7:0] SCON_gm;
  wire [7:0] SCON_gm_next;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TCON_gm_next;
  wire [7:0] TH0_gm;
  wire [7:0] TH0_gm_next;
  wire [7:0] TH1_gm;
  wire [7:0] TH1_gm_next;
  wire [7:0] TL0_gm;
  wire [7:0] TL0_gm_next;
  wire [7:0] TL1_gm;
  wire [7:0] TL1_gm_next;
  wire [7:0] TMOD_gm;
  wire [7:0] TMOD_gm_next;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IE_next ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IP_next ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [7:0] \oc8051_golden_model_1.PCON_next ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SBUF_next ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SCON_next ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TCON_next ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH0_next ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TH1_next ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL0_next ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TL1_next ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire [7:0] \oc8051_golden_model_1.TMOD_next ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire \oc8051_golden_model_1.n1046 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire \oc8051_golden_model_1.n1063 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1148 ;
  wire [3:0] \oc8051_golden_model_1.n1150 ;
  wire [3:0] \oc8051_golden_model_1.n1151 ;
  wire [3:0] \oc8051_golden_model_1.n1152 ;
  wire [3:0] \oc8051_golden_model_1.n1153 ;
  wire [3:0] \oc8051_golden_model_1.n1154 ;
  wire [3:0] \oc8051_golden_model_1.n1155 ;
  wire [3:0] \oc8051_golden_model_1.n1156 ;
  wire \oc8051_golden_model_1.n1202 ;
  wire \oc8051_golden_model_1.n1244 ;
  wire [8:0] \oc8051_golden_model_1.n1245 ;
  wire [8:0] \oc8051_golden_model_1.n1246 ;
  wire [7:0] \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire [2:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire [1:0] \oc8051_golden_model_1.n1251 ;
  wire [7:0] \oc8051_golden_model_1.n1252 ;
  wire [6:0] \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1255 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire \oc8051_golden_model_1.n1258 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire \oc8051_golden_model_1.n1260 ;
  wire \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1268 ;
  wire [7:0] \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1285 ;
  wire [7:0] \oc8051_golden_model_1.n1286 ;
  wire [15:0] \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1319 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire \oc8051_golden_model_1.n1321 ;
  wire \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire \oc8051_golden_model_1.n1324 ;
  wire \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1334 ;
  wire [7:0] \oc8051_golden_model_1.n1335 ;
  wire [8:0] \oc8051_golden_model_1.n1337 ;
  wire [8:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire [3:0] \oc8051_golden_model_1.n1343 ;
  wire [4:0] \oc8051_golden_model_1.n1344 ;
  wire [4:0] \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [8:0] \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire [7:0] \oc8051_golden_model_1.n1359 ;
  wire [6:0] \oc8051_golden_model_1.n1360 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [7:0] \oc8051_golden_model_1.n1376 ;
  wire [8:0] \oc8051_golden_model_1.n1398 ;
  wire \oc8051_golden_model_1.n1399 ;
  wire [4:0] \oc8051_golden_model_1.n1404 ;
  wire \oc8051_golden_model_1.n1405 ;
  wire \oc8051_golden_model_1.n1413 ;
  wire [7:0] \oc8051_golden_model_1.n1414 ;
  wire [6:0] \oc8051_golden_model_1.n1415 ;
  wire \oc8051_golden_model_1.n1430 ;
  wire [7:0] \oc8051_golden_model_1.n1431 ;
  wire [8:0] \oc8051_golden_model_1.n1433 ;
  wire [8:0] \oc8051_golden_model_1.n1435 ;
  wire \oc8051_golden_model_1.n1436 ;
  wire [3:0] \oc8051_golden_model_1.n1437 ;
  wire [4:0] \oc8051_golden_model_1.n1438 ;
  wire [4:0] \oc8051_golden_model_1.n1440 ;
  wire \oc8051_golden_model_1.n1441 ;
  wire [8:0] \oc8051_golden_model_1.n1442 ;
  wire \oc8051_golden_model_1.n1449 ;
  wire [7:0] \oc8051_golden_model_1.n1450 ;
  wire [6:0] \oc8051_golden_model_1.n1451 ;
  wire \oc8051_golden_model_1.n1466 ;
  wire [7:0] \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1470 ;
  wire \oc8051_golden_model_1.n1471 ;
  wire \oc8051_golden_model_1.n1478 ;
  wire [7:0] \oc8051_golden_model_1.n1479 ;
  wire [6:0] \oc8051_golden_model_1.n1480 ;
  wire [7:0] \oc8051_golden_model_1.n1481 ;
  wire [8:0] \oc8051_golden_model_1.n1483 ;
  wire [8:0] \oc8051_golden_model_1.n1485 ;
  wire \oc8051_golden_model_1.n1486 ;
  wire [4:0] \oc8051_golden_model_1.n1487 ;
  wire [4:0] \oc8051_golden_model_1.n1489 ;
  wire \oc8051_golden_model_1.n1490 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire \oc8051_golden_model_1.n1498 ;
  wire [7:0] \oc8051_golden_model_1.n1499 ;
  wire [6:0] \oc8051_golden_model_1.n1500 ;
  wire \oc8051_golden_model_1.n1515 ;
  wire [7:0] \oc8051_golden_model_1.n1516 ;
  wire [4:0] \oc8051_golden_model_1.n1518 ;
  wire \oc8051_golden_model_1.n1519 ;
  wire [7:0] \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire [8:0] \oc8051_golden_model_1.n1524 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire \oc8051_golden_model_1.n1532 ;
  wire [7:0] \oc8051_golden_model_1.n1533 ;
  wire [6:0] \oc8051_golden_model_1.n1534 ;
  wire [7:0] \oc8051_golden_model_1.n1535 ;
  wire [7:0] \oc8051_golden_model_1.n1536 ;
  wire [6:0] \oc8051_golden_model_1.n1537 ;
  wire [7:0] \oc8051_golden_model_1.n1538 ;
  wire [8:0] \oc8051_golden_model_1.n1541 ;
  wire [8:0] \oc8051_golden_model_1.n1542 ;
  wire [7:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [6:0] \oc8051_golden_model_1.n1545 ;
  wire \oc8051_golden_model_1.n1546 ;
  wire \oc8051_golden_model_1.n1547 ;
  wire \oc8051_golden_model_1.n1548 ;
  wire \oc8051_golden_model_1.n1549 ;
  wire \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1552 ;
  wire \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [8:0] \oc8051_golden_model_1.n1565 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire \oc8051_golden_model_1.n1568 ;
  wire [4:0] \oc8051_golden_model_1.n1569 ;
  wire [4:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire [7:0] \oc8051_golden_model_1.n1580 ;
  wire [6:0] \oc8051_golden_model_1.n1581 ;
  wire \oc8051_golden_model_1.n1596 ;
  wire [7:0] \oc8051_golden_model_1.n1597 ;
  wire [8:0] \oc8051_golden_model_1.n1601 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [4:0] \oc8051_golden_model_1.n1604 ;
  wire \oc8051_golden_model_1.n1605 ;
  wire \oc8051_golden_model_1.n1612 ;
  wire [7:0] \oc8051_golden_model_1.n1613 ;
  wire [6:0] \oc8051_golden_model_1.n1614 ;
  wire \oc8051_golden_model_1.n1629 ;
  wire [7:0] \oc8051_golden_model_1.n1630 ;
  wire [8:0] \oc8051_golden_model_1.n1634 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [4:0] \oc8051_golden_model_1.n1637 ;
  wire \oc8051_golden_model_1.n1638 ;
  wire \oc8051_golden_model_1.n1645 ;
  wire [7:0] \oc8051_golden_model_1.n1646 ;
  wire [6:0] \oc8051_golden_model_1.n1647 ;
  wire \oc8051_golden_model_1.n1662 ;
  wire [7:0] \oc8051_golden_model_1.n1663 ;
  wire [8:0] \oc8051_golden_model_1.n1667 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [4:0] \oc8051_golden_model_1.n1670 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire \oc8051_golden_model_1.n1678 ;
  wire [7:0] \oc8051_golden_model_1.n1679 ;
  wire [6:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1695 ;
  wire [7:0] \oc8051_golden_model_1.n1696 ;
  wire [7:0] \oc8051_golden_model_1.n1710 ;
  wire [6:0] \oc8051_golden_model_1.n1711 ;
  wire [7:0] \oc8051_golden_model_1.n1712 ;
  wire \oc8051_golden_model_1.n1756 ;
  wire [7:0] \oc8051_golden_model_1.n1757 ;
  wire \oc8051_golden_model_1.n1773 ;
  wire [7:0] \oc8051_golden_model_1.n1774 ;
  wire \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire \oc8051_golden_model_1.n1807 ;
  wire [7:0] \oc8051_golden_model_1.n1808 ;
  wire [7:0] \oc8051_golden_model_1.n1820 ;
  wire [6:0] \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1866 ;
  wire [7:0] \oc8051_golden_model_1.n1867 ;
  wire \oc8051_golden_model_1.n1883 ;
  wire [7:0] \oc8051_golden_model_1.n1884 ;
  wire \oc8051_golden_model_1.n1900 ;
  wire [7:0] \oc8051_golden_model_1.n1901 ;
  wire \oc8051_golden_model_1.n1917 ;
  wire [7:0] \oc8051_golden_model_1.n1918 ;
  wire \oc8051_golden_model_1.n1993 ;
  wire [7:0] \oc8051_golden_model_1.n1994 ;
  wire \oc8051_golden_model_1.n2010 ;
  wire [7:0] \oc8051_golden_model_1.n2011 ;
  wire \oc8051_golden_model_1.n2027 ;
  wire [7:0] \oc8051_golden_model_1.n2028 ;
  wire \oc8051_golden_model_1.n2044 ;
  wire [7:0] \oc8051_golden_model_1.n2045 ;
  wire \oc8051_golden_model_1.n2049 ;
  wire [6:0] \oc8051_golden_model_1.n2050 ;
  wire [7:0] \oc8051_golden_model_1.n2051 ;
  wire [6:0] \oc8051_golden_model_1.n2052 ;
  wire [7:0] \oc8051_golden_model_1.n2053 ;
  wire \oc8051_golden_model_1.n2068 ;
  wire [7:0] \oc8051_golden_model_1.n2069 ;
  wire \oc8051_golden_model_1.n2097 ;
  wire [7:0] \oc8051_golden_model_1.n2098 ;
  wire [6:0] \oc8051_golden_model_1.n2099 ;
  wire [7:0] \oc8051_golden_model_1.n2100 ;
  wire [3:0] \oc8051_golden_model_1.n2107 ;
  wire \oc8051_golden_model_1.n2108 ;
  wire [7:0] \oc8051_golden_model_1.n2109 ;
  wire [6:0] \oc8051_golden_model_1.n2110 ;
  wire \oc8051_golden_model_1.n2125 ;
  wire [7:0] \oc8051_golden_model_1.n2126 ;
  wire [7:0] \oc8051_golden_model_1.n2301 ;
  wire \oc8051_golden_model_1.n2304 ;
  wire \oc8051_golden_model_1.n2306 ;
  wire \oc8051_golden_model_1.n2312 ;
  wire [7:0] \oc8051_golden_model_1.n2313 ;
  wire [6:0] \oc8051_golden_model_1.n2314 ;
  wire \oc8051_golden_model_1.n2329 ;
  wire [7:0] \oc8051_golden_model_1.n2330 ;
  wire \oc8051_golden_model_1.n2334 ;
  wire \oc8051_golden_model_1.n2336 ;
  wire \oc8051_golden_model_1.n2342 ;
  wire [7:0] \oc8051_golden_model_1.n2343 ;
  wire [6:0] \oc8051_golden_model_1.n2344 ;
  wire \oc8051_golden_model_1.n2359 ;
  wire [7:0] \oc8051_golden_model_1.n2360 ;
  wire \oc8051_golden_model_1.n2364 ;
  wire \oc8051_golden_model_1.n2366 ;
  wire \oc8051_golden_model_1.n2372 ;
  wire [7:0] \oc8051_golden_model_1.n2373 ;
  wire [6:0] \oc8051_golden_model_1.n2374 ;
  wire \oc8051_golden_model_1.n2389 ;
  wire [7:0] \oc8051_golden_model_1.n2390 ;
  wire \oc8051_golden_model_1.n2394 ;
  wire \oc8051_golden_model_1.n2396 ;
  wire \oc8051_golden_model_1.n2402 ;
  wire [7:0] \oc8051_golden_model_1.n2403 ;
  wire [6:0] \oc8051_golden_model_1.n2404 ;
  wire \oc8051_golden_model_1.n2419 ;
  wire [7:0] \oc8051_golden_model_1.n2420 ;
  wire \oc8051_golden_model_1.n2422 ;
  wire [7:0] \oc8051_golden_model_1.n2423 ;
  wire [6:0] \oc8051_golden_model_1.n2424 ;
  wire [7:0] \oc8051_golden_model_1.n2425 ;
  wire [7:0] \oc8051_golden_model_1.n2426 ;
  wire [6:0] \oc8051_golden_model_1.n2427 ;
  wire [7:0] \oc8051_golden_model_1.n2428 ;
  wire [15:0] \oc8051_golden_model_1.n2432 ;
  wire \oc8051_golden_model_1.n2438 ;
  wire [7:0] \oc8051_golden_model_1.n2439 ;
  wire [6:0] \oc8051_golden_model_1.n2440 ;
  wire \oc8051_golden_model_1.n2455 ;
  wire [7:0] \oc8051_golden_model_1.n2456 ;
  wire \oc8051_golden_model_1.n2459 ;
  wire [7:0] \oc8051_golden_model_1.n2460 ;
  wire [6:0] \oc8051_golden_model_1.n2461 ;
  wire [7:0] \oc8051_golden_model_1.n2462 ;
  wire \oc8051_golden_model_1.n2490 ;
  wire [7:0] \oc8051_golden_model_1.n2491 ;
  wire [6:0] \oc8051_golden_model_1.n2492 ;
  wire [7:0] \oc8051_golden_model_1.n2493 ;
  wire \oc8051_golden_model_1.n2498 ;
  wire [7:0] \oc8051_golden_model_1.n2499 ;
  wire [6:0] \oc8051_golden_model_1.n2500 ;
  wire [7:0] \oc8051_golden_model_1.n2501 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire [7:0] \oc8051_golden_model_1.n2507 ;
  wire [6:0] \oc8051_golden_model_1.n2508 ;
  wire [7:0] \oc8051_golden_model_1.n2509 ;
  wire \oc8051_golden_model_1.n2514 ;
  wire [7:0] \oc8051_golden_model_1.n2515 ;
  wire [6:0] \oc8051_golden_model_1.n2516 ;
  wire [7:0] \oc8051_golden_model_1.n2517 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire [7:0] \oc8051_golden_model_1.n2523 ;
  wire [6:0] \oc8051_golden_model_1.n2524 ;
  wire [7:0] \oc8051_golden_model_1.n2525 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire [7:0] \oc8051_golden_model_1.n2548 ;
  wire [3:0] \oc8051_golden_model_1.n2549 ;
  wire [7:0] \oc8051_golden_model_1.n2550 ;
  wire \oc8051_golden_model_1.n2551 ;
  wire \oc8051_golden_model_1.n2552 ;
  wire \oc8051_golden_model_1.n2553 ;
  wire \oc8051_golden_model_1.n2554 ;
  wire \oc8051_golden_model_1.n2555 ;
  wire \oc8051_golden_model_1.n2556 ;
  wire \oc8051_golden_model_1.n2557 ;
  wire \oc8051_golden_model_1.n2558 ;
  wire \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [7:0] \oc8051_golden_model_1.n2575 ;
  wire [6:0] \oc8051_golden_model_1.n2576 ;
  wire \oc8051_golden_model_1.n2591 ;
  wire [7:0] \oc8051_golden_model_1.n2592 ;
  wire \oc8051_golden_model_1.n2593 ;
  wire \oc8051_golden_model_1.n2594 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2597 ;
  wire \oc8051_golden_model_1.n2598 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire \oc8051_golden_model_1.n2600 ;
  wire \oc8051_golden_model_1.n2607 ;
  wire [7:0] \oc8051_golden_model_1.n2608 ;
  wire \oc8051_golden_model_1.n2609 ;
  wire \oc8051_golden_model_1.n2610 ;
  wire \oc8051_golden_model_1.n2611 ;
  wire \oc8051_golden_model_1.n2612 ;
  wire \oc8051_golden_model_1.n2613 ;
  wire \oc8051_golden_model_1.n2614 ;
  wire \oc8051_golden_model_1.n2615 ;
  wire \oc8051_golden_model_1.n2616 ;
  wire \oc8051_golden_model_1.n2623 ;
  wire [7:0] \oc8051_golden_model_1.n2624 ;
  wire [7:0] \oc8051_golden_model_1.n2652 ;
  wire [6:0] \oc8051_golden_model_1.n2653 ;
  wire [7:0] \oc8051_golden_model_1.n2654 ;
  wire \oc8051_golden_model_1.n2673 ;
  wire [7:0] \oc8051_golden_model_1.n2674 ;
  wire [6:0] \oc8051_golden_model_1.n2675 ;
  wire \oc8051_golden_model_1.n2690 ;
  wire [7:0] \oc8051_golden_model_1.n2691 ;
  wire [7:0] \oc8051_golden_model_1.n2695 ;
  wire [3:0] \oc8051_golden_model_1.n2696 ;
  wire [7:0] \oc8051_golden_model_1.n2697 ;
  wire \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2712 ;
  wire [7:0] \oc8051_golden_model_1.n2713 ;
  wire \oc8051_golden_model_1.n2731 ;
  wire [7:0] \oc8051_golden_model_1.n2732 ;
  wire [7:0] \oc8051_golden_model_1.n2733 ;
  wire \oc8051_golden_model_1.n2749 ;
  wire [7:0] \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc_impl;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dec_rom_pc;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_rom_pc;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_36029_, rst);
  not (_14681_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_14692_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_14703_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _14692_);
  and (_14714_, _14703_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_14725_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _14692_);
  and (_14736_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _14692_);
  nor (_14747_, _14736_, _14725_);
  and (_14758_, _14747_, _14714_);
  nor (_14769_, _14758_, _14681_);
  and (_14780_, _14681_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_14790_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_14801_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _14790_);
  nor (_14812_, _14801_, _14780_);
  not (_14823_, _14812_);
  and (_14834_, _14823_, _14758_);
  or (_14845_, _14834_, _14769_);
  and (_24753_, _14845_, _36029_);
  nor (_14866_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_14877_, _14866_);
  and (_14888_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_14899_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_14910_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_14921_, _14910_);
  not (_14932_, _14801_);
  nor (_14953_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_14954_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_14965_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14954_);
  nor (_14976_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_14987_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_14998_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _14987_);
  nor (_15009_, _14998_, _14976_);
  nor (_15020_, _15009_, _14965_);
  not (_15031_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15042_, _14965_, _15031_);
  nor (_15053_, _15042_, _15020_);
  and (_15064_, _15053_, _14953_);
  not (_15075_, _15064_);
  and (_15086_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15097_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_15107_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15118_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _15107_);
  and (_15129_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_15140_, _15129_, _15097_);
  and (_15151_, _15140_, _15075_);
  nor (_15162_, _15151_, _14932_);
  not (_15173_, _14780_);
  nor (_15184_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_15195_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _14987_);
  nor (_15206_, _15195_, _15184_);
  nor (_15217_, _15206_, _14965_);
  not (_15228_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_15239_, _14965_, _15228_);
  nor (_15250_, _15239_, _15217_);
  and (_15261_, _15250_, _14953_);
  not (_15272_, _15261_);
  and (_15283_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_15294_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15305_, _15294_, _15283_);
  and (_15316_, _15305_, _15272_);
  nor (_15327_, _15316_, _15173_);
  nor (_15338_, _15327_, _15162_);
  nor (_15349_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_15360_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _14987_);
  nor (_15371_, _15360_, _15349_);
  nor (_15382_, _15371_, _14965_);
  not (_15393_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_15404_, _14965_, _15393_);
  nor (_15415_, _15404_, _15382_);
  and (_15426_, _15415_, _14953_);
  not (_15436_, _15426_);
  and (_15447_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_15458_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_15469_, _15458_, _15447_);
  and (_15480_, _15469_, _15436_);
  nor (_15491_, _15480_, _14823_);
  nor (_15502_, _15491_, _14866_);
  and (_15513_, _15502_, _15338_);
  nor (_15523_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_15534_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _14987_);
  nor (_15545_, _15534_, _15523_);
  nor (_15556_, _15545_, _14965_);
  not (_15567_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_15578_, _14965_, _15567_);
  nor (_15589_, _15578_, _15556_);
  and (_15600_, _15589_, _14953_);
  not (_15611_, _15600_);
  and (_15621_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_15632_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_15643_, _15632_, _15621_);
  and (_15654_, _15643_, _15611_);
  and (_15665_, _15654_, _14866_);
  nor (_15676_, _15665_, _15513_);
  not (_15687_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_15698_, _15687_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15708_, _15698_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15719_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_15730_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15741_, _15730_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15752_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_15763_, _15752_, _15719_);
  nor (_15774_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15785_, _15774_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_15796_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_15806_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15817_, _15698_, _15806_);
  and (_15828_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_15839_, _15828_, _15796_);
  and (_15850_, _15839_, _15763_);
  and (_15861_, _15774_, _15687_);
  and (_15872_, _15861_, _15589_);
  and (_15883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_15894_, _15883_, _15806_);
  and (_15904_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_15915_, _15883_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_15926_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_15937_, _15926_, _15904_);
  not (_15948_, _15937_);
  nor (_15959_, _15948_, _15872_);
  and (_15970_, _15959_, _15850_);
  not (_15981_, _15970_);
  and (_15991_, _15981_, _15676_);
  not (_16002_, _15991_);
  nor (_16013_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16024_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _14987_);
  nor (_16035_, _16024_, _16013_);
  nor (_16046_, _16035_, _14965_);
  not (_16057_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_16068_, _14965_, _16057_);
  nor (_16079_, _16068_, _16046_);
  and (_16089_, _16079_, _14953_);
  not (_16100_, _16089_);
  and (_16111_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_16122_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_16133_, _16122_, _16111_);
  and (_16144_, _16133_, _16100_);
  nor (_16155_, _16144_, _14932_);
  nor (_16166_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_16176_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _14987_);
  nor (_16187_, _16176_, _16166_);
  nor (_16198_, _16187_, _14965_);
  not (_16209_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_16220_, _14965_, _16209_);
  nor (_16231_, _16220_, _16198_);
  and (_16242_, _16231_, _14953_);
  not (_16253_, _16242_);
  and (_16264_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_16274_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16285_, _16274_, _16264_);
  and (_16296_, _16285_, _16253_);
  nor (_16307_, _16296_, _15173_);
  nor (_16318_, _16307_, _16155_);
  nor (_16329_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_16340_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _14987_);
  nor (_16351_, _16340_, _16329_);
  nor (_16361_, _16351_, _14965_);
  not (_16372_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_16383_, _14965_, _16372_);
  nor (_16394_, _16383_, _16361_);
  and (_16405_, _16394_, _14953_);
  not (_16416_, _16405_);
  and (_16427_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_16438_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_16449_, _16438_, _16427_);
  and (_16459_, _16449_, _16416_);
  nor (_16470_, _16459_, _14823_);
  nor (_16481_, _16470_, _14866_);
  and (_16492_, _16481_, _16318_);
  nor (_16503_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_16514_, _14987_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_16525_, _16514_, _16503_);
  nor (_16536_, _16525_, _14965_);
  not (_16547_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_16557_, _14965_, _16547_);
  nor (_16568_, _16557_, _16536_);
  and (_16579_, _16568_, _14953_);
  not (_16590_, _16579_);
  and (_16601_, _15086_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_16612_, _15118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_16623_, _16612_, _16601_);
  and (_16634_, _16623_, _16590_);
  and (_16644_, _16634_, _14866_);
  nor (_16655_, _16644_, _16492_);
  and (_16666_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_16688_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_16689_, _16688_, _16666_);
  and (_16700_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_16711_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_16722_, _16711_, _16700_);
  and (_16733_, _16722_, _16689_);
  and (_16740_, _16568_, _15861_);
  and (_16741_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_16751_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_16762_, _16751_, _16741_);
  not (_16773_, _16762_);
  nor (_16784_, _16773_, _16740_);
  and (_16795_, _16784_, _16733_);
  not (_16806_, _16795_);
  and (_16817_, _16806_, _16655_);
  and (_16828_, _16817_, _16002_);
  not (_16839_, _16828_);
  and (_16850_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_16860_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_16871_, _16860_, _16850_);
  and (_16882_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_16893_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_16904_, _16893_, _16882_);
  and (_16915_, _16904_, _16871_);
  and (_16926_, _16231_, _15861_);
  and (_16937_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_16948_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16959_, _16948_, _16937_);
  not (_16970_, _16959_);
  nor (_16981_, _16970_, _16926_);
  and (_16991_, _16981_, _16915_);
  not (_17002_, _16991_);
  and (_17013_, _17002_, _16655_);
  and (_17024_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17035_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17046_, _17035_, _17024_);
  and (_17057_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_17068_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_17079_, _17068_, _17057_);
  and (_17090_, _17079_, _17046_);
  and (_17101_, _15861_, _15250_);
  and (_17112_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_17122_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_17133_, _17122_, _17112_);
  not (_17144_, _17133_);
  nor (_17155_, _17144_, _17101_);
  and (_17166_, _17155_, _17090_);
  not (_17177_, _17166_);
  and (_17188_, _17177_, _15676_);
  and (_17199_, _17013_, _17188_);
  nor (_17210_, _15991_, _17199_);
  and (_17221_, _15981_, _17199_);
  nor (_17232_, _17221_, _17210_);
  and (_17242_, _17232_, _17013_);
  and (_17253_, _16817_, _15991_);
  and (_17264_, _15981_, _16655_);
  and (_17275_, _16806_, _15676_);
  nor (_17286_, _17275_, _17264_);
  nor (_17297_, _17286_, _17253_);
  and (_17308_, _17297_, _17242_);
  and (_17319_, _17297_, _17221_);
  nor (_17330_, _17319_, _17308_);
  nor (_17341_, _17330_, _16839_);
  and (_17352_, _16655_, _17177_);
  and (_17363_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_17373_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_17394_, _17373_, _17363_);
  and (_17395_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_17416_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_17417_, _17416_, _17395_);
  and (_17428_, _17417_, _17394_);
  and (_17439_, _16079_, _15861_);
  and (_17450_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_17461_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_17472_, _17461_, _17450_);
  not (_17483_, _17472_);
  nor (_17493_, _17483_, _17439_);
  and (_17504_, _17493_, _17428_);
  not (_17515_, _17504_);
  and (_17526_, _17515_, _15676_);
  and (_17537_, _17526_, _17352_);
  and (_17548_, _17002_, _15676_);
  nor (_17559_, _17548_, _17352_);
  nor (_17570_, _17559_, _17199_);
  and (_17581_, _17570_, _17537_);
  nor (_17592_, _15991_, _17013_);
  nor (_17603_, _17592_, _17242_);
  and (_17614_, _17603_, _17581_);
  nor (_17624_, _17297_, _17242_);
  nor (_17635_, _17624_, _17308_);
  nor (_17646_, _17635_, _17221_);
  nor (_17657_, _17646_, _17319_);
  and (_17668_, _17657_, _17614_);
  nor (_17679_, _17657_, _17614_);
  nor (_17690_, _17679_, _17668_);
  not (_17701_, _17690_);
  and (_17712_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_17722_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_17733_, _17722_, _17712_);
  and (_17744_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_17755_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_17766_, _17755_, _17744_);
  and (_17777_, _17766_, _17733_);
  and (_17788_, _16394_, _15861_);
  and (_17799_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_17810_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_17821_, _17810_, _17799_);
  not (_17832_, _17821_);
  nor (_17842_, _17832_, _17788_);
  and (_17853_, _17842_, _17777_);
  not (_17864_, _17853_);
  and (_17875_, _17864_, _16655_);
  and (_17886_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_17897_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_17908_, _17897_, _17886_);
  and (_17919_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_17930_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_17941_, _17930_, _17919_);
  and (_17951_, _17941_, _17908_);
  and (_17962_, _15861_, _15053_);
  and (_17973_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_17984_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_17995_, _17984_, _17973_);
  not (_18006_, _17995_);
  nor (_18017_, _18006_, _17962_);
  and (_18028_, _18017_, _17951_);
  not (_18039_, _18028_);
  and (_18050_, _18039_, _15676_);
  and (_18060_, _18050_, _17875_);
  and (_18071_, _17864_, _15676_);
  not (_18082_, _18071_);
  and (_18093_, _18039_, _16655_);
  and (_18104_, _18093_, _18082_);
  and (_18115_, _18104_, _17526_);
  nor (_18126_, _18115_, _18060_);
  and (_18137_, _17515_, _16655_);
  nor (_18148_, _18137_, _17188_);
  nor (_18159_, _18148_, _17537_);
  not (_18170_, _18159_);
  nor (_18180_, _18170_, _18126_);
  nor (_18191_, _17570_, _17537_);
  nor (_18202_, _18191_, _17581_);
  and (_18213_, _18202_, _18180_);
  nor (_18224_, _17603_, _17581_);
  nor (_18235_, _18224_, _17614_);
  and (_18246_, _18235_, _18213_);
  and (_18257_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_18268_, _15741_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_18279_, _18268_, _18257_);
  and (_18289_, _15785_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_18300_, _15817_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_18311_, _18300_, _18289_);
  and (_18322_, _18311_, _18279_);
  and (_18333_, _15861_, _15415_);
  and (_18344_, _15894_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18355_, _15915_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_18366_, _18355_, _18344_);
  not (_18377_, _18366_);
  nor (_18388_, _18377_, _18333_);
  and (_18398_, _18388_, _18322_);
  not (_18409_, _18398_);
  and (_18420_, _18409_, _16655_);
  and (_18431_, _18420_, _18071_);
  nor (_18442_, _18050_, _17875_);
  nor (_18453_, _18442_, _18060_);
  and (_18464_, _18453_, _18431_);
  nor (_18475_, _18104_, _17526_);
  nor (_18486_, _18475_, _18115_);
  and (_18497_, _18486_, _18464_);
  and (_18507_, _18170_, _18126_);
  nor (_18518_, _18507_, _18180_);
  and (_18529_, _18518_, _18497_);
  nor (_18540_, _18202_, _18180_);
  nor (_18551_, _18540_, _18213_);
  and (_18562_, _18551_, _18529_);
  nor (_18573_, _18235_, _18213_);
  nor (_18584_, _18573_, _18246_);
  and (_18595_, _18584_, _18562_);
  nor (_18606_, _18595_, _18246_);
  nor (_18616_, _18606_, _17701_);
  nor (_18627_, _18616_, _17668_);
  and (_18638_, _17330_, _16839_);
  nor (_18649_, _18638_, _17341_);
  not (_18660_, _18649_);
  nor (_18671_, _18660_, _18627_);
  or (_18682_, _18671_, _17253_);
  nor (_18693_, _18682_, _17341_);
  nor (_18704_, _18693_, _14921_);
  and (_18715_, _18693_, _14921_);
  nor (_18725_, _18715_, _18704_);
  not (_18736_, _18725_);
  and (_18747_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_18758_, _18660_, _18627_);
  nor (_18769_, _18758_, _18671_);
  and (_18780_, _18769_, _18747_);
  and (_18791_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_18802_, _18606_, _17701_);
  nor (_18813_, _18802_, _18616_);
  and (_18824_, _18813_, _18791_);
  nor (_18835_, _18813_, _18791_);
  nor (_18845_, _18835_, _18824_);
  not (_18856_, _18845_);
  and (_18867_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_18878_, _18584_, _18562_);
  nor (_18889_, _18878_, _18595_);
  and (_18900_, _18889_, _18867_);
  nor (_18911_, _18889_, _18867_);
  nor (_18922_, _18911_, _18900_);
  not (_18933_, _18922_);
  and (_18944_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_18954_, _18551_, _18529_);
  nor (_18965_, _18954_, _18562_);
  and (_18976_, _18965_, _18944_);
  nor (_18987_, _18965_, _18944_);
  nor (_18998_, _18987_, _18976_);
  not (_19009_, _18998_);
  and (_19020_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19031_, _18518_, _18497_);
  nor (_19042_, _19031_, _18529_);
  and (_19053_, _19042_, _19020_);
  and (_19063_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_19074_, _18486_, _18464_);
  nor (_19085_, _19074_, _18497_);
  and (_19096_, _19085_, _19063_);
  and (_19107_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_19118_, _18453_, _18431_);
  nor (_19129_, _19118_, _18464_);
  and (_19140_, _19129_, _19107_);
  nor (_19151_, _19085_, _19063_);
  nor (_19162_, _19151_, _19096_);
  and (_19172_, _19162_, _19140_);
  nor (_19183_, _19172_, _19096_);
  not (_19194_, _19183_);
  nor (_19205_, _19042_, _19020_);
  nor (_19216_, _19205_, _19053_);
  and (_19227_, _19216_, _19194_);
  nor (_19238_, _19227_, _19053_);
  nor (_19249_, _19238_, _19009_);
  nor (_19260_, _19249_, _18976_);
  nor (_19271_, _19260_, _18933_);
  nor (_19281_, _19271_, _18900_);
  nor (_19292_, _19281_, _18856_);
  nor (_19303_, _19292_, _18824_);
  nor (_19314_, _18769_, _18747_);
  nor (_19325_, _19314_, _18780_);
  not (_19336_, _19325_);
  nor (_19347_, _19336_, _19303_);
  nor (_19358_, _19347_, _18780_);
  nor (_19369_, _19358_, _18736_);
  nor (_19380_, _19369_, _18704_);
  not (_19391_, _19380_);
  and (_19401_, _19391_, _14899_);
  and (_19412_, _19401_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_19423_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_19434_, _19423_, _19412_);
  and (_19445_, _19434_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_19456_, _19445_, _14888_);
  and (_19467_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19478_, _19467_, _19456_);
  and (_19489_, _19456_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19500_, _19489_, _19478_);
  and (_26950_, _19500_, _36029_);
  nor (_19520_, _14758_, _14790_);
  and (_19531_, _14758_, _14790_);
  or (_19542_, _19531_, _19520_);
  and (_02699_, _19542_, _36029_);
  and (_19563_, _18409_, _15676_);
  and (_02900_, _19563_, _36029_);
  nor (_19584_, _18420_, _18071_);
  nor (_19595_, _19584_, _18431_);
  and (_03104_, _19595_, _36029_);
  nor (_19615_, _19129_, _19107_);
  nor (_19626_, _19615_, _19140_);
  and (_03315_, _19626_, _36029_);
  nor (_19647_, _19162_, _19140_);
  nor (_19658_, _19647_, _19172_);
  and (_03516_, _19658_, _36029_);
  nor (_19679_, _19216_, _19194_);
  nor (_19690_, _19679_, _19227_);
  and (_03717_, _19690_, _36029_);
  and (_19711_, _19238_, _19009_);
  nor (_19721_, _19711_, _19249_);
  and (_03918_, _19721_, _36029_);
  and (_19742_, _19260_, _18933_);
  nor (_19753_, _19742_, _19271_);
  and (_04119_, _19753_, _36029_);
  and (_19774_, _19281_, _18856_);
  nor (_19785_, _19774_, _19292_);
  and (_04320_, _19785_, _36029_);
  and (_19806_, _19336_, _19303_);
  nor (_19817_, _19806_, _19347_);
  and (_04434_, _19817_, _36029_);
  and (_19837_, _19358_, _18736_);
  nor (_19848_, _19837_, _19369_);
  and (_04547_, _19848_, _36029_);
  nor (_19869_, _19391_, _14899_);
  nor (_19880_, _19869_, _19401_);
  and (_04648_, _19880_, _36029_);
  and (_19901_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_19912_, _19901_, _19401_);
  nor (_19923_, _19912_, _19412_);
  and (_04749_, _19923_, _36029_);
  nor (_19943_, _19423_, _19412_);
  nor (_19954_, _19943_, _19434_);
  and (_04850_, _19954_, _36029_);
  and (_19975_, _14877_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_19986_, _19975_, _19434_);
  nor (_19997_, _19986_, _19445_);
  and (_04951_, _19997_, _36029_);
  nor (_20018_, _19445_, _14888_);
  nor (_20029_, _20018_, _19456_);
  and (_05052_, _20029_, _36029_);
  and (_20050_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _14692_);
  nor (_20061_, _20050_, _14703_);
  not (_20072_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_20083_, _14725_, _20072_);
  and (_20094_, _20083_, _20061_);
  and (_20105_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_20116_, _20105_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20127_, _20105_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20138_, _20127_, _20116_);
  and (_01053_, _20138_, _36029_);
  and (_01083_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _36029_);
  not (_20169_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_20180_, _16459_, _20169_);
  and (_20191_, _16144_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20201_, _20191_, _20180_);
  nor (_20212_, _20201_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20223_, _16296_, _20169_);
  and (_20234_, _16634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_20245_, _20234_, _20223_);
  and (_20256_, _20245_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20267_, _20256_, _20212_);
  nor (_20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20289_, _20278_, _16795_);
  nor (_20300_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_20311_, _20300_, _20289_);
  not (_20322_, _20311_);
  and (_20333_, _15480_, _20169_);
  and (_20344_, _15151_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20355_, _20344_, _20333_);
  nor (_20366_, _20355_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20377_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20388_, _15316_, _20169_);
  and (_20399_, _15654_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20410_, _20399_, _20388_);
  nor (_20421_, _20410_, _20377_);
  nor (_20432_, _20421_, _20366_);
  nor (_20443_, _20432_, _20322_);
  and (_20454_, _20432_, _20322_);
  nor (_20465_, _20454_, _20443_);
  nor (_20476_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_20487_, _20278_, _15970_);
  nor (_20498_, _20487_, _20476_);
  not (_20509_, _20498_);
  nor (_20520_, _16459_, _20169_);
  nor (_20531_, _20520_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20542_, _16144_, _20169_);
  and (_20553_, _16296_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20564_, _20553_, _20542_);
  nor (_20575_, _20564_, _20377_);
  nor (_20586_, _20575_, _20531_);
  nor (_20597_, _20586_, _20509_);
  and (_20607_, _20586_, _20509_);
  nor (_20618_, _20607_, _20597_);
  not (_20629_, _20618_);
  nor (_20640_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_20651_, _20278_, _16991_);
  nor (_20662_, _20651_, _20640_);
  not (_20673_, _20662_);
  nor (_20684_, _15480_, _20169_);
  nor (_20695_, _20684_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20706_, _15151_, _20169_);
  and (_20717_, _15316_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20728_, _20717_, _20706_);
  nor (_20739_, _20728_, _20377_);
  nor (_20750_, _20739_, _20695_);
  nor (_20761_, _20750_, _20673_);
  and (_20772_, _20750_, _20673_);
  and (_20783_, _20201_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20794_, _20783_);
  and (_20805_, _20278_, _17166_);
  nor (_20816_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  nor (_20827_, _20816_, _20805_);
  and (_20838_, _20827_, _20794_);
  and (_20849_, _20355_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20860_, _20849_);
  and (_20871_, _20278_, _17504_);
  nor (_20882_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_20893_, _20882_, _20871_);
  and (_20904_, _20893_, _20860_);
  nor (_20915_, _20893_, _20860_);
  nor (_20926_, _20915_, _20904_);
  not (_20937_, _20926_);
  and (_20948_, _20520_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20959_, _20948_);
  and (_20969_, _20278_, _18028_);
  nor (_20980_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_20991_, _20980_, _20969_);
  and (_21002_, _20991_, _20959_);
  and (_21013_, _20684_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21024_, _21013_);
  nor (_21035_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_21046_, _20278_, _17853_);
  nor (_21057_, _21046_, _21035_);
  nor (_21068_, _21057_, _21024_);
  not (_21079_, _21068_);
  nor (_21090_, _20991_, _20959_);
  nor (_21101_, _21090_, _21002_);
  and (_21112_, _21101_, _21079_);
  nor (_21123_, _21112_, _21002_);
  nor (_21134_, _21123_, _20937_);
  nor (_21145_, _21134_, _20904_);
  nor (_21156_, _20827_, _20794_);
  nor (_21167_, _21156_, _20838_);
  not (_21178_, _21167_);
  nor (_21189_, _21178_, _21145_);
  nor (_21200_, _21189_, _20838_);
  nor (_21211_, _21200_, _20772_);
  nor (_21222_, _21211_, _20761_);
  nor (_21233_, _21222_, _20629_);
  nor (_21244_, _21233_, _20597_);
  not (_21255_, _21244_);
  and (_21266_, _21255_, _20465_);
  or (_21277_, _21266_, _20443_);
  and (_21288_, _16634_, _15654_);
  or (_21299_, _21288_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_21310_, _20564_);
  and (_21321_, _20245_, _21310_);
  nor (_21331_, _20728_, _20410_);
  and (_21342_, _21331_, _21321_);
  or (_21353_, _21342_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21364_, _21353_, _21299_);
  and (_21375_, _21364_, _21277_);
  and (_21386_, _21375_, _20267_);
  nor (_21397_, _21255_, _20465_);
  or (_21408_, _21397_, _21266_);
  and (_21419_, _21408_, _21386_);
  nor (_21430_, _21386_, _20311_);
  nor (_21441_, _21430_, _21419_);
  not (_21452_, _21441_);
  and (_21463_, _21441_, _20267_);
  not (_21474_, _20432_);
  nor (_21485_, _21386_, _20509_);
  and (_21496_, _21222_, _20629_);
  nor (_21507_, _21496_, _21233_);
  and (_21518_, _21507_, _21386_);
  or (_21529_, _21518_, _21485_);
  and (_21540_, _21529_, _21474_);
  nor (_21551_, _21529_, _21474_);
  nor (_21562_, _21551_, _21540_);
  not (_21573_, _21562_);
  not (_21584_, _20586_);
  nor (_21595_, _21386_, _20673_);
  nor (_21617_, _20772_, _20761_);
  nor (_21629_, _21617_, _21200_);
  and (_21641_, _21617_, _21200_);
  or (_21653_, _21641_, _21629_);
  and (_21665_, _21653_, _21386_);
  or (_21677_, _21665_, _21595_);
  and (_21678_, _21677_, _21584_);
  nor (_21688_, _21677_, _21584_);
  nor (_21699_, _21688_, _21678_);
  not (_21710_, _21699_);
  not (_21721_, _20750_);
  and (_21732_, _21178_, _21145_);
  or (_21743_, _21732_, _21189_);
  and (_21754_, _21743_, _21386_);
  nor (_21765_, _21386_, _20827_);
  nor (_21776_, _21765_, _21754_);
  and (_21787_, _21776_, _21721_);
  and (_21798_, _21123_, _20937_);
  nor (_21809_, _21798_, _21134_);
  not (_21820_, _21809_);
  and (_21831_, _21820_, _21386_);
  nor (_21842_, _21386_, _20893_);
  nor (_21853_, _21842_, _21831_);
  and (_21864_, _21853_, _20794_);
  nor (_21875_, _21853_, _20794_);
  nor (_21886_, _21875_, _21864_);
  not (_21897_, _21886_);
  nor (_21908_, _21101_, _21079_);
  nor (_21919_, _21908_, _21112_);
  not (_21930_, _21919_);
  and (_21941_, _21930_, _21386_);
  nor (_21952_, _21386_, _20991_);
  nor (_21963_, _21952_, _21941_);
  and (_21974_, _21963_, _20860_);
  and (_21985_, _21386_, _21013_);
  nor (_21996_, _21985_, _21057_);
  and (_22007_, _21985_, _21057_);
  nor (_22018_, _22007_, _21996_);
  and (_22029_, _22018_, _20959_);
  nor (_22040_, _22018_, _20959_);
  nor (_22051_, _22040_, _22029_);
  nor (_22061_, _20278_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_22072_, _20278_, _18398_);
  nor (_22083_, _22072_, _22061_);
  nor (_22094_, _22083_, _21024_);
  not (_22105_, _22094_);
  and (_22116_, _22105_, _22051_);
  nor (_22127_, _22116_, _22029_);
  nor (_22138_, _21963_, _20860_);
  nor (_22149_, _22138_, _21974_);
  not (_22160_, _22149_);
  nor (_22171_, _22160_, _22127_);
  nor (_22192_, _22171_, _21974_);
  nor (_22193_, _22192_, _21897_);
  nor (_22204_, _22193_, _21864_);
  nor (_22215_, _21776_, _21721_);
  nor (_22226_, _22215_, _21787_);
  not (_22237_, _22226_);
  nor (_22248_, _22237_, _22204_);
  nor (_22259_, _22248_, _21787_);
  nor (_22270_, _22259_, _21710_);
  nor (_22281_, _22270_, _21678_);
  nor (_22292_, _22281_, _21573_);
  or (_22303_, _22292_, _21540_);
  or (_22314_, _22303_, _21463_);
  and (_22325_, _22314_, _21364_);
  nor (_22336_, _22325_, _21452_);
  and (_22347_, _21463_, _21364_);
  and (_22358_, _22347_, _22303_);
  or (_22369_, _22358_, _22336_);
  and (_01090_, _22369_, _36029_);
  or (_22390_, _21441_, _20267_);
  and (_22401_, _22390_, _22325_);
  and (_03061_, _22401_, _36029_);
  and (_03072_, _21386_, _36029_);
  and (_03093_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _36029_);
  and (_03115_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _36029_);
  and (_03136_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _36029_);
  or (_22462_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_22473_, _20105_, rst);
  and (_03147_, _22473_, _22462_);
  and (_22494_, _22401_, _21013_);
  or (_22505_, _22494_, _22083_);
  nand (_22516_, _22494_, _22083_);
  and (_22527_, _22516_, _22505_);
  and (_03158_, _22527_, _36029_);
  nor (_22548_, _22105_, _22051_);
  or (_22559_, _22548_, _22116_);
  nand (_22570_, _22559_, _22401_);
  or (_22581_, _22401_, _22018_);
  and (_22592_, _22581_, _22570_);
  and (_03169_, _22592_, _36029_);
  and (_22613_, _22160_, _22127_);
  or (_22624_, _22613_, _22171_);
  nand (_22635_, _22624_, _22401_);
  or (_22646_, _22401_, _21963_);
  and (_22657_, _22646_, _22635_);
  and (_03180_, _22657_, _36029_);
  and (_22678_, _22192_, _21897_);
  or (_22689_, _22678_, _22193_);
  nand (_22700_, _22689_, _22401_);
  or (_22711_, _22401_, _21853_);
  and (_22722_, _22711_, _22700_);
  and (_03191_, _22722_, _36029_);
  and (_22743_, _22237_, _22204_);
  or (_22754_, _22743_, _22248_);
  nand (_22765_, _22754_, _22401_);
  or (_22775_, _22401_, _21776_);
  and (_22786_, _22775_, _22765_);
  and (_03202_, _22786_, _36029_);
  and (_22807_, _22259_, _21710_);
  or (_22818_, _22807_, _22270_);
  nand (_22829_, _22818_, _22401_);
  or (_22840_, _22401_, _21677_);
  and (_22851_, _22840_, _22829_);
  and (_03213_, _22851_, _36029_);
  and (_22872_, _22281_, _21573_);
  or (_22883_, _22872_, _22292_);
  nand (_22894_, _22883_, _22401_);
  or (_22905_, _22401_, _21529_);
  and (_22916_, _22905_, _22894_);
  and (_03224_, _22916_, _36029_);
  and (_22937_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_22948_, _22937_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22959_, _22948_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22970_, _22959_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22981_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22992_, _22981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_23003_, _22992_);
  not (_23014_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23025_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _14692_);
  and (_23036_, _23025_, _23014_);
  and (_23047_, _23036_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_23058_, _23047_);
  nor (_23069_, _22981_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23080_, _23069_, _23058_);
  and (_23091_, _23080_, _23003_);
  not (_23102_, _23091_);
  and (_23122_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23123_, _23122_, _23025_);
  not (_23134_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_23155_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _14692_);
  and (_23156_, _23155_, _23134_);
  and (_23167_, _23156_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23188_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_23189_, _23188_, _23123_);
  not (_23200_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23221_, _23036_, _23200_);
  and (_23222_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23233_, _23156_, _23014_);
  and (_23254_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_23255_, _23254_, _23222_);
  and (_23266_, _23255_, _23189_);
  and (_23287_, _23266_, _23102_);
  not (_23288_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_23299_, _22992_, _23288_);
  and (_23320_, _22992_, _23288_);
  nor (_23321_, _23320_, _23299_);
  nor (_23332_, _23321_, _23058_);
  not (_23343_, _23332_);
  and (_23354_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_23365_, _23354_, _23123_);
  and (_23376_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_23387_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_23398_, _23387_, _23376_);
  and (_23409_, _23398_, _23365_);
  and (_23420_, _23409_, _23343_);
  nor (_23431_, _23420_, _23287_);
  and (_23442_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_23452_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_23463_, _23452_, _23442_);
  not (_23474_, _22959_);
  nor (_23485_, _22948_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_23496_, _23485_, _23058_);
  and (_23507_, _23496_, _23474_);
  or (_23518_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23529_, _23518_, _14692_);
  nor (_23540_, _23529_, _23155_);
  and (_23551_, _23540_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_23562_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_23573_, _23562_, _23551_);
  not (_23584_, _23573_);
  nor (_23595_, _23584_, _23507_);
  and (_23606_, _23595_, _23463_);
  nor (_23617_, _22959_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_23628_, _23617_);
  nor (_23639_, _23058_, _22970_);
  and (_23650_, _23639_, _23628_);
  not (_23661_, _23650_);
  and (_23672_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_23683_, _23672_, _23123_);
  and (_23694_, _23540_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_23705_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_23716_, _23705_, _23694_);
  and (_23727_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  not (_23738_, _23727_);
  and (_23749_, _23738_, _23716_);
  and (_23759_, _23749_, _23683_);
  and (_23770_, _23759_, _23661_);
  not (_23781_, _23770_);
  and (_23792_, _23781_, _23606_);
  nor (_23803_, _22970_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_23814_, _23803_);
  nor (_23825_, _23058_, _22981_);
  and (_23836_, _23825_, _23814_);
  not (_23847_, _23836_);
  and (_23858_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_23869_, _23858_, _23123_);
  and (_23880_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_23891_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_23902_, _23891_, _23880_);
  and (_23913_, _23902_, _23869_);
  and (_23924_, _23913_, _23847_);
  not (_23935_, _23924_);
  and (_23946_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_23957_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_23968_, _23957_, _23946_);
  and (_23979_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_23990_, _23979_);
  not (_24001_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24012_, _23047_, _24001_);
  and (_24023_, _23540_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24034_, _24023_, _24012_);
  and (_24045_, _24034_, _23990_);
  and (_24056_, _24045_, _23968_);
  nor (_24067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24078_, _24067_, _22937_);
  and (_24088_, _24078_, _23047_);
  and (_24099_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  nor (_24110_, _24099_, _24088_);
  and (_24121_, _23540_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  not (_24132_, _24121_);
  and (_24143_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24154_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24165_, _24154_, _24143_);
  and (_24176_, _24165_, _24132_);
  and (_24187_, _24176_, _24110_);
  nor (_24198_, _22937_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24209_, _24198_, _22948_);
  and (_24220_, _24209_, _23047_);
  and (_24231_, _23221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24242_, _24231_, _24220_);
  and (_24253_, _23167_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24264_, _23233_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_24275_, _23540_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24286_, _24275_, _24264_);
  nor (_24297_, _24286_, _24253_);
  and (_24319_, _24297_, _24242_);
  and (_24331_, _24319_, _24187_);
  and (_24343_, _24331_, _24056_);
  and (_24355_, _24343_, _23935_);
  and (_24367_, _24355_, _23792_);
  nand (_24379_, _24367_, _23431_);
  and (_24391_, _22369_, _20094_);
  not (_24392_, _24391_);
  and (_24403_, _19500_, _14758_);
  not (_24414_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_24424_, _14703_, _24414_);
  and (_24435_, _24424_, _14747_);
  not (_24446_, _24435_);
  nor (_24457_, _16795_, _16634_);
  and (_24468_, _16795_, _16634_);
  nor (_24479_, _24468_, _24457_);
  not (_24490_, _15654_);
  nor (_24501_, _15970_, _24490_);
  nor (_24512_, _15970_, _15654_);
  and (_24523_, _15970_, _15654_);
  nor (_24534_, _24523_, _24512_);
  not (_24545_, _16296_);
  nor (_24556_, _16991_, _24545_);
  nor (_24567_, _16991_, _16296_);
  and (_24578_, _16991_, _16296_);
  nor (_24589_, _24578_, _24567_);
  not (_24600_, _15316_);
  and (_24611_, _17166_, _24600_);
  nor (_24622_, _24611_, _24589_);
  nor (_24633_, _24622_, _24556_);
  nor (_24644_, _24633_, _24534_);
  nor (_24655_, _24644_, _24501_);
  and (_24666_, _24633_, _24534_);
  nor (_24677_, _24666_, _24644_);
  not (_24688_, _24677_);
  and (_24699_, _24611_, _24589_);
  nor (_24710_, _24699_, _24622_);
  not (_24721_, _24710_);
  nor (_24732_, _17166_, _15316_);
  and (_24743_, _17166_, _15316_);
  nor (_24754_, _24743_, _24732_);
  not (_24765_, _24754_);
  and (_24776_, _17504_, _16144_);
  nor (_24787_, _17504_, _16144_);
  nor (_24798_, _24787_, _24776_);
  nor (_24809_, _18028_, _15151_);
  and (_24820_, _18028_, _15151_);
  nor (_24831_, _24820_, _24809_);
  nor (_24842_, _17853_, _16459_);
  and (_24853_, _17853_, _16459_);
  nor (_24864_, _24853_, _24842_);
  not (_24875_, _15480_);
  and (_24886_, _18398_, _24875_);
  nor (_24897_, _24886_, _24864_);
  not (_24908_, _16459_);
  nor (_24919_, _17853_, _24908_);
  nor (_24930_, _24919_, _24897_);
  nor (_24941_, _24930_, _24831_);
  not (_24952_, _15151_);
  nor (_24963_, _18028_, _24952_);
  nor (_24974_, _24963_, _24941_);
  nor (_24985_, _24974_, _24798_);
  and (_24996_, _24974_, _24798_);
  nor (_25007_, _24996_, _24985_);
  not (_25018_, _25007_);
  and (_25029_, _24930_, _24831_);
  nor (_25040_, _25029_, _24941_);
  not (_25051_, _25040_);
  and (_25061_, _24886_, _24864_);
  nor (_25072_, _25061_, _24897_);
  not (_25083_, _25072_);
  nor (_25094_, _18398_, _15480_);
  and (_25105_, _18398_, _15480_);
  nor (_25116_, _25105_, _25094_);
  not (_25127_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_25138_, _14965_, _25127_);
  not (_25149_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_25160_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25171_, _25160_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25182_, _25171_, _15545_);
  nor (_25193_, _25182_, _25149_);
  nor (_25204_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25215_, _25204_, _15206_);
  not (_25226_, _25215_);
  and (_25247_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25248_, _25247_, _16525_);
  not (_25259_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25270_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25259_);
  and (_25291_, _25270_, _16187_);
  nor (_25292_, _25291_, _25248_);
  and (_25303_, _25292_, _25226_);
  and (_25324_, _25303_, _25193_);
  and (_25325_, _25171_, _15009_);
  nor (_25336_, _25325_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25347_, _25270_, _16351_);
  not (_25358_, _25347_);
  and (_25379_, _25247_, _16035_);
  and (_25380_, _25204_, _15371_);
  nor (_25391_, _25380_, _25379_);
  and (_25402_, _25391_, _25358_);
  and (_25413_, _25402_, _25336_);
  nor (_25424_, _25413_, _25324_);
  nor (_25435_, _25424_, _14965_);
  nor (_25446_, _25435_, _25138_);
  and (_25457_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25468_, _25457_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_25479_, _25468_);
  and (_25490_, _25479_, _25446_);
  and (_25511_, _25479_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_25512_, _25511_, _25490_);
  nor (_25523_, _25512_, _25116_);
  and (_25534_, _25523_, _25083_);
  and (_25545_, _25534_, _25051_);
  and (_25556_, _25545_, _25018_);
  not (_25567_, _16144_);
  or (_25578_, _17504_, _25567_);
  and (_25589_, _17504_, _25567_);
  or (_25600_, _24974_, _25589_);
  and (_25611_, _25600_, _25578_);
  or (_25622_, _25611_, _25556_);
  and (_25633_, _25622_, _24765_);
  and (_25644_, _25633_, _24721_);
  and (_25655_, _25644_, _24688_);
  nor (_25666_, _25655_, _24655_);
  nor (_25687_, _25666_, _24479_);
  and (_25688_, _25666_, _24479_);
  nor (_25699_, _25688_, _25687_);
  nor (_25710_, _25699_, _24446_);
  not (_25721_, _25710_);
  not (_25732_, _24479_);
  not (_25743_, _24534_);
  and (_25754_, _24732_, _24589_);
  nor (_25765_, _25754_, _24567_);
  nor (_25776_, _25765_, _25743_);
  not (_25787_, _24831_);
  and (_25798_, _25094_, _24864_);
  nor (_25809_, _25798_, _24842_);
  nor (_25820_, _25809_, _25787_);
  nor (_25831_, _25820_, _24809_);
  nor (_25842_, _25831_, _24798_);
  and (_25853_, _25831_, _24798_);
  nor (_25864_, _25853_, _25842_);
  not (_25885_, _25116_);
  nor (_25886_, _25512_, _25885_);
  and (_25897_, _25886_, _24864_);
  and (_25908_, _25809_, _25787_);
  nor (_25919_, _25908_, _25820_);
  and (_25930_, _25919_, _25897_);
  not (_25941_, _25930_);
  nor (_25952_, _25941_, _25864_);
  nor (_25963_, _25831_, _24776_);
  or (_25974_, _25963_, _24787_);
  or (_25985_, _25974_, _25952_);
  and (_25996_, _25985_, _24754_);
  nor (_26007_, _24732_, _24589_);
  nor (_26018_, _26007_, _25754_);
  and (_26029_, _26018_, _25996_);
  and (_26040_, _25765_, _25743_);
  nor (_26051_, _26040_, _25776_);
  and (_26062_, _26051_, _26029_);
  or (_26073_, _26062_, _25776_);
  nor (_26084_, _26073_, _24512_);
  and (_26095_, _26084_, _25732_);
  nor (_26106_, _26084_, _25732_);
  not (_26117_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_26128_, _20050_, _26117_);
  and (_26139_, _26128_, _14747_);
  not (_26150_, _26139_);
  or (_26161_, _26150_, _26106_);
  nor (_26172_, _26161_, _26095_);
  and (_26183_, _14736_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26194_, _26183_, _24424_);
  nor (_26205_, _18398_, _17853_);
  and (_26216_, _26205_, _18039_);
  and (_26237_, _26216_, _17515_);
  and (_26238_, _26237_, _17177_);
  and (_26249_, _26238_, _17002_);
  and (_26260_, _26249_, _15981_);
  and (_26271_, _26260_, _25512_);
  not (_26282_, _25512_);
  and (_26293_, _15970_, _16991_);
  and (_26304_, _18398_, _17853_);
  and (_26315_, _26304_, _18028_);
  and (_26326_, _26315_, _17504_);
  and (_26347_, _26326_, _17166_);
  and (_26348_, _26347_, _26293_);
  and (_26359_, _26348_, _26282_);
  nor (_26370_, _26359_, _26271_);
  and (_26381_, _26370_, _16795_);
  nor (_26392_, _26370_, _16795_);
  nor (_26403_, _26392_, _26381_);
  and (_26414_, _26403_, _26194_);
  not (_26425_, _16634_);
  nor (_26436_, _25512_, _26425_);
  not (_26447_, _26436_);
  and (_26458_, _25512_, _16795_);
  and (_26469_, _26183_, _14714_);
  not (_26480_, _26469_);
  nor (_26491_, _26480_, _26458_);
  and (_26502_, _26491_, _26447_);
  nor (_26513_, _26502_, _26414_);
  and (_26524_, _26128_, _20083_);
  and (_26535_, _18028_, _17853_);
  nor (_26546_, _26535_, _17504_);
  and (_26556_, _26546_, _26524_);
  and (_26567_, _26556_, _17177_);
  not (_26578_, _26567_);
  and (_26589_, _26578_, _26293_);
  nor (_26600_, _26293_, _16795_);
  nor (_26611_, _26600_, _26556_);
  and (_26622_, _26611_, _25512_);
  nor (_26633_, _26622_, _26589_);
  nor (_26644_, _26633_, _16806_);
  and (_26655_, _26633_, _16806_);
  nor (_26665_, _26655_, _26644_);
  and (_26676_, _26665_, _26524_);
  and (_26687_, _26183_, _26128_);
  not (_26698_, _26687_);
  nor (_26709_, _26698_, _25512_);
  not (_26720_, _26709_);
  not (_26731_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26742_, _14736_, _26731_);
  and (_26753_, _26742_, _26128_);
  not (_26764_, _26753_);
  nor (_26775_, _26764_, _24468_);
  and (_26796_, _26742_, _20061_);
  and (_26797_, _26796_, _24479_);
  nor (_26808_, _26797_, _26775_);
  and (_26819_, _20083_, _14714_);
  and (_26830_, _26819_, _24457_);
  and (_26841_, _24424_, _20083_);
  and (_26852_, _26841_, _16795_);
  nor (_26863_, _26852_, _26830_);
  and (_26874_, _26742_, _14703_);
  not (_26885_, _26874_);
  nor (_26896_, _26885_, _15970_);
  not (_26907_, _26896_);
  and (_26917_, _20061_, _14747_);
  not (_26928_, _26917_);
  nor (_26939_, _26928_, _16795_);
  and (_26951_, _26183_, _20061_);
  not (_26962_, _26951_);
  nor (_26973_, _26962_, _18398_);
  nor (_26984_, _26973_, _26939_);
  and (_26995_, _26984_, _26907_);
  and (_27006_, _26995_, _26863_);
  and (_27017_, _27006_, _26808_);
  and (_27027_, _27017_, _26720_);
  not (_27038_, _27027_);
  nor (_27049_, _27038_, _26676_);
  and (_27060_, _27049_, _26513_);
  not (_27071_, _27060_);
  nor (_27092_, _27071_, _26172_);
  and (_27093_, _27092_, _25721_);
  not (_27104_, _27093_);
  nor (_27115_, _27104_, _24403_);
  and (_27126_, _27115_, _24392_);
  not (_27137_, _27126_);
  or (_27147_, _27137_, _24379_);
  not (_27158_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_27169_, \oc8051_top_1.oc8051_decoder1.wr , _14692_);
  not (_27180_, _27169_);
  nor (_27201_, _27180_, _23036_);
  and (_27202_, _27201_, _27158_);
  not (_27213_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_27224_, _24379_, _27213_);
  and (_27235_, _27224_, _27202_);
  and (_27246_, _27235_, _27147_);
  nor (_27256_, _27201_, _27213_);
  nor (_27267_, _26106_, _24457_);
  nor (_27278_, _27267_, _26150_);
  not (_27289_, _27278_);
  and (_27300_, _16795_, _26425_);
  nor (_27311_, _27300_, _25687_);
  nor (_27322_, _27311_, _24446_);
  nor (_27333_, _26567_, _17002_);
  and (_27344_, _25512_, _15970_);
  and (_27355_, _27344_, _27333_);
  nor (_27366_, _27355_, _26458_);
  not (_27377_, _26524_);
  nor (_27388_, _25512_, _16795_);
  not (_27399_, _27388_);
  nor (_27420_, _27399_, _26589_);
  nor (_27421_, _27420_, _27377_);
  and (_27432_, _27421_, _27366_);
  or (_27441_, _27432_, _26556_);
  nor (_27442_, _25511_, _25446_);
  not (_27443_, _26796_);
  nor (_27454_, _27443_, _25490_);
  not (_27465_, _27454_);
  nor (_27476_, _26962_, _25446_);
  nor (_27487_, _27476_, _26753_);
  and (_27498_, _27487_, _27465_);
  nor (_27509_, _27498_, _27442_);
  not (_27520_, _27509_);
  nor (_27530_, _26928_, _25512_);
  nor (_27541_, _26698_, _18398_);
  and (_27552_, _26742_, _14714_);
  not (_27563_, _27552_);
  nor (_27574_, _27563_, _16795_);
  nor (_27585_, _27574_, _27541_);
  not (_27596_, _27585_);
  nor (_27607_, _27596_, _27530_);
  and (_27618_, _26841_, _25512_);
  and (_27629_, _25468_, _25446_);
  and (_27640_, _26742_, _24424_);
  and (_27660_, _26819_, _25446_);
  nor (_27661_, _27660_, _27640_);
  nor (_27672_, _27661_, _27629_);
  nor (_27683_, _27672_, _27618_);
  and (_27694_, _27683_, _27607_);
  and (_27705_, _27694_, _27520_);
  not (_27716_, _27705_);
  nor (_27727_, _27716_, _27441_);
  not (_27738_, _27727_);
  nor (_27749_, _27738_, _27322_);
  and (_27760_, _27749_, _27289_);
  nor (_27771_, _23924_, _23287_);
  not (_27781_, _23420_);
  and (_27792_, _23792_, _27781_);
  and (_27803_, _27792_, _27771_);
  not (_27814_, _24056_);
  nor (_27825_, _24319_, _24187_);
  and (_27836_, _27825_, _27814_);
  and (_27847_, _27836_, _27803_);
  nand (_27858_, _27847_, _27760_);
  and (_27869_, _27201_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_27880_, _27847_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_27891_, _27880_, _27869_);
  and (_27901_, _27891_, _27858_);
  or (_27912_, _27901_, _27256_);
  or (_27923_, _27912_, _27246_);
  and (_06742_, _27923_, _36029_);
  and (_27944_, _22527_, _20094_);
  not (_27955_, _27944_);
  and (_27966_, _19817_, _14758_);
  and (_27977_, _25512_, _25885_);
  nor (_27988_, _27977_, _25886_);
  nor (_27999_, _26139_, _24435_);
  not (_28010_, _27999_);
  and (_28021_, _28010_, _27988_);
  not (_28031_, _28021_);
  nor (_28042_, _27563_, _25512_);
  not (_28053_, _28042_);
  nor (_28064_, _27443_, _25094_);
  nor (_28075_, _28064_, _26753_);
  or (_28086_, _28075_, _25105_);
  and (_28097_, _26183_, _26117_);
  not (_28108_, _28097_);
  nor (_28119_, _28108_, _17853_);
  and (_28130_, _27640_, _16806_);
  nor (_28141_, _28130_, _28119_);
  and (_28152_, _26819_, _25094_);
  and (_28163_, _26841_, _18398_);
  nor (_28173_, _28163_, _28152_);
  nor (_28184_, _26480_, _15480_);
  and (_28195_, _26194_, _18398_);
  nor (_28206_, _28195_, _28184_);
  nor (_28217_, _26917_, _26524_);
  nor (_28228_, _28217_, _18398_);
  not (_28239_, _28228_);
  and (_28250_, _28239_, _28206_);
  and (_28261_, _28250_, _28173_);
  and (_28272_, _28261_, _28141_);
  and (_28283_, _28272_, _28086_);
  and (_28294_, _28283_, _28053_);
  and (_28299_, _28294_, _28031_);
  not (_28300_, _28299_);
  nor (_28301_, _28300_, _27966_);
  and (_28302_, _28301_, _27955_);
  not (_28305_, _28302_);
  or (_28313_, _28305_, _24379_);
  not (_28327_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_28328_, _24379_, _28327_);
  and (_28336_, _28328_, _27202_);
  and (_28344_, _28336_, _28313_);
  nor (_28351_, _27201_, _28327_);
  not (_28359_, _27760_);
  or (_28367_, _28359_, _24379_);
  and (_28368_, _28328_, _27869_);
  and (_28369_, _28368_, _28367_);
  or (_28371_, _28369_, _28351_);
  or (_28382_, _28371_, _28344_);
  and (_08973_, _28382_, _36029_);
  and (_28403_, _19848_, _14758_);
  not (_28413_, _28403_);
  and (_28424_, _22592_, _20094_);
  nor (_28435_, _25094_, _24864_);
  or (_28440_, _28435_, _25798_);
  and (_28461_, _28440_, _25886_);
  nor (_28462_, _28440_, _25886_);
  or (_28473_, _28462_, _28461_);
  and (_28484_, _28473_, _26139_);
  nor (_28495_, _25523_, _25083_);
  nor (_28506_, _28495_, _25534_);
  nor (_28517_, _28506_, _24446_);
  not (_28528_, _28517_);
  nor (_28539_, _26546_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_28550_, _28539_, _17864_);
  nor (_28561_, _28539_, _17864_);
  nor (_28572_, _28561_, _28550_);
  nor (_28583_, _28572_, _27377_);
  not (_28594_, _28583_);
  and (_28605_, _26796_, _24864_);
  not (_28616_, _28605_);
  nor (_28627_, _26764_, _24853_);
  not (_28638_, _28627_);
  and (_28649_, _26819_, _24842_);
  and (_28660_, _26841_, _17853_);
  nor (_28671_, _28660_, _28649_);
  and (_28682_, _28671_, _28638_);
  and (_28703_, _28682_, _28616_);
  nor (_28715_, _26885_, _18398_);
  not (_28726_, _28715_);
  nor (_28736_, _26928_, _17853_);
  nor (_28747_, _28108_, _18028_);
  nor (_28758_, _28747_, _28736_);
  and (_28768_, _28758_, _28726_);
  and (_28779_, _28768_, _28703_);
  and (_28790_, _28779_, _28594_);
  and (_28800_, _28790_, _28528_);
  nor (_28811_, _26480_, _16459_);
  nor (_28822_, _26304_, _26205_);
  not (_28833_, _28822_);
  nor (_28843_, _28833_, _25512_);
  and (_28854_, _28833_, _25512_);
  nor (_28865_, _28854_, _28843_);
  and (_28875_, _28865_, _26194_);
  nor (_28886_, _28875_, _28811_);
  nand (_28897_, _28886_, _28800_);
  nor (_28907_, _28897_, _28484_);
  not (_28918_, _28907_);
  nor (_28929_, _28918_, _28424_);
  and (_28939_, _28929_, _28413_);
  not (_28950_, _28939_);
  or (_28961_, _28950_, _24379_);
  not (_28972_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_28983_, _24379_, _28972_);
  and (_29004_, _28983_, _27202_);
  and (_29005_, _29004_, _28961_);
  nor (_29016_, _27201_, _28972_);
  and (_29027_, _24331_, _27814_);
  and (_29038_, _29027_, _27803_);
  or (_29049_, _29038_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29060_, _29049_, _27869_);
  nand (_29071_, _29038_, _27760_);
  and (_29082_, _29071_, _29060_);
  or (_29093_, _29082_, _29016_);
  or (_29104_, _29093_, _29005_);
  and (_08984_, _29104_, _36029_);
  and (_29125_, _22657_, _20094_);
  not (_29136_, _29125_);
  and (_29147_, _19880_, _14758_);
  nor (_29158_, _26480_, _15151_);
  and (_29169_, _26205_, _25512_);
  and (_29180_, _26304_, _26282_);
  nor (_29191_, _29180_, _29169_);
  and (_29202_, _29191_, _18028_);
  nor (_29213_, _29191_, _18028_);
  nor (_29224_, _29213_, _29202_);
  and (_29235_, _29224_, _26194_);
  nor (_29246_, _29235_, _29158_);
  nor (_29257_, _25534_, _25051_);
  nor (_29268_, _29257_, _25545_);
  nor (_29279_, _29268_, _24446_);
  nor (_29290_, _28108_, _17504_);
  and (_29301_, _26819_, _24809_);
  and (_29312_, _26841_, _18028_);
  nor (_29323_, _29312_, _29301_);
  nor (_29334_, _26764_, _24820_);
  and (_29345_, _26796_, _24831_);
  nor (_29356_, _29345_, _29334_);
  nor (_29367_, _26885_, _17853_);
  nor (_29378_, _26928_, _18028_);
  nor (_29389_, _29378_, _29367_);
  and (_29400_, _29389_, _29356_);
  nand (_29411_, _29400_, _29323_);
  nor (_29422_, _29411_, _29290_);
  not (_29433_, _29422_);
  nor (_29444_, _29433_, _29279_);
  nor (_29455_, _25919_, _25897_);
  nor (_29466_, _29455_, _26150_);
  and (_29477_, _29466_, _25941_);
  nor (_29488_, _28561_, _18028_);
  and (_29498_, _26535_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_29509_, _29498_, _29488_);
  nor (_29520_, _29509_, _27377_);
  nor (_29531_, _29520_, _29477_);
  and (_29551_, _29531_, _29444_);
  and (_29552_, _29551_, _29246_);
  not (_29563_, _29552_);
  nor (_29573_, _29563_, _29147_);
  and (_29584_, _29573_, _29136_);
  not (_29595_, _29584_);
  or (_29605_, _29595_, _24379_);
  not (_29616_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_29627_, _24379_, _29616_);
  and (_29637_, _29627_, _27202_);
  and (_29648_, _29637_, _29605_);
  nor (_29659_, _27201_, _29616_);
  nor (_29670_, _24187_, _24056_);
  nand (_29681_, _24319_, _27803_);
  or (_29692_, _29681_, _29670_);
  and (_29703_, _29692_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_29704_, _24187_);
  and (_29705_, _24319_, _29704_);
  and (_29706_, _29705_, _24056_);
  and (_29707_, _29706_, _28359_);
  and (_29708_, _24331_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_29709_, _29708_, _29707_);
  and (_29710_, _29709_, _27803_);
  or (_29711_, _29710_, _29703_);
  and (_29712_, _29711_, _27869_);
  or (_29713_, _29712_, _29659_);
  or (_29714_, _29713_, _29648_);
  and (_08995_, _29714_, _36029_);
  and (_29715_, _19923_, _14758_);
  not (_29716_, _29715_);
  and (_29717_, _22722_, _20094_);
  nor (_29718_, _25545_, _25018_);
  nor (_29719_, _29718_, _25556_);
  nor (_29720_, _29719_, _24446_);
  not (_29721_, _29720_);
  nor (_29722_, _26764_, _24776_);
  and (_29723_, _26796_, _24798_);
  nor (_29724_, _29723_, _29722_);
  and (_29725_, _25941_, _25864_);
  or (_29726_, _29725_, _26150_);
  nor (_29727_, _29726_, _25952_);
  nor (_29728_, _26480_, _16144_);
  nor (_29729_, _26315_, _25512_);
  nor (_29730_, _26216_, _26282_);
  nor (_29731_, _29730_, _29729_);
  and (_29732_, _29731_, _17515_);
  not (_29733_, _26194_);
  nor (_29734_, _29731_, _17515_);
  or (_29735_, _29734_, _29733_);
  nor (_29736_, _29735_, _29732_);
  nor (_29737_, _29736_, _29728_);
  nor (_29738_, _26885_, _18028_);
  nor (_29739_, _26928_, _17504_);
  nor (_29740_, _29739_, _29738_);
  not (_29741_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_29742_, _26535_, _29741_);
  nor (_29743_, _29742_, _17515_);
  or (_29744_, _29743_, _27377_);
  nor (_29745_, _29744_, _26546_);
  and (_29746_, _26819_, _24787_);
  and (_29747_, _26841_, _17504_);
  nor (_29748_, _29747_, _29746_);
  nor (_29749_, _28108_, _17166_);
  not (_29750_, _29749_);
  nand (_29751_, _29750_, _29748_);
  nor (_29752_, _29751_, _29745_);
  and (_29753_, _29752_, _29740_);
  nand (_29754_, _29753_, _29737_);
  nor (_29755_, _29754_, _29727_);
  and (_29756_, _29755_, _29724_);
  and (_29757_, _29756_, _29721_);
  not (_29758_, _29757_);
  nor (_29759_, _29758_, _29717_);
  and (_29760_, _29759_, _29716_);
  not (_29761_, _29760_);
  or (_29762_, _29761_, _24379_);
  not (_29763_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_29764_, _24379_, _29763_);
  and (_29765_, _29764_, _27202_);
  and (_29766_, _29765_, _29762_);
  nor (_29767_, _27201_, _29763_);
  and (_29768_, _29681_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_29769_, _29670_, _24319_);
  and (_29770_, _29769_, _28359_);
  not (_29771_, _24319_);
  or (_29772_, _29670_, _29771_);
  nor (_29773_, _29772_, _29763_);
  or (_29774_, _29773_, _29770_);
  and (_29775_, _29774_, _27803_);
  or (_29776_, _29775_, _29768_);
  and (_29777_, _29776_, _27869_);
  or (_29778_, _29777_, _29767_);
  or (_29779_, _29778_, _29766_);
  and (_09006_, _29779_, _36029_);
  and (_29780_, _22786_, _20094_);
  not (_29781_, _29780_);
  and (_29782_, _19954_, _14758_);
  nor (_29783_, _25622_, _24754_);
  and (_29784_, _25622_, _24754_);
  nor (_29785_, _29784_, _29783_);
  and (_29786_, _29785_, _24435_);
  not (_29787_, _29786_);
  nor (_29788_, _25985_, _24754_);
  nor (_29789_, _29788_, _25996_);
  and (_29790_, _29789_, _26139_);
  not (_29791_, _29790_);
  nor (_29792_, _26556_, _17177_);
  nor (_29793_, _29792_, _27377_);
  and (_29794_, _29793_, _26578_);
  not (_29795_, _29794_);
  and (_29796_, _26237_, _25512_);
  and (_29797_, _26326_, _26282_);
  nor (_29798_, _29797_, _29796_);
  nor (_29799_, _29798_, _17166_);
  not (_29800_, _29799_);
  and (_29801_, _29798_, _17166_);
  nor (_29802_, _29801_, _29733_);
  and (_29803_, _29802_, _29800_);
  and (_29804_, _25512_, _17177_);
  nor (_29805_, _25512_, _15316_);
  or (_29806_, _29805_, _29804_);
  and (_29807_, _29806_, _26469_);
  nor (_29808_, _29807_, _29803_);
  and (_29809_, _26819_, _24732_);
  and (_29810_, _26841_, _17166_);
  nor (_29811_, _29810_, _29809_);
  nor (_29812_, _28108_, _16991_);
  not (_29813_, _29812_);
  and (_29814_, _29813_, _29811_);
  and (_29815_, _26796_, _24754_);
  nor (_29816_, _26764_, _24743_);
  or (_29817_, _29816_, _29815_);
  nor (_29818_, _26928_, _17166_);
  nor (_29819_, _26885_, _17504_);
  nor (_29820_, _29819_, _29818_);
  not (_29821_, _29820_);
  nor (_29822_, _29821_, _29817_);
  and (_29823_, _29822_, _29814_);
  and (_29824_, _29823_, _29808_);
  and (_29825_, _29824_, _29795_);
  and (_29826_, _29825_, _29791_);
  and (_29827_, _29826_, _29787_);
  not (_29828_, _29827_);
  nor (_29829_, _29828_, _29782_);
  and (_29830_, _29829_, _29781_);
  not (_29831_, _29830_);
  or (_29832_, _29831_, _24379_);
  not (_29833_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_29834_, _24379_, _29833_);
  and (_29835_, _29834_, _27202_);
  and (_29836_, _29835_, _29832_);
  nor (_29837_, _27201_, _29833_);
  not (_29838_, _27803_);
  and (_29839_, _24187_, _24056_);
  and (_29840_, _29839_, _29771_);
  nor (_29841_, _29839_, _29771_);
  nor (_29842_, _29841_, _29840_);
  or (_29843_, _29842_, _29838_);
  and (_29844_, _29843_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_29845_, _29840_, _28359_);
  and (_29846_, _29841_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_29847_, _29846_, _29845_);
  and (_29848_, _29847_, _27803_);
  or (_29849_, _29848_, _29844_);
  and (_29850_, _29849_, _27869_);
  or (_29851_, _29850_, _29837_);
  or (_29852_, _29851_, _29836_);
  and (_09017_, _29852_, _36029_);
  and (_29853_, _22851_, _20094_);
  not (_29854_, _29853_);
  and (_29855_, _19997_, _14758_);
  nor (_29856_, _26018_, _25996_);
  nor (_29857_, _29856_, _26029_);
  and (_29858_, _29857_, _26139_);
  not (_29859_, _29858_);
  nor (_29860_, _25633_, _24721_);
  nor (_29861_, _29860_, _25644_);
  nor (_29862_, _29861_, _24446_);
  nor (_29863_, _25512_, _16296_);
  and (_29864_, _25512_, _17002_);
  nor (_29865_, _29864_, _29863_);
  nor (_29866_, _29865_, _26480_);
  nor (_29867_, _26238_, _26282_);
  nor (_29868_, _26347_, _25512_);
  nor (_29869_, _29868_, _29867_);
  and (_29870_, _29869_, _17002_);
  not (_29871_, _29870_);
  nor (_29872_, _29869_, _17002_);
  nor (_29873_, _29872_, _29733_);
  and (_29874_, _29873_, _29871_);
  nor (_29875_, _29874_, _29866_);
  not (_29876_, _26622_);
  and (_29877_, _29876_, _27333_);
  nor (_29878_, _26622_, _26567_);
  nor (_29879_, _29878_, _16991_);
  nor (_29880_, _29879_, _29877_);
  nor (_29881_, _29880_, _27377_);
  and (_29882_, _26796_, _24589_);
  and (_29883_, _26819_, _24567_);
  nor (_29884_, _26764_, _24578_);
  and (_29885_, _26841_, _16991_);
  or (_29886_, _29885_, _29884_);
  or (_29887_, _29886_, _29883_);
  nor (_29888_, _29887_, _29882_);
  nor (_29889_, _28108_, _15970_);
  nor (_29890_, _26928_, _16991_);
  nor (_29891_, _26885_, _17166_);
  or (_29892_, _29891_, _29890_);
  nor (_29893_, _29892_, _29889_);
  and (_29894_, _29893_, _29888_);
  not (_29895_, _29894_);
  nor (_29896_, _29895_, _29881_);
  and (_29897_, _29896_, _29875_);
  not (_29898_, _29897_);
  nor (_29899_, _29898_, _29862_);
  and (_29900_, _29899_, _29859_);
  not (_29901_, _29900_);
  nor (_29902_, _29901_, _29855_);
  and (_29903_, _29902_, _29854_);
  not (_29904_, _29903_);
  or (_29905_, _29904_, _24379_);
  not (_29906_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_29907_, _24379_, _29906_);
  and (_29908_, _29907_, _27202_);
  and (_29909_, _29908_, _29905_);
  nor (_29910_, _27201_, _29906_);
  and (_29911_, _29771_, _24187_);
  nor (_29912_, _29911_, _29705_);
  or (_29913_, _29912_, _29838_);
  and (_29914_, _29913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_29915_, _24187_, _27814_);
  and (_29916_, _29915_, _29771_);
  and (_29917_, _29916_, _28359_);
  or (_29918_, _29840_, _29705_);
  and (_29919_, _29918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_29920_, _29919_, _29917_);
  and (_29921_, _29920_, _27803_);
  or (_29922_, _29921_, _29914_);
  and (_29923_, _29922_, _27869_);
  or (_29924_, _29923_, _29910_);
  or (_29925_, _29924_, _29909_);
  and (_09028_, _29925_, _36029_);
  and (_29926_, _22916_, _20094_);
  not (_29927_, _29926_);
  and (_29928_, _20029_, _14758_);
  nor (_29929_, _26051_, _26029_);
  not (_29930_, _29929_);
  nor (_29931_, _26150_, _26062_);
  and (_29932_, _29931_, _29930_);
  not (_29933_, _29932_);
  nor (_29934_, _25644_, _24688_);
  nor (_29935_, _29934_, _25655_);
  nor (_29936_, _29935_, _24446_);
  nor (_29937_, _25512_, _24490_);
  or (_29938_, _29937_, _26480_);
  nor (_29939_, _29938_, _27344_);
  nor (_29940_, _25512_, _17002_);
  nand (_29941_, _29940_, _26347_);
  nand (_29942_, _26249_, _25512_);
  and (_29943_, _29942_, _29941_);
  and (_29944_, _29943_, _15970_);
  nor (_29945_, _29943_, _15970_);
  or (_29946_, _29945_, _29733_);
  nor (_29947_, _29946_, _29944_);
  nor (_29948_, _29947_, _29939_);
  nor (_29949_, _29877_, _15970_);
  and (_29950_, _29877_, _15970_);
  nor (_29951_, _29950_, _29949_);
  nor (_29952_, _29951_, _27377_);
  and (_29953_, _26796_, _24534_);
  nor (_29954_, _26764_, _24523_);
  not (_29955_, _29954_);
  and (_29956_, _26819_, _24512_);
  and (_29957_, _26841_, _15970_);
  nor (_29958_, _29957_, _29956_);
  nand (_29959_, _29958_, _29955_);
  nor (_29960_, _29959_, _29953_);
  nor (_29961_, _28108_, _16795_);
  not (_29962_, _29961_);
  nor (_29963_, _26928_, _15970_);
  nor (_29964_, _26885_, _16991_);
  nor (_29965_, _29964_, _29963_);
  and (_29966_, _29965_, _29962_);
  and (_29967_, _29966_, _29960_);
  not (_29968_, _29967_);
  nor (_29969_, _29968_, _29952_);
  and (_29970_, _29969_, _29948_);
  not (_29971_, _29970_);
  nor (_29972_, _29971_, _29936_);
  and (_29973_, _29972_, _29933_);
  not (_29974_, _29973_);
  nor (_29975_, _29974_, _29928_);
  and (_29976_, _29975_, _29927_);
  not (_29977_, _29976_);
  or (_29978_, _29977_, _24379_);
  not (_29979_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_29980_, _24379_, _29979_);
  and (_29981_, _29980_, _27202_);
  and (_29982_, _29981_, _29978_);
  nor (_29983_, _27201_, _29979_);
  not (_29984_, _27836_);
  nand (_29985_, _29984_, _27803_);
  and (_29986_, _29985_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_29987_, _27825_, _24056_);
  and (_29988_, _29987_, _28359_);
  nor (_29989_, _27825_, _29979_);
  or (_29990_, _29989_, _29988_);
  and (_29991_, _29990_, _27803_);
  or (_29992_, _29991_, _29986_);
  and (_29993_, _29992_, _27869_);
  or (_29994_, _29993_, _29983_);
  or (_29995_, _29994_, _29982_);
  and (_09039_, _29995_, _36029_);
  and (_29996_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_29997_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_29998_, _29997_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_29999_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_30000_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_30001_, _30000_, _29999_);
  and (_30002_, _29997_, _14692_);
  and (_30003_, _30002_, _30001_);
  not (_30004_, _30003_);
  and (_30005_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30006_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30007_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30008_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_30009_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_30010_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30011_, _30010_, _30009_);
  and (_30012_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_30013_, _30010_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_30014_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_30015_, _30014_, _30012_);
  and (_30016_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30017_, _30016_, _30009_);
  and (_30018_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not (_30019_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30020_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _30019_);
  and (_30021_, _30020_, _30009_);
  and (_30022_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_30023_, _30022_, _30018_);
  nor (_30024_, _30010_, _30009_);
  and (_30025_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_30026_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_30027_, _30026_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30028_, _30027_, _30009_);
  and (_30029_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_30030_, _30029_, _30025_);
  and (_30031_, _30030_, _30023_);
  and (_30032_, _30031_, _30015_);
  nor (_30033_, _30032_, _30008_);
  and (_30034_, _30033_, _30007_);
  nor (_30035_, _30034_, _30006_);
  nor (_30036_, _30035_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30037_, _30036_, _30005_);
  nor (_30038_, _30037_, _30004_);
  and (_30039_, _30001_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_30040_, _30039_, _30004_);
  nor (_30041_, _30040_, _30038_);
  not (_30042_, _30041_);
  and (_30043_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30044_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30045_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30046_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_30047_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_30048_, _30047_, _30046_);
  and (_30049_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_30050_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_30051_, _30050_, _30049_);
  and (_30052_, _30051_, _30048_);
  and (_30053_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_30054_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_30055_, _30054_, _30053_);
  and (_30056_, _30055_, _30052_);
  nor (_30057_, _30056_, _30008_);
  and (_30058_, _30057_, _30007_);
  or (_30059_, _30058_, _30045_);
  and (_30060_, _30059_, _30044_);
  nor (_30061_, _30060_, _30043_);
  nor (_30062_, _30061_, _30004_);
  and (_30063_, _30001_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_30064_, _30063_, _30004_);
  nor (_30065_, _30064_, _30062_);
  and (_30066_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_30067_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_30068_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_30069_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_30070_, _30069_, _30068_);
  and (_30071_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_30072_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_30073_, _30072_, _30071_);
  and (_30074_, _30073_, _30070_);
  and (_30075_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_30076_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_30077_, _30076_, _30075_);
  and (_30078_, _30077_, _30074_);
  nor (_30079_, _30078_, _30008_);
  and (_30080_, _30079_, _30007_);
  or (_30081_, _30080_, _30067_);
  and (_30082_, _30081_, _30044_);
  nor (_30083_, _30082_, _30066_);
  nor (_30084_, _30083_, _30004_);
  and (_30085_, _30001_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_30086_, _30085_, _30004_);
  nor (_30087_, _30086_, _30084_);
  not (_30088_, _30087_);
  and (_30089_, _30088_, _30065_);
  and (_30090_, _30089_, _30042_);
  and (_30091_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30092_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30093_, _30008_);
  and (_30094_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_30095_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_30096_, _30095_, _30094_);
  and (_30097_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_30098_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_30099_, _30098_, _30097_);
  and (_30100_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_30101_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_30102_, _30101_, _30100_);
  and (_30103_, _30102_, _30099_);
  and (_30104_, _30103_, _30096_);
  and (_30105_, _30104_, _30093_);
  nor (_30106_, _30105_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30107_, _30106_, _30092_);
  nor (_30108_, _30107_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30109_, _30108_, _30091_);
  nor (_30110_, _30109_, _30004_);
  and (_30111_, _30001_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_30112_, _30111_, _30004_);
  nor (_30113_, _30112_, _30110_);
  and (_30114_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30115_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30116_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_30117_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_30118_, _30117_, _30116_);
  and (_30119_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_30120_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_30121_, _30120_, _30119_);
  and (_30122_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_30123_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_30124_, _30123_, _30122_);
  and (_30125_, _30124_, _30121_);
  and (_30126_, _30125_, _30118_);
  nor (_30127_, _30126_, _30008_);
  and (_30128_, _30127_, _30007_);
  or (_30129_, _30128_, _30115_);
  and (_30130_, _30129_, _30044_);
  nor (_30131_, _30130_, _30114_);
  nor (_30132_, _30131_, _30004_);
  and (_30133_, _30001_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_30134_, _30133_, _30004_);
  nor (_30135_, _30134_, _30132_);
  nor (_30136_, _30135_, _30113_);
  and (_30137_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30138_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30139_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_30140_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_30141_, _30140_, _30139_);
  and (_30142_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_30143_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_30144_, _30143_, _30142_);
  and (_30145_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_30146_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_30147_, _30146_, _30145_);
  and (_30148_, _30147_, _30144_);
  and (_30149_, _30148_, _30141_);
  nor (_30150_, _30149_, _30008_);
  and (_30151_, _30150_, _30007_);
  nor (_30152_, _30151_, _30138_);
  nor (_30153_, _30152_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30154_, _30153_, _30137_);
  nor (_30155_, _30154_, _30004_);
  and (_30156_, _30001_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_30157_, _30156_, _30004_);
  nor (_30158_, _30157_, _30155_);
  nor (_30159_, _30008_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30160_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_30161_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_30162_, _30161_, _30160_);
  and (_30163_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_30164_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_30165_, _30164_, _30163_);
  and (_30166_, _30165_, _30162_);
  and (_30167_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_30168_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_30169_, _30168_, _30167_);
  and (_30170_, _30169_, _30166_);
  and (_30171_, _30170_, _30159_);
  nor (_30172_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _30007_);
  or (_30173_, _30172_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30174_, _30173_, _30171_);
  and (_30175_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_30176_, _30175_, _30174_);
  and (_30177_, _30176_, _30003_);
  and (_30178_, _30001_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_30179_, _30178_, _30004_);
  nor (_30180_, _30179_, _30177_);
  not (_30181_, _30180_);
  and (_30182_, _30181_, _30158_);
  and (_30183_, _30182_, _30136_);
  and (_30184_, _30183_, _30090_);
  and (_30185_, _30136_, _30158_);
  and (_30186_, _30087_, _30065_);
  and (_30187_, _30186_, _30041_);
  and (_30188_, _30187_, _30185_);
  nor (_30189_, _30188_, _30184_);
  and (_30190_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30191_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30192_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_30193_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_30194_, _30193_, _30192_);
  and (_30195_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_30196_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_30197_, _30196_, _30195_);
  and (_30198_, _30197_, _30194_);
  and (_30199_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_30200_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_30201_, _30200_, _30199_);
  and (_30202_, _30201_, _30198_);
  nor (_30203_, _30202_, _30008_);
  and (_30204_, _30203_, _30007_);
  or (_30205_, _30204_, _30191_);
  and (_30206_, _30205_, _30044_);
  nor (_30207_, _30206_, _30190_);
  nor (_30208_, _30207_, _30004_);
  and (_30209_, _30001_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_30210_, _30209_, _30004_);
  nor (_30211_, _30210_, _30208_);
  not (_30212_, _30113_);
  and (_30213_, _30158_, _30135_);
  and (_30214_, _30213_, _30212_);
  and (_30215_, _30214_, _30211_);
  and (_30216_, _30186_, _30042_);
  and (_30217_, _30216_, _30215_);
  and (_30218_, _30180_, _30185_);
  not (_30219_, _30065_);
  and (_30220_, _30087_, _30219_);
  and (_30221_, _30220_, _30041_);
  nor (_30222_, _30087_, _30065_);
  and (_30223_, _30222_, _30042_);
  or (_30224_, _30223_, _30221_);
  and (_30225_, _30224_, _30218_);
  nor (_30226_, _30225_, _30217_);
  and (_30227_, _30226_, _30189_);
  and (_30228_, _30222_, _30041_);
  and (_30229_, _30228_, _30185_);
  and (_30231_, _30089_, _30041_);
  and (_30232_, _30231_, _30183_);
  nor (_30234_, _30232_, _30229_);
  not (_30235_, _30234_);
  not (_30237_, _30185_);
  and (_30238_, _30221_, _30181_);
  nor (_30240_, _30238_, _30216_);
  nor (_30241_, _30240_, _30237_);
  nor (_30242_, _30241_, _30235_);
  and (_30243_, _30242_, _30227_);
  and (_30244_, _30090_, _30180_);
  not (_30245_, _30211_);
  and (_30246_, _30214_, _30245_);
  and (_30247_, _30246_, _30244_);
  not (_30248_, _30247_);
  nor (_30249_, _30065_, _30041_);
  and (_30250_, _30249_, _30087_);
  and (_30251_, _30250_, _30181_);
  and (_30252_, _30251_, _30246_);
  and (_30253_, _30231_, _30181_);
  and (_30254_, _30246_, _30253_);
  nor (_30255_, _30254_, _30252_);
  and (_30256_, _30255_, _30248_);
  and (_30257_, _30228_, _30181_);
  and (_30258_, _30211_, _30113_);
  and (_30259_, _30258_, _30213_);
  and (_30260_, _30259_, _30257_);
  not (_30261_, _30260_);
  and (_30262_, _30250_, _30180_);
  and (_30263_, _30262_, _30185_);
  and (_30264_, _30041_, _30180_);
  and (_30265_, _30264_, _30089_);
  and (_30266_, _30265_, _30185_);
  nor (_30267_, _30266_, _30263_);
  and (_30268_, _30267_, _30261_);
  and (_30269_, _30268_, _30256_);
  and (_30270_, _30269_, _30243_);
  nor (_30271_, _30270_, _29998_);
  not (_30272_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30273_, _14692_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_30274_, _30273_, _30272_);
  and (_30275_, _30274_, _30259_);
  and (_30276_, _30275_, _30250_);
  and (_30277_, _30217_, _30273_);
  and (_30278_, _30277_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_30279_, _30278_, _30276_);
  nor (_30280_, _30279_, _30271_);
  nor (_30281_, _30280_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30282_, _30281_, _29996_);
  and (_30283_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_30284_, _30135_);
  and (_30285_, _30158_, _30284_);
  and (_30286_, _30245_, _30113_);
  and (_30287_, _30286_, _30285_);
  and (_30288_, _30287_, _30257_);
  and (_30289_, _30251_, _30215_);
  and (_30290_, _30264_, _30220_);
  and (_30291_, _30290_, _30214_);
  nor (_30292_, _30291_, _30289_);
  not (_30293_, _30292_);
  nor (_30294_, _30293_, _30288_);
  and (_30295_, _30090_, _30181_);
  and (_30296_, _30215_, _30295_);
  and (_30297_, _30228_, _30180_);
  and (_30298_, _30297_, _30215_);
  nor (_30299_, _30298_, _30296_);
  and (_30300_, _30290_, _30287_);
  and (_30301_, _30259_, _30244_);
  nor (_30302_, _30301_, _30300_);
  and (_30303_, _30187_, _30181_);
  and (_30304_, _30303_, _30287_);
  and (_30305_, _30259_, _30295_);
  nor (_30306_, _30305_, _30304_);
  and (_30307_, _30306_, _30302_);
  and (_30308_, _30307_, _30299_);
  and (_30309_, _30308_, _30294_);
  and (_30310_, _30259_, _30228_);
  and (_30311_, _30262_, _30214_);
  nor (_30312_, _30311_, _30310_);
  and (_30313_, _30253_, _30215_);
  and (_30314_, _30287_, _30265_);
  nor (_30315_, _30314_, _30313_);
  and (_30316_, _30315_, _30312_);
  and (_30317_, _30265_, _30215_);
  and (_30318_, _30238_, _30214_);
  nor (_30319_, _30318_, _30317_);
  not (_30320_, _30319_);
  and (_30321_, _30089_, _30181_);
  and (_30322_, _30321_, _30287_);
  nor (_30323_, _30322_, _30320_);
  and (_30324_, _30323_, _30316_);
  not (_30325_, _30287_);
  nor (_30326_, _30325_, _30240_);
  and (_30327_, _30223_, _30180_);
  and (_30328_, _30327_, _30287_);
  nor (_30329_, _30328_, _30217_);
  not (_30330_, _30329_);
  nor (_30331_, _30330_, _30326_);
  and (_30332_, _30257_, _30215_);
  and (_30333_, _30244_, _30215_);
  nor (_30334_, _30333_, _30332_);
  and (_30335_, _30287_, _30262_);
  and (_30336_, _30297_, _30287_);
  nor (_30337_, _30336_, _30335_);
  and (_30338_, _30337_, _30334_);
  and (_30339_, _30338_, _30331_);
  and (_30340_, _30259_, _30216_);
  and (_30341_, _30340_, _30180_);
  not (_30342_, _30259_);
  and (_30343_, _30216_, _30181_);
  nor (_30344_, _30303_, _30343_);
  nor (_30345_, _30344_, _30342_);
  nor (_30346_, _30345_, _30341_);
  and (_30347_, _30264_, _30186_);
  and (_30348_, _30347_, _30287_);
  not (_30349_, _30348_);
  and (_30350_, _30218_, _30090_);
  not (_30351_, _30158_);
  and (_30352_, _30244_, _30351_);
  nor (_30353_, _30352_, _30350_);
  and (_30354_, _30353_, _30349_);
  and (_30355_, _30354_, _30346_);
  and (_30356_, _30355_, _30339_);
  and (_30357_, _30356_, _30324_);
  and (_30358_, _30357_, _30309_);
  nor (_30359_, _30358_, _29998_);
  and (_30360_, _30273_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30361_, _30360_, _30217_);
  not (_30362_, _30361_);
  and (_30363_, _30259_, _30220_);
  and (_30364_, _30363_, _30274_);
  not (_30365_, _30274_);
  nor (_30366_, _30041_, _30181_);
  and (_30367_, _30366_, _30186_);
  and (_30368_, _30259_, _30367_);
  and (_30369_, _30303_, _30259_);
  nor (_30370_, _30369_, _30368_);
  nor (_30371_, _30370_, _30365_);
  nor (_30372_, _30371_, _30364_);
  and (_30373_, _30372_, _30362_);
  not (_30374_, _30373_);
  nor (_30375_, _30374_, _30359_);
  nor (_30376_, _30375_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30377_, _30376_, _30283_);
  nor (_30378_, _30377_, _30282_);
  and (_30379_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30380_, _30258_, _30285_);
  and (_30381_, _30380_, _30265_);
  and (_30382_, _30380_, _30244_);
  nor (_30383_, _30382_, _30381_);
  and (_30384_, _30383_, _30256_);
  nor (_30385_, _30384_, _29998_);
  not (_30386_, _30385_);
  and (_30387_, _30382_, _14692_);
  and (_30388_, _30381_, _14692_);
  nor (_30389_, _30388_, _30387_);
  nor (_30390_, _30389_, _29997_);
  nor (_30391_, _30390_, _30364_);
  and (_30392_, _30391_, _30386_);
  nor (_30393_, _30392_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30394_, _30393_, _30379_);
  and (_30395_, _30394_, _36029_);
  and (_09590_, _30395_, _30378_);
  and (_30396_, _27202_, _23606_);
  and (_30397_, _23924_, _23287_);
  nor (_30398_, _23781_, _23420_);
  and (_30399_, _30398_, _30397_);
  and (_30400_, _30399_, _29027_);
  and (_30401_, _30400_, _30396_);
  nor (_30402_, _20094_, _14758_);
  and (_30403_, _26128_, _20072_);
  nor (_30404_, _26917_, _30403_);
  and (_30405_, _30404_, _26885_);
  and (_30406_, _30405_, _30402_);
  and (_30407_, _30406_, _28108_);
  nor (_30408_, _30407_, _16795_);
  not (_30409_, _30408_);
  and (_30410_, _30409_, _26863_);
  and (_30411_, _30410_, _26808_);
  and (_30412_, _30411_, _26513_);
  not (_30413_, _30412_);
  and (_30414_, _30413_, _30401_);
  and (_30415_, _23770_, _23606_);
  and (_30416_, _30415_, _27781_);
  and (_30417_, _30416_, _30397_);
  and (_30418_, _30417_, _29027_);
  and (_30419_, _30418_, _27202_);
  not (_30420_, _30419_);
  and (_30421_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_30422_, _30407_, _15970_);
  not (_30423_, _30422_);
  and (_30424_, _30423_, _29960_);
  and (_30425_, _30424_, _29948_);
  nor (_30426_, _30425_, _30420_);
  nor (_30427_, _30426_, _30421_);
  and (_30428_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_30429_, _30407_, _16991_);
  not (_30430_, _30429_);
  and (_30431_, _30430_, _29888_);
  and (_30432_, _30431_, _29875_);
  nor (_30433_, _30432_, _30420_);
  nor (_30434_, _30433_, _30428_);
  and (_30435_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_30436_, _30407_, _17166_);
  nor (_30437_, _30436_, _29817_);
  and (_30438_, _30437_, _29811_);
  and (_30439_, _30438_, _29808_);
  nor (_30440_, _30439_, _30420_);
  nor (_30441_, _30440_, _30435_);
  and (_30442_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_30443_, _30407_, _17504_);
  not (_30444_, _30443_);
  and (_30445_, _30444_, _29748_);
  and (_30446_, _30445_, _29724_);
  and (_30447_, _30446_, _29737_);
  nor (_30448_, _30447_, _30420_);
  nor (_30449_, _30448_, _30442_);
  and (_30450_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_30451_, _30407_, _18028_);
  not (_30452_, _30451_);
  and (_30453_, _30452_, _29323_);
  and (_30454_, _30453_, _29356_);
  and (_30455_, _30454_, _29246_);
  nor (_30456_, _30455_, _30420_);
  nor (_30457_, _30456_, _30450_);
  and (_30458_, _30420_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_30459_, _30407_, _17853_);
  not (_30460_, _30459_);
  and (_30461_, _30460_, _28703_);
  and (_30462_, _30461_, _28886_);
  nor (_30463_, _30462_, _30420_);
  nor (_30464_, _30463_, _30458_);
  nor (_30465_, _30401_, _24001_);
  nor (_30466_, _30407_, _18398_);
  not (_30467_, _30466_);
  and (_30468_, _30467_, _28206_);
  and (_30469_, _30468_, _28173_);
  and (_30470_, _30469_, _28086_);
  not (_30471_, _30470_);
  and (_30472_, _30471_, _30401_);
  nor (_30473_, _30472_, _30465_);
  and (_30474_, _30473_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30475_, _30474_, _30464_);
  and (_30476_, _30475_, _30457_);
  and (_30477_, _30476_, _30449_);
  and (_30478_, _30477_, _30441_);
  and (_30479_, _30478_, _30434_);
  and (_30480_, _30479_, _30427_);
  nor (_30481_, _30401_, _23288_);
  and (_30482_, _30481_, _30480_);
  nor (_30483_, _30481_, _30480_);
  nor (_30484_, _30483_, _30482_);
  and (_30485_, _30484_, _23058_);
  nor (_30486_, _30485_, _23332_);
  nor (_30487_, _30486_, _30419_);
  nor (_30488_, _30487_, _30414_);
  nor (_09611_, _30488_, rst);
  not (_30489_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30490_, _30473_, _30489_);
  nor (_30491_, _30473_, _30489_);
  nor (_30492_, _30491_, _30490_);
  and (_30493_, _30492_, _23058_);
  nor (_30494_, _30493_, _24012_);
  nor (_30495_, _30494_, _30419_);
  nor (_30496_, _30495_, _30472_);
  nand (_10725_, _30496_, _36029_);
  nor (_30497_, _30474_, _30464_);
  nor (_30498_, _30497_, _30475_);
  nor (_30499_, _30498_, _23047_);
  nor (_30500_, _30499_, _24088_);
  nor (_30501_, _30500_, _30419_);
  nor (_30502_, _30501_, _30463_);
  nand (_10736_, _30502_, _36029_);
  nor (_30503_, _30475_, _30457_);
  nor (_30504_, _30503_, _30476_);
  nor (_30505_, _30504_, _23047_);
  nor (_30506_, _30505_, _24220_);
  nor (_30507_, _30506_, _30419_);
  nor (_30508_, _30507_, _30456_);
  nand (_10747_, _30508_, _36029_);
  nor (_30509_, _30476_, _30449_);
  nor (_30510_, _30509_, _30477_);
  nor (_30511_, _30510_, _23047_);
  nor (_30512_, _30511_, _23507_);
  nor (_30513_, _30512_, _30419_);
  nor (_30514_, _30513_, _30448_);
  nor (_10758_, _30514_, rst);
  nor (_30515_, _30477_, _30441_);
  nor (_30516_, _30515_, _30478_);
  nor (_30517_, _30516_, _23047_);
  nor (_30518_, _30517_, _23650_);
  nor (_30519_, _30518_, _30419_);
  nor (_30520_, _30519_, _30440_);
  nor (_10769_, _30520_, rst);
  nor (_30521_, _30478_, _30434_);
  nor (_30522_, _30521_, _30479_);
  nor (_30523_, _30522_, _23047_);
  nor (_30524_, _30523_, _23836_);
  nor (_30525_, _30524_, _30419_);
  nor (_30526_, _30525_, _30433_);
  nor (_10780_, _30526_, rst);
  nor (_30527_, _30479_, _30427_);
  nor (_30528_, _30527_, _30480_);
  nor (_30529_, _30528_, _23047_);
  nor (_30530_, _30529_, _23091_);
  nor (_30531_, _30530_, _30419_);
  nor (_30532_, _30531_, _30426_);
  nor (_10791_, _30532_, rst);
  and (_30533_, _30396_, _29769_);
  nand (_30534_, _30533_, _30399_);
  nor (_30535_, _30534_, _27126_);
  and (_30536_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _14692_);
  and (_30537_, _30536_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_30538_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_30539_, _30538_, _30537_);
  or (_30540_, _30539_, _30535_);
  nor (_30541_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_30542_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_30543_, _30542_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30544_, _30543_, _30541_);
  nor (_30545_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_30546_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_30547_, _30546_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30548_, _30547_, _30545_);
  nor (_30549_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_30550_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_30551_, _30550_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30552_, _30551_, _30549_);
  not (_30553_, _30552_);
  nor (_30554_, _30553_, _27267_);
  nor (_30555_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_30556_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_30557_, _30556_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30558_, _30557_, _30555_);
  and (_30559_, _30558_, _30554_);
  nor (_30560_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_30561_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_30562_, _30561_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30563_, _30562_, _30560_);
  and (_30564_, _30563_, _30559_);
  and (_30565_, _30564_, _30548_);
  nor (_30566_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_30567_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_30568_, _30567_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30569_, _30568_, _30566_);
  and (_30570_, _30569_, _30565_);
  and (_30571_, _30570_, _30544_);
  nor (_30572_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_30573_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_30574_, _30573_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30575_, _30574_, _30572_);
  and (_30576_, _30575_, _30571_);
  nor (_30577_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_30578_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_30579_, _30578_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30580_, _30579_, _30577_);
  nor (_30581_, _30580_, _30576_);
  and (_30582_, _30580_, _30576_);
  or (_30583_, _30582_, _30581_);
  nor (_30584_, _30583_, _26150_);
  not (_30585_, _30584_);
  and (_30586_, _19785_, _14758_);
  and (_30587_, _25512_, _16296_);
  not (_30588_, _30587_);
  nor (_30589_, _16795_, _15480_);
  and (_30590_, _30589_, _26260_);
  and (_30591_, _30590_, _24908_);
  and (_30592_, _30591_, _24952_);
  and (_30593_, _30592_, _25567_);
  nor (_30594_, _30593_, _26282_);
  and (_30595_, _25512_, _15316_);
  nor (_30596_, _30595_, _30594_);
  and (_30597_, _30596_, _30588_);
  and (_30598_, _26348_, _16795_);
  and (_30599_, _16144_, _15151_);
  and (_30600_, _16459_, _15480_);
  and (_30601_, _30600_, _30599_);
  and (_30602_, _30601_, _30598_);
  and (_30603_, _16296_, _15316_);
  and (_30604_, _30603_, _30602_);
  nor (_30605_, _30604_, _25512_);
  not (_30606_, _30605_);
  and (_30607_, _30606_, _30597_);
  nor (_30608_, _25512_, _15654_);
  and (_30609_, _25512_, _15654_);
  nor (_30610_, _30609_, _30608_);
  and (_30611_, _30610_, _30607_);
  and (_30612_, _30611_, _26425_);
  nor (_30613_, _30611_, _26425_);
  nor (_30614_, _30613_, _30612_);
  and (_30615_, _30614_, _26194_);
  and (_30616_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_30617_, _25512_, _26425_);
  nor (_30618_, _30617_, _27388_);
  nor (_30619_, _30618_, _26480_);
  nor (_30620_, _27563_, _17504_);
  nor (_30621_, _26928_, _16634_);
  or (_30622_, _30621_, _30620_);
  or (_30623_, _30622_, _30619_);
  nor (_30624_, _30623_, _30616_);
  not (_30625_, _30624_);
  nor (_30626_, _30625_, _30615_);
  not (_30627_, _30626_);
  nor (_30628_, _30627_, _30586_);
  and (_30629_, _30628_, _30585_);
  nand (_30630_, _30629_, _30537_);
  and (_30631_, _30630_, _36029_);
  and (_12626_, _30631_, _30540_);
  and (_30632_, _30396_, _29706_);
  and (_30633_, _30632_, _30399_);
  nor (_30634_, _30633_, _30537_);
  not (_30635_, _30634_);
  nand (_30636_, _30635_, _27126_);
  not (_30637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_30638_, _30634_, _30637_);
  and (_30639_, _30638_, _36029_);
  and (_12646_, _30639_, _30636_);
  nor (_30640_, _30534_, _28302_);
  and (_30641_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_30642_, _30641_, _30537_);
  or (_30643_, _30642_, _30640_);
  and (_30644_, _22401_, _20094_);
  not (_30645_, _30644_);
  and (_30646_, _30553_, _27267_);
  nor (_30647_, _30646_, _30554_);
  and (_30648_, _30647_, _26139_);
  nor (_30649_, _27388_, _26458_);
  not (_30650_, _30649_);
  nor (_30651_, _30650_, _26370_);
  nor (_30652_, _30651_, _24875_);
  and (_30653_, _30651_, _24875_);
  nor (_30654_, _30653_, _30652_);
  and (_30655_, _30654_, _26194_);
  nor (_30656_, _26928_, _15480_);
  and (_30657_, _19563_, _14758_);
  nor (_30658_, _27563_, _17166_);
  nor (_30659_, _26480_, _18398_);
  or (_30660_, _30659_, _30658_);
  or (_30661_, _30660_, _30657_);
  nor (_30662_, _30661_, _30656_);
  not (_30663_, _30662_);
  nor (_30664_, _30663_, _30655_);
  not (_30665_, _30664_);
  nor (_30666_, _30665_, _30648_);
  and (_30667_, _30666_, _30645_);
  nand (_30668_, _30667_, _30537_);
  and (_30669_, _30668_, _36029_);
  and (_13561_, _30669_, _30643_);
  nor (_30670_, _30534_, _28939_);
  and (_30671_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_30672_, _30671_, _30537_);
  or (_30673_, _30672_, _30670_);
  nor (_30674_, _30558_, _30554_);
  nor (_30675_, _30674_, _30559_);
  and (_30676_, _30675_, _26139_);
  not (_30677_, _30676_);
  and (_30678_, _21386_, _20094_);
  and (_30679_, _30590_, _25512_);
  and (_30680_, _30598_, _15480_);
  and (_30681_, _30680_, _26282_);
  nor (_30682_, _30681_, _30679_);
  and (_30683_, _30682_, _16459_);
  nor (_30684_, _30682_, _16459_);
  or (_30685_, _30684_, _29733_);
  nor (_30686_, _30685_, _30683_);
  nor (_30687_, _26928_, _16459_);
  and (_30688_, _19595_, _14758_);
  nor (_30689_, _27563_, _16991_);
  nor (_30690_, _26480_, _17853_);
  or (_30691_, _30690_, _30689_);
  or (_30692_, _30691_, _30688_);
  nor (_30693_, _30692_, _30687_);
  not (_30694_, _30693_);
  nor (_30695_, _30694_, _30686_);
  not (_30696_, _30695_);
  nor (_30697_, _30696_, _30678_);
  and (_30698_, _30697_, _30677_);
  nand (_30699_, _30698_, _30537_);
  and (_30700_, _30699_, _36029_);
  and (_13572_, _30700_, _30673_);
  nor (_30701_, _30534_, _29584_);
  and (_30702_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_30703_, _30702_, _30537_);
  or (_30704_, _30703_, _30701_);
  nor (_30705_, _30563_, _30559_);
  nor (_30706_, _30705_, _30564_);
  and (_30707_, _30706_, _26139_);
  not (_30708_, _30707_);
  and (_30709_, _30680_, _16459_);
  and (_30710_, _30709_, _26282_);
  and (_30711_, _30591_, _25512_);
  nor (_30712_, _30711_, _30710_);
  and (_30713_, _30712_, _15151_);
  nor (_30714_, _30712_, _15151_);
  nor (_30715_, _30714_, _30713_);
  and (_30716_, _30715_, _26194_);
  not (_30717_, _30716_);
  nor (_30718_, _26480_, _18028_);
  and (_30719_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_30720_, _30719_, _30718_);
  and (_30721_, _19626_, _14758_);
  nor (_30722_, _27563_, _15970_);
  nor (_30723_, _26928_, _15151_);
  or (_30724_, _30723_, _30722_);
  nor (_30725_, _30724_, _30721_);
  and (_30726_, _30725_, _30720_);
  and (_30727_, _30726_, _30717_);
  and (_30728_, _30727_, _30708_);
  nand (_30729_, _30728_, _30537_);
  and (_30730_, _30729_, _36029_);
  and (_13582_, _30730_, _30704_);
  nor (_30731_, _30534_, _29760_);
  and (_30732_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_30733_, _30732_, _30537_);
  or (_30734_, _30733_, _30731_);
  nor (_30735_, _30564_, _30548_);
  nor (_30736_, _30735_, _30565_);
  and (_30737_, _30736_, _26139_);
  not (_30738_, _30737_);
  nor (_30739_, _30592_, _25567_);
  not (_30740_, _30739_);
  and (_30741_, _30740_, _30594_);
  and (_30742_, _30709_, _15151_);
  nor (_30743_, _30742_, _16144_);
  nor (_30744_, _30743_, _30602_);
  nor (_30745_, _30744_, _25512_);
  nor (_30746_, _30745_, _30741_);
  nor (_30747_, _30746_, _29733_);
  nor (_30748_, _26928_, _16144_);
  or (_30749_, _30748_, _27574_);
  nor (_30750_, _30749_, _30747_);
  and (_30751_, _19658_, _14758_);
  nor (_30752_, _26480_, _17504_);
  and (_30753_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_30754_, _30753_, _30752_);
  nor (_30755_, _30754_, _30751_);
  and (_30756_, _30755_, _30750_);
  and (_30757_, _30756_, _30738_);
  nand (_30758_, _30757_, _30537_);
  and (_30759_, _30758_, _36029_);
  and (_13593_, _30759_, _30734_);
  nor (_30760_, _30534_, _29830_);
  and (_30761_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_30762_, _30761_, _30537_);
  or (_30763_, _30762_, _30760_);
  nor (_30764_, _30569_, _30565_);
  not (_30765_, _30764_);
  nor (_30766_, _30570_, _26150_);
  and (_30767_, _30766_, _30765_);
  not (_30769_, _30767_);
  and (_30772_, _19690_, _14758_);
  nor (_30773_, _30602_, _25512_);
  nor (_30774_, _30773_, _30594_);
  nor (_30775_, _30774_, _24600_);
  and (_30776_, _30774_, _24600_);
  nor (_30777_, _30776_, _30775_);
  and (_30778_, _30777_, _26194_);
  nor (_30779_, _25512_, _17177_);
  not (_30780_, _30779_);
  nor (_30781_, _30595_, _26480_);
  and (_30782_, _30781_, _30780_);
  and (_30790_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_30796_, _27563_, _18398_);
  nor (_30802_, _26928_, _15316_);
  or (_30807_, _30802_, _30796_);
  nor (_30808_, _30807_, _30790_);
  not (_30809_, _30808_);
  nor (_30810_, _30809_, _30782_);
  not (_30811_, _30810_);
  nor (_30812_, _30811_, _30778_);
  not (_30813_, _30812_);
  nor (_30814_, _30813_, _30772_);
  and (_30815_, _30814_, _30769_);
  nand (_30816_, _30815_, _30537_);
  and (_30817_, _30816_, _36029_);
  and (_13604_, _30817_, _30763_);
  nor (_30818_, _30534_, _29903_);
  and (_30819_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_30820_, _30819_, _30537_);
  or (_30821_, _30820_, _30818_);
  nor (_30822_, _30570_, _30544_);
  nor (_30823_, _30822_, _30571_);
  and (_30824_, _30823_, _26139_);
  not (_30825_, _30824_);
  and (_30826_, _19721_, _14758_);
  and (_30827_, _30602_, _15316_);
  nor (_30828_, _30827_, _25512_);
  not (_30829_, _30828_);
  and (_30830_, _30829_, _30596_);
  and (_30831_, _30830_, _16296_);
  nor (_30834_, _30830_, _16296_);
  or (_30835_, _30834_, _30831_);
  and (_30836_, _30835_, _26194_);
  nor (_30837_, _29940_, _26480_);
  and (_30838_, _30837_, _30588_);
  nor (_30839_, _26928_, _16296_);
  nor (_30840_, _27563_, _17853_);
  and (_30841_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_30842_, _30841_, _30840_);
  nor (_30843_, _30842_, _30839_);
  not (_30844_, _30843_);
  nor (_30845_, _30844_, _30838_);
  not (_30846_, _30845_);
  nor (_30847_, _30846_, _30836_);
  not (_30848_, _30847_);
  nor (_30849_, _30848_, _30826_);
  and (_30850_, _30849_, _30825_);
  nand (_30851_, _30850_, _30537_);
  and (_30852_, _30851_, _36029_);
  and (_13615_, _30852_, _30821_);
  nor (_30853_, _30534_, _29976_);
  and (_30854_, _30534_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_30855_, _30854_, _30537_);
  or (_30856_, _30855_, _30853_);
  nor (_30857_, _30575_, _30571_);
  nor (_30858_, _30857_, _30576_);
  and (_30859_, _30858_, _26139_);
  not (_30860_, _30859_);
  and (_30861_, _19753_, _14758_);
  nor (_30862_, _30607_, _15654_);
  and (_30863_, _30607_, _15654_);
  nor (_30864_, _30863_, _30862_);
  nor (_30865_, _30864_, _29733_);
  nor (_30866_, _25512_, _15981_);
  not (_30867_, _30866_);
  nor (_30868_, _30609_, _26480_);
  and (_30869_, _30868_, _30867_);
  and (_30870_, _20094_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_30872_, _27563_, _18028_);
  nor (_30876_, _26928_, _15654_);
  or (_30882_, _30876_, _30872_);
  nor (_30887_, _30882_, _30870_);
  not (_30894_, _30887_);
  nor (_30902_, _30894_, _30869_);
  not (_30910_, _30902_);
  nor (_30911_, _30910_, _30865_);
  not (_30912_, _30911_);
  nor (_30913_, _30912_, _30861_);
  and (_30914_, _30913_, _30860_);
  nand (_30915_, _30914_, _30537_);
  and (_30916_, _30915_, _36029_);
  and (_13626_, _30916_, _30856_);
  nand (_30917_, _30635_, _28302_);
  not (_30918_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_30919_, _30634_, _30918_);
  and (_30920_, _30919_, _36029_);
  and (_13637_, _30920_, _30917_);
  nand (_30921_, _30635_, _28939_);
  not (_30922_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_30923_, _30634_, _30922_);
  and (_30924_, _30923_, _36029_);
  and (_13648_, _30924_, _30921_);
  nand (_30925_, _30635_, _29584_);
  not (_30926_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_30927_, _30634_, _30926_);
  and (_30928_, _30927_, _36029_);
  and (_13659_, _30928_, _30925_);
  nand (_30929_, _30635_, _29760_);
  or (_30930_, _30635_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_30931_, _30930_, _36029_);
  and (_13670_, _30931_, _30929_);
  nand (_30932_, _30635_, _29830_);
  or (_30933_, _30635_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_30934_, _30933_, _36029_);
  and (_13681_, _30934_, _30932_);
  nand (_30935_, _30635_, _29903_);
  or (_30936_, _30635_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_30937_, _30936_, _36029_);
  and (_13692_, _30937_, _30935_);
  nand (_30938_, _30635_, _29976_);
  or (_30939_, _30635_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_30940_, _30939_, _36029_);
  and (_13703_, _30940_, _30938_);
  and (_30955_, _23792_, _23924_);
  and (_30957_, _30955_, _23431_);
  and (_30958_, _30957_, _27869_);
  nor (_30959_, _29984_, _27760_);
  not (_30969_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_30976_, _27836_, _30969_);
  or (_30977_, _30976_, _30959_);
  and (_30978_, _30977_, _30958_);
  nor (_30979_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_30980_, _30979_);
  nand (_30981_, _30980_, _27760_);
  and (_30982_, _30979_, _30969_);
  not (_30983_, _23287_);
  and (_30984_, _30955_, _30983_);
  and (_30985_, _27869_, _27781_);
  and (_30986_, _30985_, _30984_);
  nor (_30987_, _30986_, _30982_);
  and (_30988_, _30987_, _30981_);
  and (_30989_, _27202_, _24343_);
  and (_30990_, _30989_, _30957_);
  or (_30991_, _30990_, _30988_);
  or (_30992_, _30991_, _30978_);
  nand (_30993_, _30990_, _30412_);
  and (_30994_, _30993_, _30992_);
  and (_16677_, _30994_, _36029_);
  not (_30995_, _30990_);
  not (_30996_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_30997_, _30958_, _29027_);
  nand (_30998_, _30997_, _30996_);
  and (_30999_, _30998_, _30995_);
  or (_31000_, _30997_, _28359_);
  and (_31001_, _31000_, _30999_);
  nor (_31002_, _30995_, _30462_);
  or (_31003_, _31002_, _31001_);
  and (_21606_, _31003_, _36029_);
  not (_31004_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_31005_, _29706_, _31004_);
  or (_31006_, _31005_, _29707_);
  and (_31007_, _31006_, _30958_);
  or (_31008_, _19848_, _19817_);
  or (_31009_, _31008_, _19880_);
  or (_31010_, _31009_, _19923_);
  or (_31011_, _31010_, _19954_);
  or (_31012_, _31011_, _19997_);
  or (_31013_, _31012_, _20029_);
  or (_31014_, _31013_, _19500_);
  and (_31015_, _31014_, _14758_);
  or (_31016_, _27311_, _25666_);
  not (_31017_, _27300_);
  nand (_31018_, _31017_, _25666_);
  and (_31019_, _31018_, _24435_);
  and (_31020_, _31019_, _31016_);
  not (_31021_, _24457_);
  nand (_31022_, _26084_, _31021_);
  or (_31023_, _26084_, _24468_);
  and (_31024_, _26139_, _31023_);
  and (_31025_, _31024_, _31022_);
  and (_31026_, _30603_, _21288_);
  and (_31027_, _30601_, _20094_);
  nand (_31028_, _31027_, _31026_);
  nand (_31029_, _31028_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_31030_, _31029_, _31025_);
  or (_31031_, _31030_, _31020_);
  or (_31032_, _31031_, _31015_);
  nor (_31033_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_31034_, _31033_, _30958_);
  and (_31035_, _31034_, _31032_);
  or (_31036_, _31035_, _31007_);
  and (_31037_, _31036_, _30995_);
  nor (_31038_, _30995_, _30455_);
  or (_31039_, _31038_, _31037_);
  and (_21618_, _31039_, _36029_);
  not (_31040_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_31041_, _30958_, _29769_);
  nand (_31042_, _31041_, _31040_);
  and (_31043_, _31042_, _30995_);
  or (_31044_, _31041_, _28359_);
  and (_31045_, _31044_, _31043_);
  nor (_31046_, _30995_, _30447_);
  or (_31047_, _31046_, _31045_);
  and (_21630_, _31047_, _36029_);
  and (_31048_, _29841_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_31049_, _31048_, _29845_);
  and (_31050_, _31049_, _30958_);
  nor (_31051_, _30995_, _30439_);
  not (_31052_, _30958_);
  or (_31053_, _31052_, _29842_);
  not (_31054_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_31055_, _30990_, _31054_);
  and (_31056_, _31055_, _31053_);
  or (_31057_, _31056_, _31051_);
  or (_31058_, _31057_, _31050_);
  and (_21642_, _31058_, _36029_);
  not (_31059_, _30986_);
  or (_31060_, _31059_, _29912_);
  and (_31061_, _31060_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31062_, _31061_, _30990_);
  and (_31063_, _29918_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31064_, _31063_, _29917_);
  and (_31065_, _31064_, _30958_);
  or (_31066_, _31065_, _31062_);
  nand (_31067_, _30990_, _30432_);
  and (_31068_, _31067_, _31066_);
  and (_21654_, _31068_, _36029_);
  and (_31069_, _25622_, _24435_);
  and (_31070_, _26139_, _25985_);
  and (_31071_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_31072_, _26917_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_31073_, _31072_, _31071_);
  or (_31074_, _31073_, _31070_);
  or (_31075_, _31074_, _31069_);
  or (_31076_, _31071_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_31077_, _31076_, _31075_);
  or (_31078_, _31077_, _30986_);
  nor (_31079_, _29987_, _29741_);
  or (_31080_, _31079_, _29988_);
  or (_31081_, _31080_, _31059_);
  and (_31082_, _31081_, _31078_);
  and (_31083_, _31082_, _30995_);
  nor (_31084_, _30995_, _30425_);
  or (_31085_, _31084_, _31083_);
  and (_21666_, _31085_, _36029_);
  not (_31086_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_31087_, _30536_, _31086_);
  and (_31088_, _31087_, _30629_);
  not (_31089_, _30536_);
  and (_31090_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _14692_);
  and (_31091_, _31090_, _31089_);
  not (_31092_, _31091_);
  not (_31093_, _27202_);
  and (_31094_, _24319_, _23606_);
  nand (_31095_, _31094_, _29839_);
  and (_31096_, _23770_, _23935_);
  nand (_31097_, _31096_, _23431_);
  or (_31098_, _31097_, _31095_);
  or (_31099_, _31098_, _31093_);
  and (_31100_, _31099_, _31092_);
  nor (_31101_, _31100_, _27126_);
  not (_31102_, _31087_);
  and (_31103_, _30415_, _27771_);
  and (_31104_, _31103_, _30985_);
  and (_31105_, _31104_, _27836_);
  and (_31106_, _31105_, _27760_);
  not (_31107_, _31100_);
  nor (_31108_, _31105_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_31109_, _31108_, _31107_);
  or (_31110_, _31109_, _31106_);
  and (_31111_, _31110_, _31102_);
  not (_31112_, _31111_);
  nor (_31113_, _31112_, _31101_);
  nor (_31114_, _31113_, _31088_);
  and (_22441_, _31114_, _36029_);
  and (_31115_, _31087_, _30667_);
  nor (_31116_, _31100_, _28302_);
  and (_31117_, _31104_, _24343_);
  and (_31118_, _31117_, _27760_);
  nor (_31119_, _31117_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_31120_, _31119_, _31107_);
  or (_31121_, _31120_, _31118_);
  and (_31122_, _31121_, _31102_);
  not (_31123_, _31122_);
  nor (_31124_, _31123_, _31116_);
  nor (_31125_, _31124_, _31115_);
  and (_24308_, _31125_, _36029_);
  and (_31126_, _31087_, _30698_);
  nor (_31127_, _31100_, _28939_);
  and (_31128_, _31104_, _29027_);
  and (_31129_, _31128_, _27760_);
  nor (_31130_, _31128_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_31131_, _31130_, _31107_);
  or (_31132_, _31131_, _31129_);
  and (_31133_, _31132_, _31102_);
  not (_31134_, _31133_);
  nor (_31135_, _31134_, _31127_);
  nor (_31136_, _31135_, _31126_);
  and (_24320_, _31136_, _36029_);
  nor (_31137_, _31102_, _30728_);
  and (_31138_, _31107_, _29584_);
  not (_31139_, _31104_);
  not (_31140_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_31141_, _29706_, _31140_);
  nor (_31142_, _31141_, _29707_);
  nor (_31143_, _31142_, _31139_);
  nor (_31144_, _31104_, _31140_);
  nor (_31145_, _31144_, _31107_);
  not (_31146_, _31145_);
  nor (_31147_, _31146_, _31143_);
  nor (_31148_, _31147_, _31087_);
  not (_31149_, _31148_);
  nor (_31150_, _31149_, _31138_);
  nor (_31151_, _31150_, _31137_);
  nor (_24332_, _31151_, rst);
  nor (_31152_, _31102_, _30757_);
  and (_31160_, _31107_, _29760_);
  not (_31171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_31182_, _29769_, _31171_);
  nor (_31192_, _31182_, _29770_);
  nor (_31198_, _31192_, _31139_);
  nor (_31208_, _31104_, _31171_);
  nor (_31219_, _31208_, _31107_);
  not (_31230_, _31219_);
  nor (_31241_, _31230_, _31198_);
  nor (_31252_, _31241_, _31087_);
  not (_31263_, _31252_);
  nor (_31274_, _31263_, _31160_);
  nor (_31285_, _31274_, _31152_);
  nor (_24344_, _31285_, rst);
  and (_31306_, _31087_, _30815_);
  nor (_31317_, _31100_, _29830_);
  and (_31328_, _31104_, _29840_);
  and (_31339_, _31328_, _27760_);
  nor (_31350_, _31328_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_31361_, _31350_, _31107_);
  or (_31366_, _31361_, _31339_);
  and (_31367_, _31366_, _31102_);
  not (_31368_, _31367_);
  nor (_31369_, _31368_, _31317_);
  nor (_31370_, _31369_, _31306_);
  and (_24356_, _31370_, _36029_);
  and (_31371_, _31087_, _30850_);
  nor (_31372_, _31100_, _29903_);
  and (_31373_, _31104_, _29916_);
  and (_31374_, _31373_, _27760_);
  nor (_31375_, _31373_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_31376_, _31375_, _31107_);
  or (_31377_, _31376_, _31374_);
  and (_31378_, _31377_, _31102_);
  not (_31379_, _31378_);
  nor (_31380_, _31379_, _31372_);
  nor (_31381_, _31380_, _31371_);
  and (_24368_, _31381_, _36029_);
  and (_31382_, _31087_, _30914_);
  nor (_31383_, _31100_, _29976_);
  and (_31384_, _31104_, _29987_);
  and (_31385_, _31384_, _27760_);
  nor (_31386_, _31384_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_31387_, _31386_, _31107_);
  or (_31388_, _31387_, _31385_);
  and (_31389_, _31388_, _31102_);
  not (_31390_, _31389_);
  nor (_31391_, _31390_, _31383_);
  nor (_31392_, _31391_, _31382_);
  and (_24380_, _31392_, _36029_);
  and (_31393_, _30417_, _27836_);
  nand (_31394_, _31393_, _27760_);
  or (_31395_, _31393_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31396_, _31395_, _27869_);
  and (_31397_, _31396_, _31394_);
  and (_31398_, _30417_, _24343_);
  nand (_31399_, _31398_, _30412_);
  or (_31400_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31401_, _31400_, _27202_);
  and (_31402_, _31401_, _31399_);
  not (_31403_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_31404_, _27201_, _31403_);
  or (_31405_, _31404_, rst);
  or (_31406_, _31405_, _31402_);
  or (_30230_, _31406_, _31397_);
  nor (_31407_, _23420_, _30983_);
  and (_31408_, _30955_, _31407_);
  and (_31409_, _31408_, _27836_);
  nand (_31410_, _31409_, _27760_);
  or (_31411_, _31409_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_31412_, _31411_, _27869_);
  and (_31413_, _31412_, _31410_);
  and (_31414_, _31408_, _24343_);
  not (_31415_, _31414_);
  nor (_31416_, _31415_, _30412_);
  not (_31417_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_31418_, _31414_, _31417_);
  or (_31419_, _31418_, _31416_);
  and (_31420_, _31419_, _27202_);
  nor (_31421_, _27201_, _31417_);
  or (_31422_, _31421_, rst);
  or (_31423_, _31422_, _31420_);
  or (_30233_, _31423_, _31413_);
  and (_31424_, _23935_, _23287_);
  and (_31425_, _31424_, _30416_);
  and (_31426_, _31425_, _27836_);
  nand (_31427_, _31426_, _27760_);
  or (_31428_, _31426_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_31429_, _31428_, _27869_);
  and (_31430_, _31429_, _31427_);
  and (_31431_, _30415_, _24355_);
  and (_31432_, _31431_, _31407_);
  not (_31433_, _31432_);
  nor (_31434_, _31433_, _30412_);
  not (_31435_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_31436_, _31432_, _31435_);
  or (_31437_, _31436_, _31434_);
  and (_31438_, _31437_, _27202_);
  nor (_31439_, _27201_, _31435_);
  or (_31440_, _31439_, rst);
  or (_31441_, _31440_, _31438_);
  or (_30236_, _31441_, _31430_);
  and (_31442_, _31424_, _27792_);
  and (_31443_, _31442_, _27836_);
  nand (_31444_, _31443_, _27760_);
  or (_31445_, _31443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_31446_, _31445_, _27869_);
  and (_31447_, _31446_, _31444_);
  and (_31448_, _31407_, _24367_);
  not (_31449_, _31448_);
  nor (_31450_, _31449_, _30412_);
  not (_31451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_31452_, _31448_, _31451_);
  or (_31453_, _31452_, _31450_);
  and (_31454_, _31453_, _27202_);
  nor (_31455_, _27201_, _31451_);
  or (_31456_, _31455_, rst);
  or (_31457_, _31456_, _31454_);
  or (_30239_, _31457_, _31447_);
  not (_31458_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_31459_, _31398_, _31458_);
  and (_31460_, _31398_, _28359_);
  or (_31461_, _31460_, _31459_);
  and (_31462_, _31461_, _27869_);
  and (_31463_, _31398_, _30471_);
  or (_31464_, _31463_, _31459_);
  and (_31465_, _31464_, _27202_);
  nor (_31466_, _27201_, _31458_);
  or (_31467_, _31466_, rst);
  or (_31468_, _31467_, _31465_);
  or (_33315_, _31468_, _31462_);
  nand (_31469_, _30418_, _27760_);
  or (_31470_, _30418_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31471_, _31470_, _27869_);
  and (_31472_, _31471_, _31469_);
  nand (_31473_, _31398_, _30462_);
  or (_31474_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31475_, _31474_, _27202_);
  and (_31476_, _31475_, _31473_);
  not (_31477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_31478_, _27201_, _31477_);
  or (_31479_, _31478_, rst);
  or (_31480_, _31479_, _31476_);
  or (_33317_, _31480_, _31472_);
  not (_31481_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not (_31482_, _29772_);
  and (_31483_, _30417_, _31482_);
  nor (_31484_, _31483_, _31481_);
  and (_31485_, _24331_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_31486_, _31485_, _29707_);
  and (_31487_, _31486_, _30417_);
  or (_31488_, _31487_, _31484_);
  and (_31489_, _31488_, _27869_);
  nand (_31490_, _31398_, _30455_);
  or (_31491_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_31492_, _31491_, _27202_);
  and (_31493_, _31492_, _31490_);
  nor (_31494_, _27201_, _31481_);
  or (_31495_, _31494_, rst);
  or (_31496_, _31495_, _31493_);
  or (_33319_, _31496_, _31489_);
  and (_31497_, _30417_, _29770_);
  nand (_31498_, _30417_, _24319_);
  or (_31499_, _31483_, _31498_);
  and (_31500_, _31499_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31501_, _31500_, _31497_);
  and (_31502_, _31501_, _27869_);
  nand (_31503_, _31398_, _30447_);
  or (_31504_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_31505_, _31504_, _27202_);
  and (_31506_, _31505_, _31503_);
  not (_31507_, _27201_);
  and (_31508_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31509_, _31508_, rst);
  or (_31510_, _31509_, _31506_);
  or (_33321_, _31510_, _31502_);
  and (_31511_, _30417_, _29840_);
  nand (_31512_, _31511_, _27760_);
  or (_31513_, _31511_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31514_, _31513_, _27869_);
  and (_31515_, _31514_, _31512_);
  nand (_31516_, _31398_, _30439_);
  or (_31517_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31518_, _31517_, _27202_);
  and (_31519_, _31518_, _31516_);
  and (_31520_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_31521_, _31520_, rst);
  or (_31522_, _31521_, _31519_);
  or (_33322_, _31522_, _31515_);
  and (_31523_, _30417_, _29916_);
  nand (_31524_, _31523_, _27760_);
  or (_31525_, _31523_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31526_, _31525_, _27869_);
  and (_31527_, _31526_, _31524_);
  nand (_31528_, _31398_, _30432_);
  or (_31529_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31530_, _31529_, _27202_);
  and (_31531_, _31530_, _31528_);
  and (_31532_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_31533_, _31532_, rst);
  or (_31534_, _31533_, _31531_);
  or (_33324_, _31534_, _31527_);
  nand (_31535_, _30417_, _29984_);
  and (_31536_, _31535_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_31537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_31538_, _27825_, _31537_);
  or (_31539_, _31538_, _29988_);
  and (_31540_, _31539_, _30417_);
  or (_31541_, _31540_, _31536_);
  and (_31542_, _31541_, _27869_);
  nand (_31543_, _31398_, _30425_);
  or (_31544_, _31398_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_31545_, _31544_, _27202_);
  and (_31546_, _31545_, _31543_);
  nor (_31547_, _27201_, _31537_);
  or (_31548_, _31547_, rst);
  or (_31549_, _31548_, _31546_);
  or (_33326_, _31549_, _31542_);
  nand (_31550_, _31414_, _27760_);
  or (_31551_, _31414_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_31552_, _31551_, _27869_);
  and (_31553_, _31552_, _31550_);
  and (_31554_, _31414_, _30471_);
  not (_31555_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_31556_, _31414_, _31555_);
  or (_31557_, _31556_, _31554_);
  and (_31558_, _31557_, _27202_);
  nor (_31559_, _27201_, _31555_);
  or (_31560_, _31559_, rst);
  or (_31561_, _31560_, _31558_);
  or (_33328_, _31561_, _31553_);
  and (_31562_, _31408_, _29027_);
  nand (_31563_, _31562_, _27760_);
  or (_31564_, _31562_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_31565_, _31564_, _27869_);
  and (_31566_, _31565_, _31563_);
  nor (_31567_, _31415_, _30462_);
  not (_31568_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_31569_, _31414_, _31568_);
  or (_31570_, _31569_, _31567_);
  and (_31571_, _31570_, _27202_);
  nor (_31572_, _27201_, _31568_);
  or (_31574_, _31572_, rst);
  or (_31575_, _31574_, _31571_);
  or (_33330_, _31575_, _31566_);
  and (_31576_, _31408_, _29706_);
  nand (_31577_, _31576_, _27760_);
  or (_31578_, _31576_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_31579_, _31578_, _27869_);
  and (_31580_, _31579_, _31577_);
  nor (_31581_, _31415_, _30455_);
  not (_31582_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_31583_, _31414_, _31582_);
  or (_31584_, _31583_, _31581_);
  and (_31585_, _31584_, _27202_);
  nor (_31586_, _27201_, _31582_);
  or (_31587_, _31586_, rst);
  or (_31588_, _31587_, _31585_);
  or (_33332_, _31588_, _31580_);
  and (_31589_, _31408_, _29769_);
  nand (_31590_, _31589_, _27760_);
  or (_31591_, _31589_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_31592_, _31591_, _27869_);
  and (_31593_, _31592_, _31590_);
  nor (_31594_, _31415_, _30447_);
  and (_31595_, _31415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31596_, _31595_, _31594_);
  and (_31597_, _31596_, _27202_);
  and (_31598_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31599_, _31598_, rst);
  or (_31600_, _31599_, _31597_);
  or (_33333_, _31600_, _31593_);
  and (_31602_, _31408_, _29840_);
  nand (_31606_, _31602_, _27760_);
  or (_31607_, _31602_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_31608_, _31607_, _27869_);
  and (_31609_, _31608_, _31606_);
  nor (_31610_, _31415_, _30439_);
  and (_31611_, _31415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31612_, _31611_, _31610_);
  and (_31613_, _31612_, _27202_);
  and (_31614_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31615_, _31614_, rst);
  or (_31616_, _31615_, _31613_);
  or (_33335_, _31616_, _31609_);
  and (_31617_, _31408_, _29916_);
  nand (_31618_, _31617_, _27760_);
  or (_31619_, _31617_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_31620_, _31619_, _27869_);
  and (_31621_, _31620_, _31618_);
  nor (_31622_, _31415_, _30432_);
  and (_31623_, _31415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31624_, _31623_, _31622_);
  and (_31625_, _31624_, _27202_);
  and (_31626_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31627_, _31626_, rst);
  or (_31628_, _31627_, _31625_);
  or (_33337_, _31628_, _31621_);
  and (_31629_, _31408_, _29987_);
  nand (_31630_, _31629_, _27760_);
  or (_31631_, _31629_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_31632_, _31631_, _27869_);
  and (_31633_, _31632_, _31630_);
  nor (_31634_, _31415_, _30425_);
  not (_31635_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_31636_, _31414_, _31635_);
  or (_31637_, _31636_, _31634_);
  and (_31638_, _31637_, _27202_);
  nor (_31639_, _27201_, _31635_);
  or (_31640_, _31639_, rst);
  or (_31641_, _31640_, _31638_);
  or (_33339_, _31641_, _31633_);
  and (_31642_, _31425_, _24343_);
  nand (_31643_, _31642_, _27760_);
  or (_31644_, _31642_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_31645_, _31644_, _27869_);
  and (_31646_, _31645_, _31643_);
  nor (_31647_, _31433_, _30470_);
  not (_31648_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_31649_, _31432_, _31648_);
  or (_31650_, _31649_, _31647_);
  and (_31651_, _31650_, _27202_);
  nor (_31652_, _27201_, _31648_);
  or (_31653_, _31652_, rst);
  or (_31654_, _31653_, _31651_);
  or (_33341_, _31654_, _31646_);
  and (_31655_, _31425_, _29027_);
  nand (_31656_, _31655_, _27760_);
  or (_31657_, _31655_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_31658_, _31657_, _27869_);
  and (_31659_, _31658_, _31656_);
  nor (_31660_, _31433_, _30462_);
  not (_31661_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_31662_, _31432_, _31661_);
  or (_31663_, _31662_, _31660_);
  and (_31665_, _31663_, _27202_);
  nor (_31672_, _27201_, _31661_);
  or (_31673_, _31672_, rst);
  or (_31674_, _31673_, _31665_);
  or (_33343_, _31674_, _31659_);
  and (_31675_, _31425_, _29706_);
  nand (_31676_, _31675_, _27760_);
  or (_31677_, _31675_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_31678_, _31677_, _27869_);
  and (_31679_, _31678_, _31676_);
  nor (_31680_, _31433_, _30455_);
  not (_31681_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_31682_, _31432_, _31681_);
  or (_31683_, _31682_, _31680_);
  and (_31684_, _31683_, _27202_);
  nor (_31685_, _27201_, _31681_);
  or (_31686_, _31685_, rst);
  or (_31687_, _31686_, _31684_);
  or (_33344_, _31687_, _31679_);
  and (_31688_, _31425_, _29769_);
  nand (_31689_, _31688_, _27760_);
  or (_31690_, _31688_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_31691_, _31690_, _27869_);
  and (_31692_, _31691_, _31689_);
  nor (_31693_, _31433_, _30447_);
  and (_31694_, _31433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31695_, _31694_, _31693_);
  and (_31696_, _31695_, _27202_);
  and (_31697_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31698_, _31697_, rst);
  or (_31699_, _31698_, _31696_);
  or (_33346_, _31699_, _31692_);
  and (_31700_, _31425_, _29840_);
  nand (_31701_, _31700_, _27760_);
  or (_31702_, _31700_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_31703_, _31702_, _27869_);
  and (_31704_, _31703_, _31701_);
  nor (_31705_, _31433_, _30439_);
  and (_31706_, _31433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31707_, _31706_, _31705_);
  and (_31708_, _31707_, _27202_);
  and (_31709_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31710_, _31709_, rst);
  or (_31711_, _31710_, _31708_);
  or (_33348_, _31711_, _31704_);
  and (_31712_, _31425_, _29916_);
  nand (_31713_, _31712_, _27760_);
  or (_31714_, _31712_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_31719_, _31714_, _27869_);
  and (_31720_, _31719_, _31713_);
  nor (_31721_, _31433_, _30432_);
  and (_31722_, _31433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31723_, _31722_, _31721_);
  and (_31724_, _31723_, _27202_);
  and (_31725_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31726_, _31725_, rst);
  or (_31727_, _31726_, _31724_);
  or (_33350_, _31727_, _31720_);
  and (_31728_, _31425_, _29987_);
  nand (_31729_, _31728_, _27760_);
  or (_31730_, _31728_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_31731_, _31730_, _27869_);
  and (_31732_, _31731_, _31729_);
  nor (_31735_, _31433_, _30425_);
  not (_31743_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_31744_, _31432_, _31743_);
  or (_31745_, _31744_, _31735_);
  and (_31746_, _31745_, _27202_);
  nor (_31747_, _27201_, _31743_);
  or (_31748_, _31747_, rst);
  or (_31749_, _31748_, _31746_);
  or (_33352_, _31749_, _31732_);
  and (_31750_, _31442_, _24343_);
  nand (_31751_, _31750_, _27760_);
  or (_31752_, _31750_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_31753_, _31752_, _27869_);
  and (_31754_, _31753_, _31751_);
  nor (_31755_, _31449_, _30470_);
  not (_31756_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_31757_, _31448_, _31756_);
  or (_31758_, _31757_, _31755_);
  and (_31759_, _31758_, _27202_);
  nor (_31760_, _27201_, _31756_);
  or (_31761_, _31760_, rst);
  or (_31762_, _31761_, _31759_);
  or (_33354_, _31762_, _31754_);
  and (_31763_, _31442_, _29027_);
  nand (_31764_, _31763_, _27760_);
  or (_31765_, _31763_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_31766_, _31765_, _27869_);
  and (_31767_, _31766_, _31764_);
  nor (_31768_, _31449_, _30462_);
  not (_31769_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_31770_, _31448_, _31769_);
  or (_31771_, _31770_, _31768_);
  and (_31772_, _31771_, _27202_);
  nor (_31773_, _27201_, _31769_);
  or (_31774_, _31773_, rst);
  or (_31775_, _31774_, _31772_);
  or (_33355_, _31775_, _31767_);
  and (_31776_, _31442_, _29706_);
  nand (_31777_, _31776_, _27760_);
  or (_31778_, _31776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_31779_, _31778_, _27869_);
  and (_31780_, _31779_, _31777_);
  nor (_31781_, _31449_, _30455_);
  not (_31782_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_31783_, _31448_, _31782_);
  or (_31784_, _31783_, _31781_);
  and (_31785_, _31784_, _27202_);
  nor (_31786_, _27201_, _31782_);
  or (_31787_, _31786_, rst);
  or (_31788_, _31787_, _31785_);
  or (_33357_, _31788_, _31780_);
  and (_31789_, _31442_, _29769_);
  nand (_31790_, _31789_, _27760_);
  or (_31791_, _31789_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_31792_, _31791_, _27869_);
  and (_31793_, _31792_, _31790_);
  nor (_31794_, _31449_, _30447_);
  and (_31795_, _31449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31796_, _31795_, _31794_);
  and (_31797_, _31796_, _27202_);
  and (_31798_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31799_, _31798_, rst);
  or (_31800_, _31799_, _31797_);
  or (_33359_, _31800_, _31793_);
  and (_31801_, _31442_, _29840_);
  nand (_31802_, _31801_, _27760_);
  or (_31803_, _31801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_31804_, _31803_, _27869_);
  and (_31805_, _31804_, _31802_);
  nor (_31806_, _31449_, _30439_);
  and (_31807_, _31449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31808_, _31807_, _31806_);
  and (_31809_, _31808_, _27202_);
  and (_31810_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31811_, _31810_, rst);
  or (_31812_, _31811_, _31809_);
  or (_33361_, _31812_, _31805_);
  and (_31813_, _31442_, _29916_);
  nand (_31814_, _31813_, _27760_);
  or (_31815_, _31813_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_31816_, _31815_, _27869_);
  and (_31817_, _31816_, _31814_);
  nor (_31818_, _31449_, _30432_);
  and (_31819_, _31449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31820_, _31819_, _31818_);
  and (_31821_, _31820_, _27202_);
  and (_31822_, _31507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31823_, _31822_, rst);
  or (_31824_, _31823_, _31821_);
  or (_33363_, _31824_, _31817_);
  and (_31825_, _31442_, _29987_);
  nand (_31826_, _31825_, _27760_);
  or (_31827_, _31825_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_31828_, _31827_, _27869_);
  and (_31829_, _31828_, _31826_);
  nor (_31830_, _31449_, _30425_);
  not (_31831_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_31832_, _31448_, _31831_);
  or (_31833_, _31832_, _31830_);
  and (_31834_, _31833_, _27202_);
  nor (_31835_, _27201_, _31831_);
  or (_31836_, _31835_, rst);
  or (_31837_, _31836_, _31834_);
  or (_33365_, _31837_, _31829_);
  and (_31838_, _30345_, _30274_);
  nor (_31839_, _30301_, _30289_);
  nor (_31840_, _30317_, _30305_);
  and (_31841_, _31840_, _30299_);
  and (_31842_, _31841_, _31839_);
  not (_31843_, _30313_);
  and (_31844_, _30334_, _31843_);
  and (_31845_, _31844_, _30346_);
  and (_31846_, _31845_, _31842_);
  nor (_31847_, _31846_, _29998_);
  nor (_31848_, _31847_, _31838_);
  not (_31849_, _31848_);
  and (_31850_, _30394_, _30282_);
  and (_31851_, _31850_, _30377_);
  and (_31852_, _31851_, _30284_);
  not (_31853_, _30282_);
  nor (_31854_, _30377_, _31853_);
  and (_31855_, _31854_, _30394_);
  not (_31856_, _30002_);
  and (_31857_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_31858_, _30093_, _30002_);
  not (_31859_, _31858_);
  and (_31860_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_31861_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_31862_, _31861_, _31860_);
  and (_31863_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_31864_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_31865_, _31864_, _31863_);
  and (_31866_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_31867_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_31868_, _31867_, _31866_);
  and (_31869_, _31868_, _31865_);
  and (_31870_, _31869_, _31862_);
  nor (_31871_, _31870_, _31859_);
  nor (_31872_, _31871_, _31857_);
  not (_31873_, _31872_);
  and (_31874_, _31873_, _31855_);
  nor (_31875_, _31874_, _31852_);
  and (_31876_, _30394_, _30378_);
  not (_31877_, _30508_);
  and (_31878_, _31877_, _31876_);
  and (_31879_, _30377_, _31853_);
  and (_31880_, _31879_, _30394_);
  and (_31881_, _30211_, _27814_);
  nor (_31882_, _31881_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_31883_, _23420_, _23036_);
  nor (_31884_, _31883_, _27180_);
  not (_31885_, _24331_);
  nor (_31886_, _30211_, _27814_);
  nor (_31887_, _31886_, _31885_);
  and (_31888_, _31887_, _31884_);
  and (_31889_, _31888_, _31882_);
  not (_31890_, _23606_);
  nor (_31891_, _30990_, _31040_);
  nor (_31892_, _31891_, _31046_);
  nor (_31893_, _31892_, _31890_);
  and (_31894_, _31892_, _31890_);
  nor (_31895_, _31894_, _31893_);
  and (_31896_, _31895_, _31889_);
  nor (_31897_, _31892_, _30211_);
  and (_31898_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_31899_, _31892_, _30245_);
  and (_31900_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_31901_, _31900_, _31898_);
  and (_31902_, _31892_, _30211_);
  and (_31903_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_31904_, _31892_, _30245_);
  and (_31905_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_31906_, _31905_, _31903_);
  and (_31907_, _31906_, _31901_);
  nor (_31908_, _31907_, _31896_);
  not (_31909_, _30455_);
  and (_31910_, _31896_, _31909_);
  nor (_31911_, _31910_, _31908_);
  not (_31912_, _31911_);
  and (_31913_, _31912_, _31880_);
  nor (_31914_, _31913_, _31878_);
  and (_31915_, _31914_, _31875_);
  nor (_31916_, _31915_, _31849_);
  not (_31917_, _30526_);
  and (_31918_, _31917_, _31876_);
  and (_31919_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_31920_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_31921_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_31922_, _31921_, _31920_);
  and (_31923_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_31924_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_31925_, _31924_, _31923_);
  and (_31926_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_31927_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_31928_, _31927_, _31926_);
  and (_31929_, _31928_, _31925_);
  and (_31930_, _31929_, _31922_);
  nor (_31931_, _31930_, _31859_);
  nor (_31932_, _31931_, _31919_);
  not (_31933_, _31932_);
  and (_31934_, _31933_, _31855_);
  nor (_31935_, _31934_, _31918_);
  and (_31936_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_31937_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_31938_, _31937_, _31936_);
  and (_31939_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_31940_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_31941_, _31940_, _31939_);
  and (_31942_, _31941_, _31938_);
  nor (_31943_, _31942_, _31896_);
  not (_31944_, _30432_);
  and (_31945_, _31896_, _31944_);
  nor (_31946_, _31945_, _31943_);
  not (_31947_, _31946_);
  and (_31948_, _31947_, _31880_);
  not (_31949_, _31854_);
  nor (_31950_, _31879_, _30394_);
  and (_31951_, _31950_, _31949_);
  nor (_31952_, _31951_, _31948_);
  and (_31953_, _31952_, _31935_);
  not (_31954_, _31953_);
  and (_31955_, _30259_, _30343_);
  nor (_31956_, _30369_, _31955_);
  nor (_31957_, _31956_, _30365_);
  not (_31958_, _30332_);
  and (_31959_, _30366_, _30089_);
  and (_31960_, _31959_, _30259_);
  nor (_31961_, _31960_, _30289_);
  and (_31962_, _31961_, _31958_);
  and (_31963_, _31962_, _31843_);
  and (_31964_, _31959_, _30215_);
  not (_31965_, _31964_);
  and (_31966_, _31965_, _31956_);
  not (_31967_, _30368_);
  and (_31968_, _30264_, _30222_);
  and (_31969_, _31968_, _30215_);
  nor (_31970_, _31969_, _30296_);
  and (_31971_, _31970_, _31967_);
  and (_31972_, _31971_, _31966_);
  and (_31973_, _31972_, _31963_);
  and (_31974_, _31973_, _31840_);
  nor (_31975_, _31974_, _29998_);
  nor (_31976_, _31975_, _31957_);
  not (_31977_, _30488_);
  and (_31978_, _31977_, _31876_);
  not (_31979_, _31978_);
  and (_31980_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_31981_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_31982_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_31983_, _31982_, _31981_);
  and (_31984_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_31985_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_31986_, _31985_, _31984_);
  and (_31987_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_31988_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_31989_, _31988_, _31987_);
  and (_31990_, _31989_, _31986_);
  and (_31991_, _31990_, _31983_);
  nor (_31992_, _31991_, _31859_);
  nor (_31993_, _31992_, _31980_);
  not (_31994_, _31993_);
  and (_31995_, _31994_, _31854_);
  not (_31996_, _31995_);
  not (_31997_, _30394_);
  and (_31998_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  not (_31999_, _31998_);
  and (_32000_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_32001_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_32002_, _32001_, _32000_);
  and (_32003_, _32002_, _31999_);
  and (_32004_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_32005_, _32004_, _31896_);
  and (_32006_, _32005_, _32003_);
  and (_32007_, _31896_, _30412_);
  or (_32008_, _32007_, _32006_);
  not (_32009_, _32008_);
  and (_32010_, _32009_, _31879_);
  nor (_32011_, _32010_, _31997_);
  and (_32012_, _32011_, _31996_);
  and (_32013_, _32012_, _31979_);
  not (_32014_, _32013_);
  nor (_32015_, _32014_, _31976_);
  and (_32016_, _32015_, _31954_);
  nor (_32017_, _32016_, _31916_);
  and (_32018_, _23420_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32019_, _32018_, _23935_);
  nor (_32020_, _24319_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32021_, _32020_, _32019_);
  not (_32022_, _32021_);
  and (_32023_, _32022_, _32017_);
  and (_32024_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  not (_32025_, _32024_);
  and (_32026_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_32027_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_32028_, _32027_, _32026_);
  and (_32029_, _32028_, _32025_);
  and (_32030_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_32031_, _32030_, _31896_);
  and (_32032_, _32031_, _32029_);
  and (_32033_, _31896_, _30470_);
  or (_32034_, _32033_, _32032_);
  not (_32035_, _32034_);
  and (_32036_, _32035_, _31880_);
  and (_32037_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_32038_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_32039_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_32040_, _32039_, _32038_);
  and (_32041_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_32042_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_32043_, _32042_, _32041_);
  and (_32044_, _32043_, _32040_);
  and (_32045_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_32046_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_32047_, _32046_, _32045_);
  and (_32048_, _32047_, _32044_);
  nor (_32049_, _32048_, _31859_);
  nor (_32050_, _32049_, _32037_);
  not (_32051_, _32050_);
  and (_32052_, _32051_, _31855_);
  nor (_32053_, _32052_, _32036_);
  not (_32054_, _30496_);
  and (_32055_, _32054_, _31876_);
  and (_32056_, _31851_, _30245_);
  nor (_32057_, _32056_, _32055_);
  and (_32058_, _32057_, _32053_);
  nor (_32059_, _32058_, _31849_);
  not (_32060_, _31892_);
  and (_32061_, _32060_, _31851_);
  and (_32062_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_32063_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_32064_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_32065_, _32064_, _32063_);
  and (_32066_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_32067_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_32068_, _32067_, _32066_);
  and (_32069_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_32070_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_32071_, _32070_, _32069_);
  and (_32072_, _32071_, _32068_);
  and (_32073_, _32072_, _32065_);
  nor (_32074_, _32073_, _31859_);
  nor (_32075_, _32074_, _32062_);
  not (_32076_, _32075_);
  and (_32077_, _32076_, _31855_);
  nor (_32078_, _32077_, _32061_);
  not (_32079_, _30514_);
  and (_32080_, _32079_, _31876_);
  and (_32081_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_32082_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_32083_, _32082_, _32081_);
  and (_32084_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_32085_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_32086_, _32085_, _32084_);
  and (_32087_, _32086_, _32083_);
  nor (_32088_, _32087_, _31896_);
  not (_32089_, _30447_);
  and (_32090_, _31896_, _32089_);
  nor (_32091_, _32090_, _32088_);
  not (_32092_, _32091_);
  and (_32093_, _32092_, _31880_);
  nor (_32094_, _32093_, _32080_);
  and (_32095_, _32094_, _32078_);
  not (_32096_, _32095_);
  and (_32097_, _32096_, _32015_);
  nor (_32098_, _32097_, _32059_);
  and (_32099_, _32018_, _31890_);
  nor (_32100_, _24056_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32101_, _32100_, _32099_);
  not (_32102_, _32101_);
  nor (_32103_, _32102_, _32098_);
  nor (_32104_, _32103_, _32023_);
  nor (_32105_, _32022_, _32017_);
  not (_32106_, _32105_);
  and (_32107_, _32013_, _31849_);
  nor (_32108_, _32096_, _32107_);
  not (_32109_, _30532_);
  and (_32110_, _32109_, _31876_);
  not (_32111_, _30425_);
  and (_32112_, _31896_, _32111_);
  and (_32113_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_32114_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_32115_, _32114_, _32113_);
  and (_32116_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_32117_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_32118_, _32117_, _32116_);
  and (_32119_, _32118_, _32115_);
  nor (_32120_, _32119_, _31896_);
  nor (_32121_, _32120_, _32112_);
  not (_32122_, _32121_);
  and (_32123_, _32122_, _31880_);
  and (_32124_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_32125_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_32126_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_32127_, _32126_, _32125_);
  and (_32128_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_32129_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_32130_, _32129_, _32128_);
  and (_32131_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_32132_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_32133_, _32132_, _32131_);
  and (_32134_, _32133_, _32130_);
  and (_32135_, _32134_, _32127_);
  nor (_32136_, _32135_, _31859_);
  nor (_32137_, _32136_, _32124_);
  not (_32138_, _32137_);
  and (_32139_, _32138_, _31854_);
  or (_32140_, _32139_, _32123_);
  or (_32141_, _32140_, _32110_);
  nor (_32142_, _32141_, _31950_);
  and (_32143_, _32142_, _32107_);
  nor (_32144_, _32143_, _32108_);
  and (_32145_, _32018_, _23287_);
  nor (_32146_, _32018_, _31890_);
  nor (_32147_, _32146_, _32145_);
  not (_32148_, _32147_);
  and (_32149_, _32148_, _32144_);
  nor (_32150_, _32148_, _32144_);
  nor (_32151_, _32150_, _32149_);
  and (_32152_, _32151_, _32106_);
  and (_32153_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_32154_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_32155_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_32156_, _32155_, _32154_);
  and (_32157_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_32158_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_32159_, _32158_, _32157_);
  and (_32160_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_32161_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_32162_, _32161_, _32160_);
  and (_32163_, _32162_, _32159_);
  and (_32164_, _32163_, _32156_);
  nor (_32165_, _32164_, _31859_);
  nor (_32166_, _32165_, _32153_);
  not (_32167_, _32166_);
  and (_32168_, _32167_, _31855_);
  and (_32169_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  not (_32170_, _32169_);
  and (_32171_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_32172_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32173_, _32172_, _32171_);
  and (_32174_, _32173_, _32170_);
  and (_32175_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_32176_, _32175_, _31896_);
  and (_32177_, _32176_, _32174_);
  and (_32178_, _31896_, _30462_);
  or (_32179_, _32178_, _32177_);
  not (_32180_, _32179_);
  and (_32181_, _32180_, _31880_);
  nor (_32182_, _32181_, _32168_);
  not (_32183_, _30502_);
  and (_32184_, _32183_, _31876_);
  not (_32185_, _32184_);
  and (_32186_, _31879_, _31997_);
  and (_32187_, _31851_, _30212_);
  nor (_32188_, _32187_, _32186_);
  and (_32189_, _32188_, _32185_);
  and (_32190_, _32189_, _32182_);
  nor (_32191_, _32190_, _31849_);
  and (_32192_, _31856_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_32193_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_32194_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_32195_, _32194_, _32193_);
  and (_32196_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_32197_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_32198_, _32197_, _32196_);
  and (_32199_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_32200_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_32201_, _32200_, _32199_);
  and (_32202_, _32201_, _32198_);
  and (_32203_, _32202_, _32195_);
  nor (_32204_, _32203_, _31859_);
  nor (_32205_, _32204_, _32192_);
  not (_32206_, _32205_);
  and (_32207_, _32206_, _31855_);
  or (_32208_, _31055_, _31051_);
  and (_32209_, _32208_, _31851_);
  nor (_32210_, _32209_, _32207_);
  and (_32211_, _31897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_32212_, _31899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_32213_, _32212_, _32211_);
  and (_32214_, _31902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_32215_, _31904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_32216_, _32215_, _32214_);
  and (_32217_, _32216_, _32213_);
  nor (_32218_, _32217_, _31896_);
  not (_32219_, _30439_);
  and (_32220_, _31896_, _32219_);
  nor (_32221_, _32220_, _32218_);
  not (_32222_, _32221_);
  and (_32223_, _32222_, _31880_);
  not (_32224_, _32223_);
  and (_32225_, _31997_, _30282_);
  not (_32226_, _30520_);
  and (_32227_, _32226_, _31876_);
  nor (_32228_, _32227_, _32225_);
  and (_32229_, _32228_, _32224_);
  and (_32230_, _32229_, _32210_);
  not (_32231_, _32230_);
  and (_32232_, _32231_, _32015_);
  nor (_32233_, _32232_, _32191_);
  and (_32234_, _32018_, _23781_);
  nor (_32235_, _24187_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_32236_, _32235_, _32234_);
  nand (_32237_, _32236_, _32233_);
  or (_32238_, _32236_, _32233_);
  and (_32239_, _32238_, _32237_);
  not (_32240_, _32239_);
  not (_32241_, _31884_);
  and (_32242_, _32102_, _32098_);
  nor (_32243_, _32242_, _32241_);
  and (_32244_, _32243_, _32240_);
  and (_32245_, _32244_, _32152_);
  and (_32246_, _32245_, _32104_);
  not (_32247_, _32017_);
  and (_32248_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_32249_, _32098_);
  and (_32250_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_32251_, _32250_, _32248_);
  and (_32252_, _32251_, _32233_);
  not (_32253_, _32233_);
  not (_32254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_32255_, _32098_, _32254_);
  and (_32256_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_32257_, _32256_, _32255_);
  and (_32258_, _32257_, _32253_);
  or (_32259_, _32258_, _32252_);
  or (_32260_, _32259_, _32247_);
  not (_32261_, _32144_);
  and (_32262_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_32263_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_32264_, _32263_, _32262_);
  and (_32265_, _32264_, _32233_);
  not (_32266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_32267_, _32098_, _32266_);
  and (_32268_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_32269_, _32268_, _32267_);
  and (_32270_, _32269_, _32253_);
  or (_32271_, _32270_, _32265_);
  or (_32272_, _32271_, _32017_);
  and (_32273_, _32272_, _32261_);
  and (_32274_, _32273_, _32260_);
  or (_32275_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_32276_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_32277_, _32276_, _32275_);
  and (_32278_, _32277_, _32233_);
  or (_32279_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_32280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_32281_, _32098_, _32280_);
  and (_32282_, _32281_, _32279_);
  and (_32283_, _32282_, _32253_);
  or (_32284_, _32283_, _32278_);
  or (_32285_, _32284_, _32247_);
  or (_32286_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_32287_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_32288_, _32287_, _32286_);
  and (_32289_, _32288_, _32233_);
  or (_32290_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_32291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_32292_, _32098_, _32291_);
  and (_32293_, _32292_, _32290_);
  and (_32294_, _32293_, _32253_);
  or (_32295_, _32294_, _32289_);
  or (_32296_, _32295_, _32017_);
  and (_32297_, _32296_, _32144_);
  and (_32298_, _32297_, _32285_);
  or (_32299_, _32298_, _32274_);
  or (_32300_, _32299_, _32246_);
  not (_32301_, _32246_);
  or (_32302_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_32303_, _32302_, _36029_);
  and (_33440_, _32303_, _32300_);
  nor (_32304_, _32101_, _32241_);
  nor (_32305_, _32236_, _32241_);
  and (_32306_, _32305_, _32304_);
  and (_32307_, _32147_, _31884_);
  nor (_32308_, _32021_, _32241_);
  and (_32309_, _32308_, _32307_);
  and (_32310_, _32309_, _32306_);
  and (_32311_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_32312_, _32311_, _25247_);
  nor (_32313_, _32312_, _27760_);
  nand (_32314_, _25247_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32315_, _16525_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32316_, _32315_, _32314_);
  nor (_32317_, _30412_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32318_, _32317_, _32316_);
  or (_32319_, _32318_, _32313_);
  and (_32320_, _32319_, _31884_);
  and (_32321_, _32320_, _32310_);
  not (_32322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_32323_, _32310_, _32322_);
  or (_33450_, _32323_, _32321_);
  nor (_32324_, _32308_, _32307_);
  nor (_32325_, _32305_, _32304_);
  and (_32326_, _32325_, _31884_);
  and (_32327_, _32326_, _32324_);
  and (_32328_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25149_);
  and (_32329_, _32328_, _25204_);
  not (_32330_, _32329_);
  nor (_32331_, _32330_, _27760_);
  not (_32332_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_32333_, _30470_, _32332_);
  or (_32334_, _15371_, _32332_);
  and (_32335_, _32334_, _32330_);
  and (_32336_, _32335_, _32333_);
  or (_32337_, _32336_, _32331_);
  and (_32338_, _32337_, _32327_);
  not (_32339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_32340_, _32327_, _32339_);
  or (_33693_, _32340_, _32338_);
  nand (_32341_, _32328_, _25270_);
  nor (_32342_, _32341_, _27760_);
  nor (_32343_, _30462_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32344_, _32328_, _25160_);
  and (_32345_, _32328_, _25247_);
  or (_32346_, _32345_, _32311_);
  or (_32347_, _32346_, _32344_);
  and (_32348_, _32347_, _16351_);
  or (_32349_, _32348_, _32343_);
  or (_32350_, _32349_, _32342_);
  and (_32351_, _32350_, _32327_);
  not (_32352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_32353_, _32327_, _32352_);
  or (_33698_, _32353_, _32351_);
  not (_32354_, _32327_);
  and (_32355_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_32356_, _32328_, _25171_);
  nor (_32357_, _32356_, _27760_);
  nor (_32358_, _30455_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32359_, _32328_, _25259_);
  or (_32360_, _32359_, _32346_);
  and (_32361_, _32360_, _15009_);
  or (_32362_, _32361_, _32358_);
  or (_32363_, _32362_, _32357_);
  and (_32364_, _32363_, _32327_);
  or (_33703_, _32364_, _32355_);
  and (_32365_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_32366_, _32345_, _28359_);
  nor (_32367_, _30447_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32368_, _32344_, _32311_);
  or (_32369_, _32368_, _32359_);
  and (_32370_, _32369_, _16035_);
  or (_32371_, _32370_, _32367_);
  or (_32372_, _32371_, _32366_);
  and (_32373_, _32372_, _32327_);
  or (_33709_, _32373_, _32365_);
  and (_32374_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_32375_, _32311_, _25204_);
  nor (_32376_, _32375_, _27760_);
  nor (_32377_, _30439_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_32378_, _25204_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32379_, _15206_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32380_, _32379_, _32378_);
  or (_32381_, _32380_, _32377_);
  or (_32382_, _32381_, _32376_);
  and (_32383_, _32382_, _32327_);
  or (_33714_, _32383_, _32374_);
  nand (_32384_, _32311_, _25270_);
  nor (_32385_, _32384_, _27760_);
  nor (_32386_, _30432_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_32387_, _25270_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32388_, _16187_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32389_, _32388_, _32387_);
  or (_32390_, _32389_, _32386_);
  or (_32391_, _32390_, _32385_);
  and (_32392_, _32391_, _32327_);
  and (_32393_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_33719_, _32393_, _32392_);
  and (_32394_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_32395_, _32311_, _25171_);
  nor (_32396_, _32395_, _27760_);
  nor (_32397_, _30425_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_32398_, _25171_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_32399_, _15545_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32400_, _32399_, _32398_);
  or (_32401_, _32400_, _32397_);
  or (_32402_, _32401_, _32396_);
  and (_32403_, _32402_, _32327_);
  or (_33724_, _32403_, _32394_);
  and (_32404_, _32327_, _32319_);
  and (_32405_, _32354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_33727_, _32405_, _32404_);
  and (_32406_, _32337_, _31884_);
  and (_32407_, _32304_, _32236_);
  and (_32408_, _32407_, _32324_);
  and (_32409_, _32408_, _32406_);
  not (_32410_, _32408_);
  and (_32411_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_33734_, _32411_, _32409_);
  and (_32412_, _32350_, _31884_);
  and (_32413_, _32408_, _32412_);
  and (_32414_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_33737_, _32414_, _32413_);
  and (_32415_, _32363_, _31884_);
  and (_32416_, _32408_, _32415_);
  and (_32417_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_33741_, _32417_, _32416_);
  and (_32418_, _32372_, _31884_);
  and (_32419_, _32408_, _32418_);
  and (_32420_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_33744_, _32420_, _32419_);
  and (_32421_, _32382_, _31884_);
  and (_32422_, _32408_, _32421_);
  not (_32423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_32424_, _32408_, _32423_);
  or (_33748_, _32424_, _32422_);
  and (_32425_, _32391_, _31884_);
  and (_32426_, _32408_, _32425_);
  not (_32427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_32428_, _32408_, _32427_);
  or (_33751_, _32428_, _32426_);
  and (_32429_, _32402_, _31884_);
  and (_32430_, _32408_, _32429_);
  and (_32431_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_33755_, _32431_, _32430_);
  and (_32432_, _32408_, _32320_);
  and (_32433_, _32410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_33757_, _32433_, _32432_);
  and (_32434_, _32305_, _32101_);
  and (_32435_, _32434_, _32324_);
  and (_32436_, _32435_, _32406_);
  not (_32437_, _32435_);
  and (_32438_, _32437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_33764_, _32438_, _32436_);
  and (_32439_, _32435_, _32412_);
  and (_32440_, _32437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_33768_, _32440_, _32439_);
  and (_32441_, _32435_, _32415_);
  not (_32442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_32443_, _32435_, _32442_);
  or (_33771_, _32443_, _32441_);
  and (_32444_, _32435_, _32418_);
  and (_32445_, _32437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_33775_, _32445_, _32444_);
  and (_32446_, _32435_, _32421_);
  not (_32447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_32448_, _32435_, _32447_);
  or (_33778_, _32448_, _32446_);
  and (_32449_, _32435_, _32425_);
  not (_32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_32451_, _32435_, _32450_);
  or (_33782_, _32451_, _32449_);
  and (_32452_, _32435_, _32429_);
  and (_32453_, _32437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_33785_, _32453_, _32452_);
  and (_32454_, _32435_, _32320_);
  not (_32455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_32456_, _32435_, _32455_);
  or (_33788_, _32456_, _32454_);
  and (_32457_, _32324_, _32306_);
  and (_32458_, _32457_, _32406_);
  not (_32459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_32460_, _32457_, _32459_);
  or (_33793_, _32460_, _32458_);
  and (_32461_, _32457_, _32412_);
  not (_32462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_32463_, _32457_, _32462_);
  or (_33797_, _32463_, _32461_);
  and (_32464_, _32457_, _32415_);
  not (_32465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_32466_, _32457_, _32465_);
  or (_33800_, _32466_, _32464_);
  and (_32467_, _32457_, _32418_);
  not (_32468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_32469_, _32457_, _32468_);
  or (_33804_, _32469_, _32467_);
  and (_32470_, _32457_, _32421_);
  not (_32471_, _32457_);
  and (_32472_, _32471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_33807_, _32472_, _32470_);
  and (_32473_, _32457_, _32425_);
  and (_32474_, _32471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_33811_, _32474_, _32473_);
  and (_32475_, _32457_, _32429_);
  and (_32476_, _32471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_33814_, _32476_, _32475_);
  and (_32477_, _32457_, _32320_);
  nor (_32478_, _32457_, _32254_);
  or (_33817_, _32478_, _32477_);
  and (_32479_, _32308_, _32148_);
  and (_32480_, _32479_, _32325_);
  and (_32481_, _32480_, _32406_);
  not (_32482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_32483_, _32480_, _32482_);
  or (_33824_, _32483_, _32481_);
  and (_32494_, _32480_, _32412_);
  not (_32502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_32511_, _32480_, _32502_);
  or (_33827_, _32511_, _32494_);
  and (_32514_, _32480_, _32415_);
  not (_32515_, _32480_);
  and (_32516_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_33831_, _32516_, _32514_);
  and (_32517_, _32480_, _32418_);
  and (_32518_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_33834_, _32518_, _32517_);
  and (_32519_, _32480_, _32421_);
  and (_32520_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_33838_, _32520_, _32519_);
  and (_32521_, _32480_, _32425_);
  and (_32522_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_33841_, _32522_, _32521_);
  and (_32523_, _32480_, _32429_);
  and (_32524_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_33845_, _32524_, _32523_);
  and (_32525_, _32480_, _32320_);
  and (_32526_, _32515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_33848_, _32526_, _32525_);
  and (_32527_, _32479_, _32407_);
  and (_32528_, _32527_, _32406_);
  not (_32529_, _32527_);
  and (_32530_, _32529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_33852_, _32530_, _32528_);
  and (_32531_, _32527_, _32412_);
  and (_32532_, _32529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_33855_, _32532_, _32531_);
  and (_32533_, _32527_, _32415_);
  and (_32534_, _32529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_33859_, _32534_, _32533_);
  and (_32535_, _32527_, _32418_);
  not (_32536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_32537_, _32527_, _32536_);
  or (_33862_, _32537_, _32535_);
  and (_32538_, _32527_, _32421_);
  not (_32539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_32542_, _32527_, _32539_);
  or (_33866_, _32542_, _32538_);
  and (_32548_, _32527_, _32425_);
  not (_32550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_32551_, _32527_, _32550_);
  or (_33869_, _32551_, _32548_);
  and (_32555_, _32527_, _32429_);
  not (_32561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_32562_, _32527_, _32561_);
  or (_33873_, _32562_, _32555_);
  and (_32563_, _32527_, _32320_);
  and (_32569_, _32529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_33876_, _32569_, _32563_);
  and (_32573_, _32479_, _32434_);
  and (_32574_, _32573_, _32406_);
  not (_32578_, _32573_);
  and (_32584_, _32578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_33880_, _32584_, _32574_);
  and (_32585_, _32573_, _32412_);
  and (_32586_, _32578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_33884_, _32586_, _32585_);
  and (_32595_, _32573_, _32415_);
  not (_32596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_32597_, _32573_, _32596_);
  or (_33887_, _32597_, _32595_);
  and (_32606_, _32573_, _32418_);
  and (_32607_, _32578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_33891_, _32607_, _32606_);
  and (_32612_, _32573_, _32421_);
  not (_32617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_32618_, _32573_, _32617_);
  or (_33894_, _32618_, _32612_);
  and (_32622_, _32573_, _32425_);
  not (_32628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_32629_, _32573_, _32628_);
  or (_33898_, _32629_, _32622_);
  and (_32630_, _32573_, _32429_);
  and (_32636_, _32578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_33901_, _32636_, _32630_);
  and (_32640_, _32573_, _32320_);
  not (_32641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_32646_, _32573_, _32641_);
  or (_33904_, _32646_, _32640_);
  and (_32651_, _32479_, _32306_);
  and (_32652_, _32651_, _32406_);
  not (_32657_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_32662_, _32651_, _32657_);
  or (_33908_, _32662_, _32652_);
  and (_32663_, _32651_, _32412_);
  not (_32667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_32673_, _32651_, _32667_);
  or (_33912_, _32673_, _32663_);
  and (_32674_, _32651_, _32415_);
  not (_32677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_32683_, _32651_, _32677_);
  or (_33915_, _32683_, _32674_);
  and (_32685_, _32651_, _32418_);
  not (_32687_, _32651_);
  and (_32693_, _32687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_33919_, _32693_, _32685_);
  and (_32696_, _32651_, _32421_);
  and (_32698_, _32687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_33922_, _32698_, _32696_);
  and (_32706_, _32651_, _32425_);
  and (_32707_, _32687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_33926_, _32707_, _32706_);
  and (_32714_, _32651_, _32429_);
  not (_32716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_32717_, _32651_, _32716_);
  or (_33929_, _32717_, _32714_);
  and (_32718_, _32651_, _32320_);
  nor (_32719_, _32651_, _32266_);
  or (_33932_, _32719_, _32718_);
  and (_32720_, _32307_, _32021_);
  and (_32721_, _32720_, _32325_);
  and (_32722_, _32721_, _32406_);
  not (_32723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_32724_, _32721_, _32723_);
  or (_33939_, _32724_, _32722_);
  and (_32725_, _32721_, _32412_);
  not (_32726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32727_, _32721_, _32726_);
  or (_33942_, _32727_, _32725_);
  and (_32728_, _32721_, _32415_);
  not (_32729_, _32721_);
  and (_32730_, _32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_33946_, _32730_, _32728_);
  and (_32731_, _32721_, _32418_);
  not (_32732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_32733_, _32721_, _32732_);
  or (_33949_, _32733_, _32731_);
  and (_32734_, _32721_, _32421_);
  and (_32735_, _32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_33953_, _32735_, _32734_);
  and (_32736_, _32721_, _32425_);
  and (_32737_, _32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_33956_, _32737_, _32736_);
  and (_32738_, _32721_, _32429_);
  and (_32739_, _32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_33960_, _32739_, _32738_);
  and (_32740_, _32721_, _32320_);
  and (_32741_, _32729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_33962_, _32741_, _32740_);
  and (_32742_, _32720_, _32407_);
  and (_32743_, _32742_, _32406_);
  not (_32744_, _32742_);
  and (_32745_, _32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_33967_, _32745_, _32743_);
  and (_32746_, _32742_, _32412_);
  and (_32747_, _32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_33970_, _32747_, _32746_);
  and (_32748_, _32742_, _32415_);
  and (_32749_, _32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_33974_, _32749_, _32748_);
  and (_32750_, _32742_, _32418_);
  and (_32751_, _32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_33977_, _32751_, _32750_);
  and (_32752_, _32742_, _32421_);
  not (_32753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_32754_, _32742_, _32753_);
  or (_33981_, _32754_, _32752_);
  and (_32755_, _32742_, _32425_);
  not (_32756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_32757_, _32742_, _32756_);
  or (_33984_, _32757_, _32755_);
  and (_32758_, _32742_, _32429_);
  not (_32759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_32760_, _32742_, _32759_);
  or (_33988_, _32760_, _32758_);
  and (_32761_, _32742_, _32320_);
  and (_32762_, _32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_33990_, _32762_, _32761_);
  and (_32763_, _32720_, _32434_);
  and (_32764_, _32763_, _32406_);
  not (_32765_, _32763_);
  and (_32766_, _32765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_33994_, _32766_, _32764_);
  and (_32767_, _32763_, _32412_);
  and (_32768_, _32765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_33997_, _32768_, _32767_);
  and (_32769_, _32763_, _32415_);
  not (_32770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_32771_, _32763_, _32770_);
  or (_34001_, _32771_, _32769_);
  and (_32772_, _32763_, _32418_);
  and (_32773_, _32765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_34005_, _32773_, _32772_);
  and (_32774_, _32763_, _32421_);
  not (_32775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_32776_, _32763_, _32775_);
  or (_34009_, _32776_, _32774_);
  and (_32777_, _32763_, _32425_);
  not (_32778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_32779_, _32763_, _32778_);
  or (_34013_, _32779_, _32777_);
  and (_32780_, _32763_, _32429_);
  not (_32781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_32782_, _32763_, _32781_);
  or (_34017_, _32782_, _32780_);
  and (_32783_, _32763_, _32320_);
  nor (_32784_, _32763_, _32280_);
  or (_34020_, _32784_, _32783_);
  and (_32785_, _32720_, _32306_);
  and (_32786_, _32785_, _32406_);
  not (_32787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_32788_, _32785_, _32787_);
  or (_34025_, _32788_, _32786_);
  and (_32789_, _32785_, _32412_);
  not (_32790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_32791_, _32785_, _32790_);
  or (_34029_, _32791_, _32789_);
  and (_32792_, _32785_, _32415_);
  not (_32793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_32794_, _32785_, _32793_);
  or (_34033_, _32794_, _32792_);
  and (_32795_, _32785_, _32418_);
  not (_32796_, _32785_);
  and (_32797_, _32796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_34037_, _32797_, _32795_);
  and (_32798_, _32785_, _32421_);
  and (_32799_, _32796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_34041_, _32799_, _32798_);
  and (_32800_, _32785_, _32425_);
  and (_32801_, _32796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_34045_, _32801_, _32800_);
  and (_32802_, _32785_, _32429_);
  and (_32803_, _32796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_34049_, _32803_, _32802_);
  and (_32804_, _32785_, _32320_);
  not (_32805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_32806_, _32785_, _32805_);
  or (_34052_, _32806_, _32804_);
  and (_32807_, _32325_, _32309_);
  and (_32808_, _32807_, _32406_);
  not (_32809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_32810_, _32807_, _32809_);
  or (_34058_, _32810_, _32808_);
  and (_32811_, _32807_, _32412_);
  not (_32812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_32813_, _32807_, _32812_);
  or (_34062_, _32813_, _32811_);
  and (_32814_, _32807_, _32415_);
  not (_32815_, _32807_);
  and (_32816_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_34066_, _32816_, _32814_);
  and (_32817_, _32807_, _32418_);
  and (_32818_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_34070_, _32818_, _32817_);
  and (_32819_, _32807_, _32421_);
  and (_32820_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_34074_, _32820_, _32819_);
  and (_32821_, _32807_, _32425_);
  and (_32822_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_34078_, _32822_, _32821_);
  and (_32823_, _32807_, _32429_);
  and (_32824_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_34082_, _32824_, _32823_);
  and (_32825_, _32807_, _32320_);
  and (_32826_, _32815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_34085_, _32826_, _32825_);
  and (_32827_, _32407_, _32309_);
  and (_32828_, _32827_, _32406_);
  not (_32829_, _32827_);
  and (_32830_, _32829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_34090_, _32830_, _32828_);
  and (_32831_, _32827_, _32412_);
  and (_32832_, _32829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_34094_, _32832_, _32831_);
  and (_32833_, _32827_, _32415_);
  and (_32834_, _32829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_34098_, _32834_, _32833_);
  and (_32835_, _32827_, _32418_);
  and (_32836_, _32829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_34102_, _32836_, _32835_);
  and (_32837_, _32827_, _32421_);
  not (_32838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_32839_, _32827_, _32838_);
  or (_34106_, _32839_, _32837_);
  and (_32840_, _32827_, _32425_);
  not (_32841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_32842_, _32827_, _32841_);
  or (_34109_, _32842_, _32840_);
  and (_32843_, _32827_, _32429_);
  not (_32844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_32845_, _32827_, _32844_);
  or (_34113_, _32845_, _32843_);
  and (_32846_, _32827_, _32320_);
  and (_32847_, _32829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_34115_, _32847_, _32846_);
  and (_32848_, _32434_, _32309_);
  and (_32849_, _32848_, _32406_);
  not (_32850_, _32848_);
  and (_32851_, _32850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_34120_, _32851_, _32849_);
  and (_32852_, _32848_, _32412_);
  and (_32853_, _32850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_34124_, _32853_, _32852_);
  and (_32854_, _32848_, _32415_);
  not (_32855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_32856_, _32848_, _32855_);
  or (_34128_, _32856_, _32854_);
  and (_32857_, _32848_, _32418_);
  not (_32858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_32859_, _32848_, _32858_);
  or (_34132_, _32859_, _32857_);
  and (_32860_, _32848_, _32421_);
  not (_32861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_32862_, _32848_, _32861_);
  or (_34136_, _32862_, _32860_);
  and (_32863_, _32848_, _32425_);
  not (_32864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_32865_, _32848_, _32864_);
  or (_34139_, _32865_, _32863_);
  and (_32866_, _32848_, _32429_);
  not (_32867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_32868_, _32848_, _32867_);
  or (_34143_, _32868_, _32866_);
  and (_32869_, _32848_, _32320_);
  nor (_32870_, _32848_, _32291_);
  or (_34146_, _32870_, _32869_);
  and (_32871_, _32406_, _32310_);
  not (_32872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_32873_, _32310_, _32872_);
  or (_34151_, _32873_, _32871_);
  and (_32874_, _32412_, _32310_);
  not (_32875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_32876_, _32310_, _32875_);
  or (_34155_, _32876_, _32874_);
  and (_32877_, _32415_, _32310_);
  not (_32878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_32879_, _32310_, _32878_);
  or (_34159_, _32879_, _32877_);
  and (_32880_, _32418_, _32310_);
  not (_32881_, _32310_);
  and (_32882_, _32881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_34162_, _32882_, _32880_);
  and (_32883_, _32421_, _32310_);
  and (_32884_, _32881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_34166_, _32884_, _32883_);
  and (_32885_, _32425_, _32310_);
  and (_32886_, _32881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_34170_, _32886_, _32885_);
  and (_32887_, _32429_, _32310_);
  and (_32888_, _32881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_34174_, _32888_, _32887_);
  or (_32889_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_32890_, _32098_, _32339_);
  and (_32891_, _32890_, _32233_);
  and (_32892_, _32891_, _32889_);
  nor (_32893_, _32098_, _32459_);
  and (_32894_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_32895_, _32894_, _32893_);
  and (_32896_, _32895_, _32253_);
  or (_32897_, _32896_, _32892_);
  or (_32898_, _32897_, _32247_);
  or (_32899_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_32900_, _32098_, _32482_);
  and (_32901_, _32900_, _32233_);
  and (_32902_, _32901_, _32899_);
  nor (_32903_, _32098_, _32657_);
  and (_32904_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_32905_, _32904_, _32903_);
  and (_32906_, _32905_, _32253_);
  or (_32907_, _32906_, _32902_);
  or (_32908_, _32907_, _32017_);
  and (_32909_, _32908_, _32261_);
  and (_32910_, _32909_, _32898_);
  nand (_32911_, _32098_, _32723_);
  or (_32912_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_32913_, _32912_, _32911_);
  and (_32914_, _32913_, _32233_);
  and (_32915_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_32916_, _32098_, _32787_);
  or (_32917_, _32916_, _32915_);
  and (_32918_, _32917_, _32253_);
  or (_32919_, _32918_, _32914_);
  or (_32920_, _32919_, _32247_);
  nand (_32921_, _32098_, _32809_);
  or (_32922_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_32923_, _32922_, _32921_);
  and (_32924_, _32923_, _32233_);
  and (_32925_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_32926_, _32098_, _32872_);
  or (_32927_, _32926_, _32925_);
  and (_32928_, _32927_, _32253_);
  or (_32929_, _32928_, _32924_);
  or (_32930_, _32929_, _32017_);
  and (_32931_, _32930_, _32144_);
  and (_32932_, _32931_, _32920_);
  or (_32933_, _32932_, _32910_);
  or (_32934_, _32933_, _32246_);
  or (_32935_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_32936_, _32935_, _36029_);
  and (_36008_, _32936_, _32934_);
  or (_32937_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_32938_, _32098_, _32352_);
  and (_32939_, _32938_, _32233_);
  and (_32940_, _32939_, _32937_);
  nor (_32941_, _32098_, _32462_);
  and (_32942_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_32943_, _32942_, _32941_);
  and (_32944_, _32943_, _32253_);
  or (_32945_, _32944_, _32940_);
  or (_32946_, _32945_, _32247_);
  or (_32947_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_32948_, _32098_, _32502_);
  and (_32949_, _32948_, _32233_);
  and (_32950_, _32949_, _32947_);
  nor (_32951_, _32098_, _32667_);
  and (_32952_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_32953_, _32952_, _32951_);
  and (_32954_, _32953_, _32253_);
  or (_32955_, _32954_, _32950_);
  or (_32956_, _32955_, _32017_);
  and (_32957_, _32956_, _32261_);
  and (_32958_, _32957_, _32946_);
  nand (_32959_, _32098_, _32726_);
  or (_32960_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_32961_, _32960_, _32959_);
  and (_32962_, _32961_, _32233_);
  and (_32963_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_32964_, _32098_, _32790_);
  or (_32965_, _32964_, _32963_);
  and (_32966_, _32965_, _32253_);
  or (_32967_, _32966_, _32962_);
  or (_32968_, _32967_, _32247_);
  nand (_32969_, _32098_, _32812_);
  or (_32970_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_32971_, _32970_, _32969_);
  and (_32972_, _32971_, _32233_);
  and (_32973_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_32974_, _32098_, _32875_);
  or (_32975_, _32974_, _32973_);
  and (_32976_, _32975_, _32253_);
  or (_32977_, _32976_, _32972_);
  or (_32978_, _32977_, _32017_);
  and (_32979_, _32978_, _32144_);
  and (_32980_, _32979_, _32968_);
  or (_32981_, _32980_, _32958_);
  or (_32982_, _32981_, _32246_);
  or (_32983_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_32984_, _32983_, _36029_);
  and (_36010_, _32984_, _32982_);
  and (_32985_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_32986_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_32987_, _32986_, _32985_);
  and (_32988_, _32987_, _32233_);
  nor (_32989_, _32098_, _32465_);
  and (_32990_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_32991_, _32990_, _32989_);
  and (_32992_, _32991_, _32253_);
  or (_32993_, _32992_, _32988_);
  or (_32994_, _32993_, _32247_);
  and (_32995_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_32996_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_32997_, _32996_, _32995_);
  and (_32998_, _32997_, _32233_);
  nor (_32999_, _32098_, _32677_);
  and (_33000_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_33001_, _33000_, _32999_);
  and (_33002_, _33001_, _32253_);
  or (_33003_, _33002_, _32998_);
  or (_33004_, _33003_, _32017_);
  and (_33005_, _33004_, _32261_);
  and (_33006_, _33005_, _32994_);
  or (_33007_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_33008_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_33009_, _33008_, _33007_);
  and (_33010_, _33009_, _32233_);
  or (_33011_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_33012_, _32098_, _32770_);
  and (_33013_, _33012_, _33011_);
  and (_33014_, _33013_, _32253_);
  or (_33015_, _33014_, _33010_);
  or (_33016_, _33015_, _32247_);
  or (_33017_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_33018_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_33019_, _33018_, _33017_);
  and (_33020_, _33019_, _32233_);
  or (_33021_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_33022_, _32098_, _32855_);
  and (_33023_, _33022_, _33021_);
  and (_33024_, _33023_, _32253_);
  or (_33025_, _33024_, _33020_);
  or (_33026_, _33025_, _32017_);
  and (_33027_, _33026_, _32144_);
  and (_33028_, _33027_, _33016_);
  or (_33029_, _33028_, _33006_);
  or (_33030_, _33029_, _32246_);
  or (_33031_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_33032_, _33031_, _36029_);
  and (_36012_, _33032_, _33030_);
  or (_33033_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_33034_, _32098_, _32858_);
  and (_33035_, _33034_, _33033_);
  or (_33036_, _33035_, _32233_);
  or (_33037_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_33038_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_33039_, _33038_, _33037_);
  or (_33040_, _33039_, _32253_);
  and (_33041_, _33040_, _32144_);
  and (_33042_, _33041_, _33036_);
  and (_33043_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_33044_, _32098_, _32536_);
  or (_33045_, _33044_, _32253_);
  or (_33046_, _33045_, _33043_);
  and (_33047_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_33048_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_33049_, _33048_, _32233_);
  or (_33050_, _33049_, _33047_);
  and (_33051_, _33050_, _32261_);
  and (_33052_, _33051_, _33046_);
  or (_33053_, _33052_, _33042_);
  and (_33054_, _33053_, _32247_);
  or (_33055_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_33056_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_33057_, _33056_, _33055_);
  or (_33058_, _33057_, _32233_);
  nand (_33059_, _32098_, _32732_);
  or (_33060_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_33061_, _33060_, _33059_);
  or (_33062_, _33061_, _32253_);
  and (_33063_, _33062_, _32144_);
  and (_33064_, _33063_, _33058_);
  and (_33065_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_33066_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_33067_, _33066_, _32253_);
  or (_33068_, _33067_, _33065_);
  nor (_33069_, _32098_, _32468_);
  and (_33070_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_33071_, _33070_, _32233_);
  or (_33072_, _33071_, _33069_);
  and (_33073_, _33072_, _32261_);
  and (_33074_, _33073_, _33068_);
  or (_33075_, _33074_, _33064_);
  and (_33076_, _33075_, _32017_);
  or (_33077_, _33076_, _32246_);
  or (_33078_, _33077_, _33054_);
  or (_33079_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_33080_, _33079_, _36029_);
  and (_36013_, _33080_, _33078_);
  and (_33081_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_33082_, _32098_, _32423_);
  or (_33083_, _33082_, _33081_);
  and (_33084_, _33083_, _32233_);
  or (_33085_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_33086_, _32098_, _32447_);
  and (_33087_, _33086_, _33085_);
  and (_33088_, _33087_, _32253_);
  or (_33089_, _33088_, _33084_);
  or (_33090_, _33089_, _32247_);
  and (_33091_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_33092_, _32098_, _32539_);
  or (_33093_, _33092_, _33091_);
  and (_33094_, _33093_, _32233_);
  or (_33095_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_33096_, _32098_, _32617_);
  and (_33097_, _33096_, _33095_);
  and (_33098_, _33097_, _32253_);
  or (_33099_, _33098_, _33094_);
  or (_33100_, _33099_, _32017_);
  and (_33101_, _33100_, _32261_);
  and (_33102_, _33101_, _33090_);
  and (_33103_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_33104_, _32098_, _32753_);
  or (_33105_, _33104_, _33103_);
  and (_33106_, _33105_, _32233_);
  or (_33107_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_33108_, _32098_, _32775_);
  and (_33109_, _33108_, _33107_);
  and (_33110_, _33109_, _32253_);
  or (_33111_, _33110_, _33106_);
  or (_33112_, _33111_, _32247_);
  and (_33113_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_33114_, _32098_, _32838_);
  or (_33115_, _33114_, _33113_);
  and (_33116_, _33115_, _32233_);
  or (_33117_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_33118_, _32098_, _32861_);
  and (_33119_, _33118_, _33117_);
  and (_33120_, _33119_, _32253_);
  or (_33121_, _33120_, _33116_);
  or (_33122_, _33121_, _32017_);
  and (_33123_, _33122_, _32144_);
  and (_33124_, _33123_, _33112_);
  or (_33125_, _33124_, _33102_);
  or (_33126_, _33125_, _32246_);
  or (_33127_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_33128_, _33127_, _36029_);
  and (_36015_, _33128_, _33126_);
  and (_33129_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_33130_, _32098_, _32427_);
  or (_33131_, _33130_, _33129_);
  and (_33132_, _33131_, _32233_);
  or (_33133_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_33134_, _32098_, _32450_);
  and (_33135_, _33134_, _33133_);
  and (_33136_, _33135_, _32253_);
  or (_33137_, _33136_, _33132_);
  or (_33138_, _33137_, _32247_);
  and (_33139_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_33140_, _32098_, _32550_);
  or (_33141_, _33140_, _33139_);
  and (_33142_, _33141_, _32233_);
  or (_33143_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_33144_, _32098_, _32628_);
  and (_33145_, _33144_, _33143_);
  and (_33146_, _33145_, _32253_);
  or (_33147_, _33146_, _33142_);
  or (_33148_, _33147_, _32017_);
  and (_33149_, _33148_, _32261_);
  and (_33150_, _33149_, _33138_);
  and (_33151_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_33152_, _32098_, _32756_);
  or (_33153_, _33152_, _33151_);
  and (_33154_, _33153_, _32233_);
  or (_33155_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_33156_, _32098_, _32778_);
  and (_33157_, _33156_, _33155_);
  and (_33158_, _33157_, _32253_);
  or (_33159_, _33158_, _33154_);
  or (_33160_, _33159_, _32247_);
  and (_33161_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_33162_, _32098_, _32841_);
  or (_33163_, _33162_, _33161_);
  and (_33164_, _33163_, _32233_);
  or (_33165_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_33166_, _32098_, _32864_);
  and (_33167_, _33166_, _33165_);
  and (_33168_, _33167_, _32253_);
  or (_33169_, _33168_, _33164_);
  or (_33170_, _33169_, _32017_);
  and (_33171_, _33170_, _32144_);
  and (_33172_, _33171_, _33160_);
  or (_33173_, _33172_, _33150_);
  or (_33174_, _33173_, _32246_);
  or (_33175_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_33176_, _33175_, _36029_);
  and (_36017_, _33176_, _33174_);
  and (_33177_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_33178_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_33179_, _33178_, _33177_);
  and (_33180_, _33179_, _32233_);
  and (_33181_, _32249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_33182_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_33183_, _33182_, _33181_);
  and (_33184_, _33183_, _32253_);
  or (_33185_, _33184_, _33180_);
  or (_33186_, _33185_, _32247_);
  and (_33187_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_33188_, _32098_, _32561_);
  or (_33189_, _33188_, _33187_);
  and (_33190_, _33189_, _32233_);
  nor (_33191_, _32098_, _32716_);
  and (_33192_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_33193_, _33192_, _33191_);
  and (_33194_, _33193_, _32253_);
  or (_33195_, _33194_, _33190_);
  or (_33196_, _33195_, _32017_);
  and (_33197_, _33196_, _32261_);
  and (_33198_, _33197_, _33186_);
  and (_33199_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_33200_, _32098_, _32759_);
  or (_33201_, _33200_, _33199_);
  and (_33202_, _33201_, _32233_);
  or (_33203_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_33204_, _32098_, _32781_);
  and (_33205_, _33204_, _33203_);
  and (_33206_, _33205_, _32253_);
  or (_33207_, _33206_, _33202_);
  or (_33208_, _33207_, _32247_);
  and (_33209_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_33210_, _32098_, _32844_);
  or (_33211_, _33210_, _33209_);
  and (_33212_, _33211_, _32233_);
  or (_33213_, _32098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_33214_, _32098_, _32867_);
  and (_33215_, _33214_, _33213_);
  and (_33216_, _33215_, _32253_);
  or (_33217_, _33216_, _33212_);
  or (_33218_, _33217_, _32017_);
  and (_33219_, _33218_, _32144_);
  and (_33220_, _33219_, _33208_);
  or (_33221_, _33220_, _33198_);
  or (_33222_, _33221_, _32246_);
  or (_33223_, _32301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_33224_, _33223_, _36029_);
  and (_36019_, _33224_, _33222_);
  or (_33225_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_33226_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_33227_, _33226_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_33228_, _33227_, _33225_);
  nand (_33229_, _33228_, _36029_);
  or (_33230_, \oc8051_gm_cxrom_1.cell0.data [7], _36029_);
  and (_36026_, _33230_, _33229_);
  or (_33231_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33232_, \oc8051_gm_cxrom_1.cell0.data [0], _33226_);
  nand (_33233_, _33232_, _33231_);
  nand (_33234_, _33233_, _36029_);
  or (_33235_, \oc8051_gm_cxrom_1.cell0.data [0], _36029_);
  and (_36033_, _33235_, _33234_);
  or (_33236_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33237_, \oc8051_gm_cxrom_1.cell0.data [1], _33226_);
  nand (_33238_, _33237_, _33236_);
  nand (_33239_, _33238_, _36029_);
  or (_33240_, \oc8051_gm_cxrom_1.cell0.data [1], _36029_);
  and (_36036_, _33240_, _33239_);
  or (_33241_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33242_, \oc8051_gm_cxrom_1.cell0.data [2], _33226_);
  nand (_33243_, _33242_, _33241_);
  nand (_33244_, _33243_, _36029_);
  or (_33245_, \oc8051_gm_cxrom_1.cell0.data [2], _36029_);
  and (_36040_, _33245_, _33244_);
  or (_33246_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33247_, \oc8051_gm_cxrom_1.cell0.data [3], _33226_);
  nand (_33248_, _33247_, _33246_);
  nand (_33249_, _33248_, _36029_);
  or (_33250_, \oc8051_gm_cxrom_1.cell0.data [3], _36029_);
  and (_36043_, _33250_, _33249_);
  or (_33251_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33252_, \oc8051_gm_cxrom_1.cell0.data [4], _33226_);
  nand (_33253_, _33252_, _33251_);
  nand (_33254_, _33253_, _36029_);
  or (_33255_, \oc8051_gm_cxrom_1.cell0.data [4], _36029_);
  and (_36047_, _33255_, _33254_);
  or (_33256_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33257_, \oc8051_gm_cxrom_1.cell0.data [5], _33226_);
  nand (_33258_, _33257_, _33256_);
  nand (_33259_, _33258_, _36029_);
  or (_33260_, \oc8051_gm_cxrom_1.cell0.data [5], _36029_);
  and (_36051_, _33260_, _33259_);
  or (_33261_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33262_, \oc8051_gm_cxrom_1.cell0.data [6], _33226_);
  nand (_33263_, _33262_, _33261_);
  nand (_33264_, _33263_, _36029_);
  or (_33265_, \oc8051_gm_cxrom_1.cell0.data [6], _36029_);
  and (_36054_, _33265_, _33264_);
  or (_33266_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_33267_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_33268_, _33267_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_33269_, _33268_, _33266_);
  nand (_33270_, _33269_, _36029_);
  or (_33271_, \oc8051_gm_cxrom_1.cell1.data [7], _36029_);
  and (_36074_, _33271_, _33270_);
  or (_33272_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33273_, \oc8051_gm_cxrom_1.cell1.data [0], _33267_);
  nand (_33274_, _33273_, _33272_);
  nand (_33275_, _33274_, _36029_);
  or (_33276_, \oc8051_gm_cxrom_1.cell1.data [0], _36029_);
  and (_36080_, _33276_, _33275_);
  or (_33277_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33278_, \oc8051_gm_cxrom_1.cell1.data [1], _33267_);
  nand (_33279_, _33278_, _33277_);
  nand (_33280_, _33279_, _36029_);
  or (_33281_, \oc8051_gm_cxrom_1.cell1.data [1], _36029_);
  and (_36084_, _33281_, _33280_);
  or (_33282_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33283_, \oc8051_gm_cxrom_1.cell1.data [2], _33267_);
  nand (_33284_, _33283_, _33282_);
  nand (_33285_, _33284_, _36029_);
  or (_33286_, \oc8051_gm_cxrom_1.cell1.data [2], _36029_);
  and (_36087_, _33286_, _33285_);
  or (_33287_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33288_, \oc8051_gm_cxrom_1.cell1.data [3], _33267_);
  nand (_33289_, _33288_, _33287_);
  nand (_33290_, _33289_, _36029_);
  or (_33291_, \oc8051_gm_cxrom_1.cell1.data [3], _36029_);
  and (_36091_, _33291_, _33290_);
  or (_33292_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33293_, \oc8051_gm_cxrom_1.cell1.data [4], _33267_);
  nand (_33294_, _33293_, _33292_);
  nand (_33295_, _33294_, _36029_);
  or (_33296_, \oc8051_gm_cxrom_1.cell1.data [4], _36029_);
  and (_36095_, _33296_, _33295_);
  or (_33297_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33298_, \oc8051_gm_cxrom_1.cell1.data [5], _33267_);
  nand (_33299_, _33298_, _33297_);
  nand (_33300_, _33299_, _36029_);
  or (_33301_, \oc8051_gm_cxrom_1.cell1.data [5], _36029_);
  and (_36098_, _33301_, _33300_);
  or (_33302_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33303_, \oc8051_gm_cxrom_1.cell1.data [6], _33267_);
  nand (_33304_, _33303_, _33302_);
  nand (_33305_, _33304_, _36029_);
  or (_33306_, \oc8051_gm_cxrom_1.cell1.data [6], _36029_);
  and (_36102_, _33306_, _33305_);
  or (_33307_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_33308_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_33309_, _33308_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_33310_, _33309_, _33307_);
  nand (_33311_, _33310_, _36029_);
  or (_33312_, \oc8051_gm_cxrom_1.cell2.data [7], _36029_);
  and (_36115_, _33312_, _33311_);
  or (_33313_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33314_, \oc8051_gm_cxrom_1.cell2.data [0], _33308_);
  nand (_33316_, _33314_, _33313_);
  nand (_33318_, _33316_, _36029_);
  or (_33320_, \oc8051_gm_cxrom_1.cell2.data [0], _36029_);
  and (_36121_, _33320_, _33318_);
  or (_33323_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33325_, \oc8051_gm_cxrom_1.cell2.data [1], _33308_);
  nand (_33327_, _33325_, _33323_);
  nand (_33329_, _33327_, _36029_);
  or (_33331_, \oc8051_gm_cxrom_1.cell2.data [1], _36029_);
  and (_36125_, _33331_, _33329_);
  or (_33334_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33336_, \oc8051_gm_cxrom_1.cell2.data [2], _33308_);
  nand (_33338_, _33336_, _33334_);
  nand (_33340_, _33338_, _36029_);
  or (_33342_, \oc8051_gm_cxrom_1.cell2.data [2], _36029_);
  and (_36128_, _33342_, _33340_);
  or (_33345_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33347_, \oc8051_gm_cxrom_1.cell2.data [3], _33308_);
  nand (_33349_, _33347_, _33345_);
  nand (_33351_, _33349_, _36029_);
  or (_33353_, \oc8051_gm_cxrom_1.cell2.data [3], _36029_);
  and (_00009_, _33353_, _33351_);
  or (_33356_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33358_, \oc8051_gm_cxrom_1.cell2.data [4], _33308_);
  nand (_33360_, _33358_, _33356_);
  nand (_33362_, _33360_, _36029_);
  or (_33364_, \oc8051_gm_cxrom_1.cell2.data [4], _36029_);
  and (_00012_, _33364_, _33362_);
  or (_33366_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33367_, \oc8051_gm_cxrom_1.cell2.data [5], _33308_);
  nand (_33368_, _33367_, _33366_);
  nand (_33369_, _33368_, _36029_);
  or (_33370_, \oc8051_gm_cxrom_1.cell2.data [5], _36029_);
  and (_00016_, _33370_, _33369_);
  or (_33371_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33372_, \oc8051_gm_cxrom_1.cell2.data [6], _33308_);
  nand (_33373_, _33372_, _33371_);
  nand (_33374_, _33373_, _36029_);
  or (_33375_, \oc8051_gm_cxrom_1.cell2.data [6], _36029_);
  and (_00019_, _33375_, _33374_);
  or (_33376_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_33377_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_33378_, _33377_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_33379_, _33378_, _33376_);
  nand (_33380_, _33379_, _36029_);
  or (_33381_, \oc8051_gm_cxrom_1.cell3.data [7], _36029_);
  and (_00033_, _33381_, _33380_);
  or (_33382_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33383_, \oc8051_gm_cxrom_1.cell3.data [0], _33377_);
  nand (_33384_, _33383_, _33382_);
  nand (_33385_, _33384_, _36029_);
  or (_33386_, \oc8051_gm_cxrom_1.cell3.data [0], _36029_);
  and (_00039_, _33386_, _33385_);
  or (_33387_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33388_, \oc8051_gm_cxrom_1.cell3.data [1], _33377_);
  nand (_33389_, _33388_, _33387_);
  nand (_33390_, _33389_, _36029_);
  or (_33391_, \oc8051_gm_cxrom_1.cell3.data [1], _36029_);
  and (_00042_, _33391_, _33390_);
  or (_33392_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33393_, \oc8051_gm_cxrom_1.cell3.data [2], _33377_);
  nand (_33394_, _33393_, _33392_);
  nand (_33395_, _33394_, _36029_);
  or (_33396_, \oc8051_gm_cxrom_1.cell3.data [2], _36029_);
  and (_00045_, _33396_, _33395_);
  or (_33397_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33398_, \oc8051_gm_cxrom_1.cell3.data [3], _33377_);
  nand (_33399_, _33398_, _33397_);
  nand (_33400_, _33399_, _36029_);
  or (_33401_, \oc8051_gm_cxrom_1.cell3.data [3], _36029_);
  and (_00049_, _33401_, _33400_);
  or (_33402_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33403_, \oc8051_gm_cxrom_1.cell3.data [4], _33377_);
  nand (_33404_, _33403_, _33402_);
  nand (_33405_, _33404_, _36029_);
  or (_33406_, \oc8051_gm_cxrom_1.cell3.data [4], _36029_);
  and (_00052_, _33406_, _33405_);
  or (_33407_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33408_, \oc8051_gm_cxrom_1.cell3.data [5], _33377_);
  nand (_33409_, _33408_, _33407_);
  nand (_33410_, _33409_, _36029_);
  or (_33411_, \oc8051_gm_cxrom_1.cell3.data [5], _36029_);
  and (_00055_, _33411_, _33410_);
  or (_33412_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33413_, \oc8051_gm_cxrom_1.cell3.data [6], _33377_);
  nand (_33414_, _33413_, _33412_);
  nand (_33415_, _33414_, _36029_);
  or (_33416_, \oc8051_gm_cxrom_1.cell3.data [6], _36029_);
  and (_00058_, _33416_, _33415_);
  or (_33417_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_33418_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_33419_, _33418_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_33420_, _33419_, _33417_);
  nand (_33421_, _33420_, _36029_);
  or (_33422_, \oc8051_gm_cxrom_1.cell4.data [7], _36029_);
  and (_00075_, _33422_, _33421_);
  or (_33423_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33424_, \oc8051_gm_cxrom_1.cell4.data [0], _33418_);
  nand (_33425_, _33424_, _33423_);
  nand (_33426_, _33425_, _36029_);
  or (_33427_, \oc8051_gm_cxrom_1.cell4.data [0], _36029_);
  and (_00081_, _33427_, _33426_);
  or (_33428_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33429_, \oc8051_gm_cxrom_1.cell4.data [1], _33418_);
  nand (_33430_, _33429_, _33428_);
  nand (_33431_, _33430_, _36029_);
  or (_33432_, \oc8051_gm_cxrom_1.cell4.data [1], _36029_);
  and (_00084_, _33432_, _33431_);
  or (_33433_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33434_, \oc8051_gm_cxrom_1.cell4.data [2], _33418_);
  nand (_33435_, _33434_, _33433_);
  nand (_33436_, _33435_, _36029_);
  or (_33437_, \oc8051_gm_cxrom_1.cell4.data [2], _36029_);
  and (_00087_, _33437_, _33436_);
  or (_33438_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33439_, \oc8051_gm_cxrom_1.cell4.data [3], _33418_);
  nand (_33441_, _33439_, _33438_);
  nand (_33442_, _33441_, _36029_);
  or (_33443_, \oc8051_gm_cxrom_1.cell4.data [3], _36029_);
  and (_00091_, _33443_, _33442_);
  or (_33444_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33445_, \oc8051_gm_cxrom_1.cell4.data [4], _33418_);
  nand (_33446_, _33445_, _33444_);
  nand (_33447_, _33446_, _36029_);
  or (_33448_, \oc8051_gm_cxrom_1.cell4.data [4], _36029_);
  and (_00094_, _33448_, _33447_);
  or (_33449_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33451_, \oc8051_gm_cxrom_1.cell4.data [5], _33418_);
  nand (_33452_, _33451_, _33449_);
  nand (_33453_, _33452_, _36029_);
  or (_33454_, \oc8051_gm_cxrom_1.cell4.data [5], _36029_);
  and (_00097_, _33454_, _33453_);
  or (_33455_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33456_, \oc8051_gm_cxrom_1.cell4.data [6], _33418_);
  nand (_33457_, _33456_, _33455_);
  nand (_33458_, _33457_, _36029_);
  or (_33459_, \oc8051_gm_cxrom_1.cell4.data [6], _36029_);
  and (_00100_, _33459_, _33458_);
  or (_33460_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_33461_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_33462_, _33461_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_33463_, _33462_, _33460_);
  nand (_33464_, _33463_, _36029_);
  or (_33465_, \oc8051_gm_cxrom_1.cell5.data [7], _36029_);
  and (_00117_, _33465_, _33464_);
  or (_33466_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33467_, \oc8051_gm_cxrom_1.cell5.data [0], _33461_);
  nand (_33468_, _33467_, _33466_);
  nand (_33469_, _33468_, _36029_);
  or (_33470_, \oc8051_gm_cxrom_1.cell5.data [0], _36029_);
  and (_00123_, _33470_, _33469_);
  or (_33471_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33472_, \oc8051_gm_cxrom_1.cell5.data [1], _33461_);
  nand (_33473_, _33472_, _33471_);
  nand (_33474_, _33473_, _36029_);
  or (_33475_, \oc8051_gm_cxrom_1.cell5.data [1], _36029_);
  and (_00126_, _33475_, _33474_);
  or (_33476_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33477_, \oc8051_gm_cxrom_1.cell5.data [2], _33461_);
  nand (_33478_, _33477_, _33476_);
  nand (_33479_, _33478_, _36029_);
  or (_33480_, \oc8051_gm_cxrom_1.cell5.data [2], _36029_);
  and (_00129_, _33480_, _33479_);
  or (_33481_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33482_, \oc8051_gm_cxrom_1.cell5.data [3], _33461_);
  nand (_33483_, _33482_, _33481_);
  nand (_33484_, _33483_, _36029_);
  or (_33485_, \oc8051_gm_cxrom_1.cell5.data [3], _36029_);
  and (_00133_, _33485_, _33484_);
  or (_33486_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33487_, \oc8051_gm_cxrom_1.cell5.data [4], _33461_);
  nand (_33488_, _33487_, _33486_);
  nand (_33489_, _33488_, _36029_);
  or (_33490_, \oc8051_gm_cxrom_1.cell5.data [4], _36029_);
  and (_00136_, _33490_, _33489_);
  or (_33491_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33492_, \oc8051_gm_cxrom_1.cell5.data [5], _33461_);
  nand (_33493_, _33492_, _33491_);
  nand (_33494_, _33493_, _36029_);
  or (_33495_, \oc8051_gm_cxrom_1.cell5.data [5], _36029_);
  and (_00139_, _33495_, _33494_);
  or (_33496_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33497_, \oc8051_gm_cxrom_1.cell5.data [6], _33461_);
  nand (_33498_, _33497_, _33496_);
  nand (_33499_, _33498_, _36029_);
  or (_33500_, \oc8051_gm_cxrom_1.cell5.data [6], _36029_);
  and (_00142_, _33500_, _33499_);
  or (_33501_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_33502_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_33503_, _33502_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_33504_, _33503_, _33501_);
  nand (_33505_, _33504_, _36029_);
  or (_33506_, \oc8051_gm_cxrom_1.cell6.data [7], _36029_);
  and (_00159_, _33506_, _33505_);
  or (_33507_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33508_, \oc8051_gm_cxrom_1.cell6.data [0], _33502_);
  nand (_33509_, _33508_, _33507_);
  nand (_33510_, _33509_, _36029_);
  or (_33511_, \oc8051_gm_cxrom_1.cell6.data [0], _36029_);
  and (_00165_, _33511_, _33510_);
  or (_33512_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33513_, \oc8051_gm_cxrom_1.cell6.data [1], _33502_);
  nand (_33514_, _33513_, _33512_);
  nand (_33515_, _33514_, _36029_);
  or (_33516_, \oc8051_gm_cxrom_1.cell6.data [1], _36029_);
  and (_00168_, _33516_, _33515_);
  or (_33517_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33518_, \oc8051_gm_cxrom_1.cell6.data [2], _33502_);
  nand (_33519_, _33518_, _33517_);
  nand (_33520_, _33519_, _36029_);
  or (_33521_, \oc8051_gm_cxrom_1.cell6.data [2], _36029_);
  and (_00171_, _33521_, _33520_);
  or (_33522_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33523_, \oc8051_gm_cxrom_1.cell6.data [3], _33502_);
  nand (_33524_, _33523_, _33522_);
  nand (_33525_, _33524_, _36029_);
  or (_33526_, \oc8051_gm_cxrom_1.cell6.data [3], _36029_);
  and (_00175_, _33526_, _33525_);
  or (_33527_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33528_, \oc8051_gm_cxrom_1.cell6.data [4], _33502_);
  nand (_33529_, _33528_, _33527_);
  nand (_33530_, _33529_, _36029_);
  or (_33531_, \oc8051_gm_cxrom_1.cell6.data [4], _36029_);
  and (_00178_, _33531_, _33530_);
  or (_33532_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33533_, \oc8051_gm_cxrom_1.cell6.data [5], _33502_);
  nand (_33534_, _33533_, _33532_);
  nand (_33535_, _33534_, _36029_);
  or (_33536_, \oc8051_gm_cxrom_1.cell6.data [5], _36029_);
  and (_00182_, _33536_, _33535_);
  or (_33537_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33538_, \oc8051_gm_cxrom_1.cell6.data [6], _33502_);
  nand (_33539_, _33538_, _33537_);
  nand (_33540_, _33539_, _36029_);
  or (_33541_, \oc8051_gm_cxrom_1.cell6.data [6], _36029_);
  and (_00185_, _33541_, _33540_);
  or (_33542_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_33543_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_33544_, _33543_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_33545_, _33544_, _33542_);
  nand (_33546_, _33545_, _36029_);
  or (_33547_, \oc8051_gm_cxrom_1.cell7.data [7], _36029_);
  and (_00204_, _33547_, _33546_);
  or (_33548_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33549_, \oc8051_gm_cxrom_1.cell7.data [0], _33543_);
  nand (_33550_, _33549_, _33548_);
  nand (_33551_, _33550_, _36029_);
  or (_33552_, \oc8051_gm_cxrom_1.cell7.data [0], _36029_);
  and (_00211_, _33552_, _33551_);
  or (_33553_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33554_, \oc8051_gm_cxrom_1.cell7.data [1], _33543_);
  nand (_33555_, _33554_, _33553_);
  nand (_33556_, _33555_, _36029_);
  or (_33557_, \oc8051_gm_cxrom_1.cell7.data [1], _36029_);
  and (_00214_, _33557_, _33556_);
  or (_33558_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33559_, \oc8051_gm_cxrom_1.cell7.data [2], _33543_);
  nand (_33560_, _33559_, _33558_);
  nand (_33561_, _33560_, _36029_);
  or (_33562_, \oc8051_gm_cxrom_1.cell7.data [2], _36029_);
  and (_00218_, _33562_, _33561_);
  or (_33563_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33564_, \oc8051_gm_cxrom_1.cell7.data [3], _33543_);
  nand (_33565_, _33564_, _33563_);
  nand (_33566_, _33565_, _36029_);
  or (_33567_, \oc8051_gm_cxrom_1.cell7.data [3], _36029_);
  and (_00221_, _33567_, _33566_);
  or (_33568_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33569_, \oc8051_gm_cxrom_1.cell7.data [4], _33543_);
  nand (_33570_, _33569_, _33568_);
  nand (_33571_, _33570_, _36029_);
  or (_33572_, \oc8051_gm_cxrom_1.cell7.data [4], _36029_);
  and (_00225_, _33572_, _33571_);
  or (_33573_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33574_, \oc8051_gm_cxrom_1.cell7.data [5], _33543_);
  nand (_33575_, _33574_, _33573_);
  nand (_33576_, _33575_, _36029_);
  or (_33577_, \oc8051_gm_cxrom_1.cell7.data [5], _36029_);
  and (_00228_, _33577_, _33576_);
  or (_33578_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33579_, \oc8051_gm_cxrom_1.cell7.data [6], _33543_);
  nand (_33580_, _33579_, _33578_);
  nand (_33581_, _33580_, _36029_);
  or (_33582_, \oc8051_gm_cxrom_1.cell7.data [6], _36029_);
  and (_00232_, _33582_, _33581_);
  or (_33583_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_33584_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_33585_, _33584_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_33586_, _33585_, _33583_);
  nand (_33587_, _33586_, _36029_);
  or (_33588_, \oc8051_gm_cxrom_1.cell8.data [7], _36029_);
  and (_00250_, _33588_, _33587_);
  or (_33589_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33590_, \oc8051_gm_cxrom_1.cell8.data [0], _33584_);
  nand (_33591_, _33590_, _33589_);
  nand (_33592_, _33591_, _36029_);
  or (_33593_, \oc8051_gm_cxrom_1.cell8.data [0], _36029_);
  and (_00256_, _33593_, _33592_);
  or (_33594_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33595_, \oc8051_gm_cxrom_1.cell8.data [1], _33584_);
  nand (_33596_, _33595_, _33594_);
  nand (_33597_, _33596_, _36029_);
  or (_33598_, \oc8051_gm_cxrom_1.cell8.data [1], _36029_);
  and (_00259_, _33598_, _33597_);
  or (_33599_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33600_, \oc8051_gm_cxrom_1.cell8.data [2], _33584_);
  nand (_33601_, _33600_, _33599_);
  nand (_33602_, _33601_, _36029_);
  or (_33603_, \oc8051_gm_cxrom_1.cell8.data [2], _36029_);
  and (_00263_, _33603_, _33602_);
  or (_33604_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33605_, \oc8051_gm_cxrom_1.cell8.data [3], _33584_);
  nand (_33606_, _33605_, _33604_);
  nand (_33607_, _33606_, _36029_);
  or (_33608_, \oc8051_gm_cxrom_1.cell8.data [3], _36029_);
  and (_00266_, _33608_, _33607_);
  or (_33609_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33610_, \oc8051_gm_cxrom_1.cell8.data [4], _33584_);
  nand (_33611_, _33610_, _33609_);
  nand (_33612_, _33611_, _36029_);
  or (_33613_, \oc8051_gm_cxrom_1.cell8.data [4], _36029_);
  and (_00270_, _33613_, _33612_);
  or (_33614_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33615_, \oc8051_gm_cxrom_1.cell8.data [5], _33584_);
  nand (_33616_, _33615_, _33614_);
  nand (_33617_, _33616_, _36029_);
  or (_33618_, \oc8051_gm_cxrom_1.cell8.data [5], _36029_);
  and (_00273_, _33618_, _33617_);
  or (_33619_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33620_, \oc8051_gm_cxrom_1.cell8.data [6], _33584_);
  nand (_33621_, _33620_, _33619_);
  nand (_33622_, _33621_, _36029_);
  or (_33623_, \oc8051_gm_cxrom_1.cell8.data [6], _36029_);
  and (_00276_, _33623_, _33622_);
  or (_33624_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_33625_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_33626_, _33625_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_33627_, _33626_, _33624_);
  nand (_33628_, _33627_, _36029_);
  or (_33629_, \oc8051_gm_cxrom_1.cell9.data [7], _36029_);
  and (_00293_, _33629_, _33628_);
  or (_33630_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33631_, \oc8051_gm_cxrom_1.cell9.data [0], _33625_);
  nand (_33632_, _33631_, _33630_);
  nand (_33633_, _33632_, _36029_);
  or (_33634_, \oc8051_gm_cxrom_1.cell9.data [0], _36029_);
  and (_00299_, _33634_, _33633_);
  or (_33635_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33636_, \oc8051_gm_cxrom_1.cell9.data [1], _33625_);
  nand (_33637_, _33636_, _33635_);
  nand (_33638_, _33637_, _36029_);
  or (_33639_, \oc8051_gm_cxrom_1.cell9.data [1], _36029_);
  and (_00302_, _33639_, _33638_);
  or (_33640_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33641_, \oc8051_gm_cxrom_1.cell9.data [2], _33625_);
  nand (_33642_, _33641_, _33640_);
  nand (_33643_, _33642_, _36029_);
  or (_33644_, \oc8051_gm_cxrom_1.cell9.data [2], _36029_);
  and (_00305_, _33644_, _33643_);
  or (_33645_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33646_, \oc8051_gm_cxrom_1.cell9.data [3], _33625_);
  nand (_33647_, _33646_, _33645_);
  nand (_33648_, _33647_, _36029_);
  or (_33649_, \oc8051_gm_cxrom_1.cell9.data [3], _36029_);
  and (_00308_, _33649_, _33648_);
  or (_33650_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33651_, \oc8051_gm_cxrom_1.cell9.data [4], _33625_);
  nand (_33652_, _33651_, _33650_);
  nand (_33653_, _33652_, _36029_);
  or (_33654_, \oc8051_gm_cxrom_1.cell9.data [4], _36029_);
  and (_00312_, _33654_, _33653_);
  or (_33655_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33656_, \oc8051_gm_cxrom_1.cell9.data [5], _33625_);
  nand (_33657_, _33656_, _33655_);
  nand (_33658_, _33657_, _36029_);
  or (_33659_, \oc8051_gm_cxrom_1.cell9.data [5], _36029_);
  and (_00315_, _33659_, _33658_);
  or (_33660_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33661_, \oc8051_gm_cxrom_1.cell9.data [6], _33625_);
  nand (_33662_, _33661_, _33660_);
  nand (_33663_, _33662_, _36029_);
  or (_33664_, \oc8051_gm_cxrom_1.cell9.data [6], _36029_);
  and (_00318_, _33664_, _33663_);
  or (_33665_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_33666_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_33667_, _33666_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_33668_, _33667_, _33665_);
  nand (_33669_, _33668_, _36029_);
  or (_33670_, \oc8051_gm_cxrom_1.cell10.data [7], _36029_);
  and (_00336_, _33670_, _33669_);
  or (_33671_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33672_, \oc8051_gm_cxrom_1.cell10.data [0], _33666_);
  nand (_33673_, _33672_, _33671_);
  nand (_33674_, _33673_, _36029_);
  or (_33675_, \oc8051_gm_cxrom_1.cell10.data [0], _36029_);
  and (_00343_, _33675_, _33674_);
  or (_33676_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33677_, \oc8051_gm_cxrom_1.cell10.data [1], _33666_);
  nand (_33678_, _33677_, _33676_);
  nand (_33679_, _33678_, _36029_);
  or (_33680_, \oc8051_gm_cxrom_1.cell10.data [1], _36029_);
  and (_00347_, _33680_, _33679_);
  or (_33681_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33682_, \oc8051_gm_cxrom_1.cell10.data [2], _33666_);
  nand (_33683_, _33682_, _33681_);
  nand (_33684_, _33683_, _36029_);
  or (_33685_, \oc8051_gm_cxrom_1.cell10.data [2], _36029_);
  and (_00351_, _33685_, _33684_);
  or (_33686_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33687_, \oc8051_gm_cxrom_1.cell10.data [3], _33666_);
  nand (_33688_, _33687_, _33686_);
  nand (_33689_, _33688_, _36029_);
  or (_33690_, \oc8051_gm_cxrom_1.cell10.data [3], _36029_);
  and (_00355_, _33690_, _33689_);
  or (_33691_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33692_, \oc8051_gm_cxrom_1.cell10.data [4], _33666_);
  nand (_33694_, _33692_, _33691_);
  nand (_33695_, _33694_, _36029_);
  or (_33696_, \oc8051_gm_cxrom_1.cell10.data [4], _36029_);
  and (_00359_, _33696_, _33695_);
  or (_33697_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33699_, \oc8051_gm_cxrom_1.cell10.data [5], _33666_);
  nand (_33700_, _33699_, _33697_);
  nand (_33701_, _33700_, _36029_);
  or (_33702_, \oc8051_gm_cxrom_1.cell10.data [5], _36029_);
  and (_00363_, _33702_, _33701_);
  or (_33704_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33705_, \oc8051_gm_cxrom_1.cell10.data [6], _33666_);
  nand (_33706_, _33705_, _33704_);
  nand (_33707_, _33706_, _36029_);
  or (_33708_, \oc8051_gm_cxrom_1.cell10.data [6], _36029_);
  and (_00367_, _33708_, _33707_);
  or (_33710_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_33711_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_33712_, _33711_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_33713_, _33712_, _33710_);
  nand (_33715_, _33713_, _36029_);
  or (_33716_, \oc8051_gm_cxrom_1.cell11.data [7], _36029_);
  and (_00389_, _33716_, _33715_);
  or (_33717_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33718_, \oc8051_gm_cxrom_1.cell11.data [0], _33711_);
  nand (_33720_, _33718_, _33717_);
  nand (_33721_, _33720_, _36029_);
  or (_33722_, \oc8051_gm_cxrom_1.cell11.data [0], _36029_);
  and (_00396_, _33722_, _33721_);
  or (_33723_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33725_, \oc8051_gm_cxrom_1.cell11.data [1], _33711_);
  nand (_33726_, _33725_, _33723_);
  nand (_33728_, _33726_, _36029_);
  or (_33729_, \oc8051_gm_cxrom_1.cell11.data [1], _36029_);
  and (_00400_, _33729_, _33728_);
  or (_33730_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33731_, \oc8051_gm_cxrom_1.cell11.data [2], _33711_);
  nand (_33732_, _33731_, _33730_);
  nand (_33733_, _33732_, _36029_);
  or (_33735_, \oc8051_gm_cxrom_1.cell11.data [2], _36029_);
  and (_00404_, _33735_, _33733_);
  or (_33736_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33738_, \oc8051_gm_cxrom_1.cell11.data [3], _33711_);
  nand (_33739_, _33738_, _33736_);
  nand (_33740_, _33739_, _36029_);
  or (_33742_, \oc8051_gm_cxrom_1.cell11.data [3], _36029_);
  and (_00408_, _33742_, _33740_);
  or (_33743_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33745_, \oc8051_gm_cxrom_1.cell11.data [4], _33711_);
  nand (_33746_, _33745_, _33743_);
  nand (_33747_, _33746_, _36029_);
  or (_33749_, \oc8051_gm_cxrom_1.cell11.data [4], _36029_);
  and (_00412_, _33749_, _33747_);
  or (_33750_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33752_, \oc8051_gm_cxrom_1.cell11.data [5], _33711_);
  nand (_33753_, _33752_, _33750_);
  nand (_33754_, _33753_, _36029_);
  or (_33756_, \oc8051_gm_cxrom_1.cell11.data [5], _36029_);
  and (_00416_, _33756_, _33754_);
  or (_33758_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33759_, \oc8051_gm_cxrom_1.cell11.data [6], _33711_);
  nand (_33760_, _33759_, _33758_);
  nand (_33761_, _33760_, _36029_);
  or (_33762_, \oc8051_gm_cxrom_1.cell11.data [6], _36029_);
  and (_00420_, _33762_, _33761_);
  or (_33763_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_33765_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_33766_, _33765_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_33767_, _33766_, _33763_);
  nand (_33769_, _33767_, _36029_);
  or (_33770_, \oc8051_gm_cxrom_1.cell12.data [7], _36029_);
  and (_00442_, _33770_, _33769_);
  or (_33772_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33773_, \oc8051_gm_cxrom_1.cell12.data [0], _33765_);
  nand (_33774_, _33773_, _33772_);
  nand (_33776_, _33774_, _36029_);
  or (_33777_, \oc8051_gm_cxrom_1.cell12.data [0], _36029_);
  and (_00449_, _33777_, _33776_);
  or (_33779_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33780_, \oc8051_gm_cxrom_1.cell12.data [1], _33765_);
  nand (_33781_, _33780_, _33779_);
  nand (_33783_, _33781_, _36029_);
  or (_33784_, \oc8051_gm_cxrom_1.cell12.data [1], _36029_);
  and (_00453_, _33784_, _33783_);
  or (_33786_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33787_, \oc8051_gm_cxrom_1.cell12.data [2], _33765_);
  nand (_33789_, _33787_, _33786_);
  nand (_33790_, _33789_, _36029_);
  or (_33791_, \oc8051_gm_cxrom_1.cell12.data [2], _36029_);
  and (_00457_, _33791_, _33790_);
  or (_33792_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33794_, \oc8051_gm_cxrom_1.cell12.data [3], _33765_);
  nand (_33795_, _33794_, _33792_);
  nand (_33796_, _33795_, _36029_);
  or (_33798_, \oc8051_gm_cxrom_1.cell12.data [3], _36029_);
  and (_00461_, _33798_, _33796_);
  or (_33799_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33801_, \oc8051_gm_cxrom_1.cell12.data [4], _33765_);
  nand (_33802_, _33801_, _33799_);
  nand (_33803_, _33802_, _36029_);
  or (_33805_, \oc8051_gm_cxrom_1.cell12.data [4], _36029_);
  and (_00465_, _33805_, _33803_);
  or (_33806_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33808_, \oc8051_gm_cxrom_1.cell12.data [5], _33765_);
  nand (_33809_, _33808_, _33806_);
  nand (_33810_, _33809_, _36029_);
  or (_33812_, \oc8051_gm_cxrom_1.cell12.data [5], _36029_);
  and (_00469_, _33812_, _33810_);
  or (_33813_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33815_, \oc8051_gm_cxrom_1.cell12.data [6], _33765_);
  nand (_33816_, _33815_, _33813_);
  nand (_33818_, _33816_, _36029_);
  or (_33819_, \oc8051_gm_cxrom_1.cell12.data [6], _36029_);
  and (_00473_, _33819_, _33818_);
  or (_33820_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_33821_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_33822_, _33821_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_33823_, _33822_, _33820_);
  nand (_33825_, _33823_, _36029_);
  or (_33826_, \oc8051_gm_cxrom_1.cell13.data [7], _36029_);
  and (_00495_, _33826_, _33825_);
  or (_33828_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33829_, \oc8051_gm_cxrom_1.cell13.data [0], _33821_);
  nand (_33830_, _33829_, _33828_);
  nand (_33832_, _33830_, _36029_);
  or (_33833_, \oc8051_gm_cxrom_1.cell13.data [0], _36029_);
  and (_00502_, _33833_, _33832_);
  or (_33835_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33836_, \oc8051_gm_cxrom_1.cell13.data [1], _33821_);
  nand (_33837_, _33836_, _33835_);
  nand (_33839_, _33837_, _36029_);
  or (_33840_, \oc8051_gm_cxrom_1.cell13.data [1], _36029_);
  and (_00506_, _33840_, _33839_);
  or (_33842_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33843_, \oc8051_gm_cxrom_1.cell13.data [2], _33821_);
  nand (_33844_, _33843_, _33842_);
  nand (_33846_, _33844_, _36029_);
  or (_33847_, \oc8051_gm_cxrom_1.cell13.data [2], _36029_);
  and (_00510_, _33847_, _33846_);
  or (_33849_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33850_, \oc8051_gm_cxrom_1.cell13.data [3], _33821_);
  nand (_33851_, _33850_, _33849_);
  nand (_33853_, _33851_, _36029_);
  or (_33854_, \oc8051_gm_cxrom_1.cell13.data [3], _36029_);
  and (_00514_, _33854_, _33853_);
  or (_33856_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33857_, \oc8051_gm_cxrom_1.cell13.data [4], _33821_);
  nand (_33858_, _33857_, _33856_);
  nand (_33860_, _33858_, _36029_);
  or (_33861_, \oc8051_gm_cxrom_1.cell13.data [4], _36029_);
  and (_00518_, _33861_, _33860_);
  or (_33863_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33864_, \oc8051_gm_cxrom_1.cell13.data [5], _33821_);
  nand (_33865_, _33864_, _33863_);
  nand (_33867_, _33865_, _36029_);
  or (_33868_, \oc8051_gm_cxrom_1.cell13.data [5], _36029_);
  and (_00522_, _33868_, _33867_);
  or (_33870_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33871_, \oc8051_gm_cxrom_1.cell13.data [6], _33821_);
  nand (_33872_, _33871_, _33870_);
  nand (_33874_, _33872_, _36029_);
  or (_33875_, \oc8051_gm_cxrom_1.cell13.data [6], _36029_);
  and (_00526_, _33875_, _33874_);
  or (_33877_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_33878_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_33879_, _33878_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_33881_, _33879_, _33877_);
  nand (_33882_, _33881_, _36029_);
  or (_33883_, \oc8051_gm_cxrom_1.cell14.data [7], _36029_);
  and (_00548_, _33883_, _33882_);
  or (_33885_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33886_, \oc8051_gm_cxrom_1.cell14.data [0], _33878_);
  nand (_33888_, _33886_, _33885_);
  nand (_33889_, _33888_, _36029_);
  or (_33890_, \oc8051_gm_cxrom_1.cell14.data [0], _36029_);
  and (_00555_, _33890_, _33889_);
  or (_33892_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33893_, \oc8051_gm_cxrom_1.cell14.data [1], _33878_);
  nand (_33895_, _33893_, _33892_);
  nand (_33896_, _33895_, _36029_);
  or (_33897_, \oc8051_gm_cxrom_1.cell14.data [1], _36029_);
  and (_00559_, _33897_, _33896_);
  or (_33899_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33900_, \oc8051_gm_cxrom_1.cell14.data [2], _33878_);
  nand (_33902_, _33900_, _33899_);
  nand (_33903_, _33902_, _36029_);
  or (_33905_, \oc8051_gm_cxrom_1.cell14.data [2], _36029_);
  and (_00563_, _33905_, _33903_);
  or (_33906_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33907_, \oc8051_gm_cxrom_1.cell14.data [3], _33878_);
  nand (_33909_, _33907_, _33906_);
  nand (_33910_, _33909_, _36029_);
  or (_33911_, \oc8051_gm_cxrom_1.cell14.data [3], _36029_);
  and (_00567_, _33911_, _33910_);
  or (_33913_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33914_, \oc8051_gm_cxrom_1.cell14.data [4], _33878_);
  nand (_33916_, _33914_, _33913_);
  nand (_33917_, _33916_, _36029_);
  or (_33918_, \oc8051_gm_cxrom_1.cell14.data [4], _36029_);
  and (_00571_, _33918_, _33917_);
  or (_33920_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33921_, \oc8051_gm_cxrom_1.cell14.data [5], _33878_);
  nand (_33923_, _33921_, _33920_);
  nand (_33924_, _33923_, _36029_);
  or (_33925_, \oc8051_gm_cxrom_1.cell14.data [5], _36029_);
  and (_00575_, _33925_, _33924_);
  or (_33927_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33928_, \oc8051_gm_cxrom_1.cell14.data [6], _33878_);
  nand (_33930_, _33928_, _33927_);
  nand (_33931_, _33930_, _36029_);
  or (_33933_, \oc8051_gm_cxrom_1.cell14.data [6], _36029_);
  and (_00579_, _33933_, _33931_);
  or (_33934_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_33935_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_33936_, _33935_, \oc8051_gm_cxrom_1.cell15.data [7]);
  and (_33937_, _33936_, _33934_);
  or (_33938_, _33937_, rst);
  or (_33940_, \oc8051_gm_cxrom_1.cell15.data [7], _36029_);
  and (_00601_, _33940_, _33938_);
  or (_33941_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33943_, \oc8051_gm_cxrom_1.cell15.data [0], _33935_);
  and (_33944_, _33943_, _33941_);
  or (_33945_, _33944_, rst);
  or (_33947_, \oc8051_gm_cxrom_1.cell15.data [0], _36029_);
  and (_00608_, _33947_, _33945_);
  or (_33948_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33950_, \oc8051_gm_cxrom_1.cell15.data [1], _33935_);
  and (_33951_, _33950_, _33948_);
  or (_33952_, _33951_, rst);
  or (_33954_, \oc8051_gm_cxrom_1.cell15.data [1], _36029_);
  and (_00612_, _33954_, _33952_);
  or (_33955_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33957_, \oc8051_gm_cxrom_1.cell15.data [2], _33935_);
  and (_33958_, _33957_, _33955_);
  or (_33959_, _33958_, rst);
  or (_33961_, \oc8051_gm_cxrom_1.cell15.data [2], _36029_);
  and (_00616_, _33961_, _33959_);
  or (_33963_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33964_, \oc8051_gm_cxrom_1.cell15.data [3], _33935_);
  and (_33965_, _33964_, _33963_);
  or (_33966_, _33965_, rst);
  or (_33968_, \oc8051_gm_cxrom_1.cell15.data [3], _36029_);
  and (_00620_, _33968_, _33966_);
  or (_33969_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33971_, \oc8051_gm_cxrom_1.cell15.data [4], _33935_);
  and (_33972_, _33971_, _33969_);
  or (_33973_, _33972_, rst);
  or (_33975_, \oc8051_gm_cxrom_1.cell15.data [4], _36029_);
  and (_00624_, _33975_, _33973_);
  or (_33976_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33978_, \oc8051_gm_cxrom_1.cell15.data [5], _33935_);
  and (_33979_, _33978_, _33976_);
  or (_33980_, _33979_, rst);
  or (_33982_, \oc8051_gm_cxrom_1.cell15.data [5], _36029_);
  and (_00628_, _33982_, _33980_);
  or (_33983_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33985_, \oc8051_gm_cxrom_1.cell15.data [6], _33935_);
  and (_33986_, _33985_, _33983_);
  or (_33987_, _33986_, rst);
  or (_33989_, \oc8051_gm_cxrom_1.cell15.data [6], _36029_);
  and (_00632_, _33989_, _33987_);
  nor (_04368_, _30392_, rst);
  and (_33991_, _30002_, _36029_);
  nand (_33992_, _33991_, _30223_);
  nor (_33993_, _30259_, _30214_);
  or (_04371_, _33993_, _33992_);
  not (_33995_, _30037_);
  and (_33996_, _30083_, _30061_);
  and (_33998_, _33996_, _33995_);
  not (_33999_, _30109_);
  and (_34000_, _30154_, _30131_);
  and (_34002_, _34000_, _33999_);
  and (_34003_, _34002_, _30207_);
  and (_34004_, _34003_, _33998_);
  not (_34006_, _30083_);
  and (_34007_, _34006_, _30061_);
  not (_34008_, _30176_);
  not (_34010_, _30154_);
  nor (_34011_, _34010_, _30131_);
  and (_34012_, _30207_, _30109_);
  and (_34014_, _34012_, _34011_);
  and (_34015_, _34014_, _34008_);
  not (_34016_, _30207_);
  and (_34018_, _34002_, _34016_);
  and (_34019_, _34018_, _30037_);
  or (_34021_, _34019_, _34015_);
  and (_34022_, _34021_, _34007_);
  or (_34023_, _34022_, _34004_);
  nor (_34024_, _30083_, _30061_);
  and (_34026_, _34024_, _33995_);
  and (_34027_, _34012_, _34000_);
  and (_34028_, _30131_, _33999_);
  and (_34030_, _34008_, _30154_);
  and (_34031_, _34030_, _34028_);
  or (_34032_, _34031_, _34027_);
  and (_34034_, _34032_, _34026_);
  nor (_34035_, _30037_, _34008_);
  and (_34036_, _34007_, _34035_);
  not (_34038_, _34036_);
  nor (_34039_, _34038_, _34000_);
  and (_34040_, _30176_, _30154_);
  and (_34042_, _34026_, _34028_);
  and (_34043_, _34042_, _34040_);
  and (_34044_, _30037_, _30176_);
  and (_34046_, _34024_, _34044_);
  and (_34047_, _34046_, _34010_);
  or (_34048_, _34047_, _34043_);
  or (_34050_, _34048_, _34039_);
  and (_34051_, _30037_, _34008_);
  nor (_34053_, _34051_, _34035_);
  and (_34054_, _34053_, _33996_);
  and (_34055_, _34054_, _34027_);
  and (_34056_, _34051_, _34007_);
  and (_34057_, _34027_, _34056_);
  or (_34059_, _34057_, _34055_);
  or (_34060_, _34059_, _34050_);
  or (_34061_, _34060_, _34034_);
  not (_34063_, _30061_);
  and (_34064_, _30083_, _34063_);
  and (_34065_, _34064_, _34051_);
  and (_34067_, _34065_, _34027_);
  and (_34068_, _34035_, _33996_);
  and (_34069_, _34027_, _34068_);
  and (_34071_, _34000_, _30109_);
  not (_34072_, _34071_);
  nor (_34073_, _30037_, _30176_);
  and (_34075_, _34064_, _34073_);
  nor (_34076_, _34075_, _34016_);
  nor (_34077_, _34076_, _34072_);
  or (_34079_, _34077_, _34069_);
  nor (_34080_, _34079_, _34067_);
  and (_34081_, _34064_, _34035_);
  and (_34083_, _34081_, _34018_);
  and (_34084_, _34011_, _30109_);
  and (_34086_, _34084_, _34016_);
  and (_34087_, _34086_, _34046_);
  or (_34088_, _34087_, _34083_);
  and (_34089_, _34064_, _30176_);
  and (_34091_, _34089_, _34027_);
  and (_34092_, _33996_, _30037_);
  and (_34093_, _34092_, _34003_);
  or (_34095_, _34093_, _34091_);
  nor (_34096_, _34095_, _34088_);
  nand (_34097_, _34096_, _34080_);
  or (_34099_, _34097_, _34061_);
  or (_34100_, _34099_, _34023_);
  and (_34101_, _34100_, _30003_);
  not (_34103_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_34104_, _30001_, _14692_);
  and (_34105_, _34104_, _30272_);
  nor (_34107_, _34105_, _34103_);
  or (_34108_, _34107_, rst);
  or (_04374_, _34108_, _34101_);
  nand (_34110_, _30083_, _29997_);
  or (_34111_, _29997_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_34112_, _34111_, _36029_);
  and (_04377_, _34112_, _34110_);
  and (_34114_, \oc8051_top_1.oc8051_sfr1.wait_data , _36029_);
  and (_34116_, _34114_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_34117_, _30363_, _30298_);
  and (_34118_, _30297_, _30246_);
  and (_34119_, _30265_, _30259_);
  and (_34121_, _30257_, _30214_);
  or (_34122_, _34121_, _34119_);
  or (_34123_, _34122_, _34118_);
  or (_34125_, _34123_, _34117_);
  not (_34126_, _30346_);
  and (_34127_, _30380_, _30327_);
  and (_34129_, _30246_, _30231_);
  and (_34130_, _34129_, _30180_);
  or (_34131_, _34130_, _34127_);
  or (_34133_, _34131_, _34126_);
  or (_34134_, _34133_, _34125_);
  and (_34135_, _34134_, _33991_);
  or (_04380_, _34135_, _34116_);
  and (_34137_, _30219_, _30041_);
  nor (_34138_, _30181_, _30158_);
  and (_34140_, _34138_, _34137_);
  and (_34141_, _34140_, _30088_);
  or (_34142_, _34141_, _30229_);
  and (_34144_, _30285_, _30113_);
  and (_34145_, _34144_, _30297_);
  or (_34147_, _34145_, _34142_);
  and (_34148_, _30259_, _30253_);
  or (_34149_, _34148_, _30247_);
  or (_34150_, _34149_, _34147_);
  and (_34152_, _34150_, _30002_);
  and (_34153_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34154_, \oc8051_top_1.oc8051_decoder1.state [0], _14692_);
  and (_34156_, _34154_, _34103_);
  not (_34157_, _30383_);
  and (_34158_, _34157_, _34156_);
  or (_34160_, _34158_, _34153_);
  or (_34161_, _34160_, _34152_);
  and (_04383_, _34161_, _36029_);
  and (_34163_, _34114_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_34164_, _30380_, _30347_);
  nor (_34165_, _30347_, _30257_);
  nor (_34167_, _34165_, _30325_);
  or (_34168_, _34167_, _34164_);
  and (_34169_, _34144_, _30303_);
  or (_34171_, _34169_, _34168_);
  not (_34172_, _30189_);
  nor (_34173_, _34165_, _30158_);
  nor (_34175_, _30180_, _30158_);
  and (_34176_, _34175_, _30187_);
  or (_34177_, _34176_, _34173_);
  or (_34178_, _34177_, _34172_);
  and (_34179_, _30380_, _30321_);
  and (_34180_, _30295_, _30351_);
  or (_34181_, _34180_, _34179_);
  or (_34182_, _34181_, _34149_);
  or (_34183_, _34182_, _34178_);
  or (_34184_, _34183_, _34171_);
  and (_34185_, _34184_, _33991_);
  or (_04386_, _34185_, _34163_);
  and (_34186_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34187_, _30314_, _30002_);
  or (_34188_, _34187_, _34186_);
  or (_34189_, _34188_, _34158_);
  and (_04389_, _34189_, _36029_);
  and (_34190_, _30135_, _30212_);
  and (_34191_, _30245_, _30158_);
  and (_34192_, _34191_, _34190_);
  and (_34193_, _34192_, _30231_);
  and (_34194_, _30327_, _30259_);
  and (_34195_, _30327_, _30214_);
  or (_34196_, _34195_, _34194_);
  or (_34197_, _34196_, _34193_);
  and (_34198_, _34197_, _34156_);
  or (_34199_, _34198_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34200_, _30286_, _30213_);
  and (_34201_, _30215_, _30187_);
  nor (_34202_, _34201_, _34200_);
  nor (_34203_, _34202_, _30180_);
  not (_34204_, _29998_);
  and (_34205_, _34130_, _34204_);
  or (_34206_, _34205_, _34203_);
  and (_34207_, _34206_, _30272_);
  or (_34208_, _34207_, _34199_);
  or (_34209_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _14692_);
  and (_34210_, _34209_, _36029_);
  and (_04392_, _34210_, _34208_);
  and (_34211_, _34114_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_34212_, _34175_, _30228_);
  or (_34213_, _34176_, _34212_);
  or (_34214_, _30303_, _30297_);
  and (_34215_, _34214_, _30185_);
  or (_34216_, _34215_, _34213_);
  and (_34217_, _30215_, _30090_);
  or (_34218_, _34169_, _34121_);
  or (_34219_, _34218_, _34217_);
  or (_34220_, _34141_, _30336_);
  or (_34221_, _30288_, _30247_);
  or (_34222_, _34221_, _34220_);
  or (_34223_, _34222_, _34219_);
  or (_34224_, _34223_, _34216_);
  and (_34225_, _34224_, _33991_);
  or (_04395_, _34225_, _34211_);
  and (_34226_, _34114_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_34227_, _34145_, _30305_);
  and (_34228_, _30246_, _30186_);
  and (_34229_, _34144_, _30262_);
  or (_34230_, _34229_, _34228_);
  or (_34231_, _34230_, _34227_);
  or (_34232_, _34231_, _34177_);
  and (_34233_, _30228_, _30183_);
  and (_34234_, _34137_, _30218_);
  or (_34235_, _34234_, _30263_);
  or (_34236_, _34235_, _34233_);
  and (_34237_, _30380_, _30290_);
  or (_34238_, _34237_, _30293_);
  or (_34239_, _34238_, _34236_);
  or (_34240_, _34239_, _34232_);
  nor (_34241_, _30311_, _30188_);
  not (_34242_, _34241_);
  not (_34243_, _30302_);
  and (_34244_, _34138_, _30250_);
  or (_34245_, _34244_, _34140_);
  or (_34246_, _34245_, _34243_);
  or (_34247_, _34246_, _34242_);
  or (_34248_, _34247_, _34171_);
  or (_34249_, _34248_, _34240_);
  and (_34250_, _34249_, _33991_);
  or (_04398_, _34250_, _34226_);
  and (_34251_, _34144_, _30216_);
  or (_34252_, _34251_, _30232_);
  and (_34253_, _30216_, _30185_);
  and (_34254_, _34175_, _30231_);
  or (_34255_, _34254_, _34253_);
  and (_34256_, _30216_, _30351_);
  or (_34257_, _34256_, _34255_);
  or (_34258_, _34257_, _34252_);
  and (_34259_, _34144_, _30253_);
  or (_34260_, _34259_, _34258_);
  and (_34261_, _34260_, _30002_);
  nand (_34262_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_34263_, _34262_, _30389_);
  or (_34264_, _34263_, _34261_);
  and (_04401_, _34264_, _36029_);
  or (_34265_, _30336_, _30332_);
  not (_34266_, _30299_);
  or (_34267_, _34167_, _34266_);
  or (_34268_, _34267_, _34265_);
  and (_34269_, _30249_, _30181_);
  and (_34270_, _34269_, _30287_);
  or (_34271_, _34270_, _30304_);
  and (_34272_, _30303_, _30215_);
  or (_34273_, _34272_, _30291_);
  nor (_34274_, _34273_, _34271_);
  nand (_34275_, _34274_, _30316_);
  or (_34276_, _34275_, _34268_);
  and (_34277_, _34175_, _30249_);
  or (_34278_, _34277_, _30352_);
  and (_34279_, _34200_, _30181_);
  and (_34280_, _34138_, _30231_);
  or (_34281_, _34280_, _34279_);
  or (_34282_, _34281_, _34142_);
  or (_34283_, _34282_, _34278_);
  and (_34284_, _34269_, _30185_);
  or (_34285_, _34284_, _30188_);
  or (_34286_, _34285_, _30350_);
  or (_34287_, _30318_, _30266_);
  or (_34288_, _34287_, _34286_);
  or (_34289_, _34288_, _34283_);
  or (_34290_, _34289_, _34177_);
  or (_34291_, _34290_, _34276_);
  and (_34292_, _34291_, _30002_);
  and (_34293_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34294_, _30369_, _30274_);
  or (_34295_, _34272_, _34279_);
  and (_34296_, _34295_, _30274_);
  or (_34297_, _34296_, _34158_);
  or (_34298_, _34297_, _34294_);
  or (_34299_, _34298_, _34293_);
  or (_34300_, _34299_, _34292_);
  and (_04404_, _34300_, _36029_);
  nor (_04464_, _30280_, rst);
  nor (_04466_, _30375_, rst);
  not (_34301_, _33991_);
  not (_34302_, _33993_);
  and (_34303_, _34302_, _30327_);
  nor (_34304_, _34303_, _34129_);
  or (_04469_, _34304_, _34301_);
  nand (_34305_, _34129_, _33991_);
  or (_34306_, _33992_, _30342_);
  and (_04472_, _34306_, _34305_);
  or (_34307_, _34023_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_34308_, _34307_, _34105_);
  nor (_34309_, _34104_, _30272_);
  or (_34310_, _34309_, rst);
  or (_04475_, _34310_, _34308_);
  nand (_34311_, _30207_, _29997_);
  or (_34312_, _29997_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_34313_, _34312_, _36029_);
  and (_04478_, _34313_, _34311_);
  nand (_34314_, _30109_, _29997_);
  or (_34315_, _29997_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_34316_, _34315_, _36029_);
  and (_04481_, _34316_, _34314_);
  nand (_34317_, _30131_, _29997_);
  or (_34318_, _29997_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_34319_, _34318_, _36029_);
  and (_04484_, _34319_, _34317_);
  nand (_34320_, _30154_, _29997_);
  or (_34321_, _29997_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_34322_, _34321_, _36029_);
  and (_04487_, _34322_, _34320_);
  nand (_34323_, _34008_, _29997_);
  or (_34324_, _29997_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_34325_, _34324_, _36029_);
  and (_04490_, _34325_, _34323_);
  nand (_34326_, _30037_, _29997_);
  or (_34327_, _29997_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34328_, _34327_, _36029_);
  and (_04493_, _34328_, _34326_);
  nand (_34329_, _30061_, _29997_);
  or (_34330_, _29997_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34331_, _34330_, _36029_);
  and (_04496_, _34331_, _34329_);
  or (_34332_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _14692_);
  and (_34333_, _34332_, _34199_);
  or (_34334_, _34148_, _30300_);
  or (_34335_, _34334_, _34237_);
  and (_34336_, _30223_, _30181_);
  and (_34337_, _34336_, _30380_);
  and (_34338_, _34144_, _30238_);
  or (_34339_, _34338_, _34337_);
  and (_34340_, _30380_, _30251_);
  and (_34341_, _30327_, _30351_);
  or (_34342_, _34341_, _34340_);
  or (_34343_, _34342_, _34339_);
  or (_34344_, _34244_, _34127_);
  and (_34345_, _30238_, _30185_);
  or (_34346_, _34345_, _34229_);
  or (_34347_, _34346_, _34344_);
  or (_34348_, _34347_, _34343_);
  or (_34349_, _34348_, _34335_);
  or (_34350_, _30257_, _30187_);
  and (_34351_, _34350_, _30380_);
  and (_34352_, _34175_, _30221_);
  or (_34353_, _34352_, _34256_);
  or (_34354_, _34259_, _34228_);
  or (_34355_, _34354_, _34353_);
  or (_34356_, _34355_, _34351_);
  and (_34357_, _30253_, _30185_);
  or (_34358_, _30263_, _34357_);
  or (_34359_, _30328_, _30247_);
  or (_34360_, _34359_, _34358_);
  and (_34361_, _34138_, _30221_);
  or (_34362_, _34251_, _34361_);
  or (_34363_, _34362_, _30225_);
  or (_34364_, _34363_, _34255_);
  or (_34365_, _34364_, _34360_);
  or (_34366_, _34365_, _34356_);
  or (_34367_, _34366_, _34349_);
  and (_34368_, _34367_, _30002_);
  or (_34369_, _34368_, _34333_);
  and (_28683_, _34369_, _36029_);
  and (_34370_, _34114_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_34371_, _30290_, _30262_);
  and (_34372_, _34371_, _30215_);
  or (_34373_, _34372_, _34245_);
  and (_34374_, _30065_, _30042_);
  and (_34375_, _34175_, _34374_);
  and (_34376_, _34375_, _30088_);
  nor (_34377_, _34376_, _30184_);
  not (_34378_, _30380_);
  or (_34379_, _34378_, _30240_);
  nand (_34380_, _34379_, _34377_);
  or (_34381_, _34380_, _34373_);
  or (_34382_, _34335_, _34236_);
  and (_34383_, _30380_, _30262_);
  nor (_34384_, _34383_, _34179_);
  nand (_34385_, _34384_, _30337_);
  or (_34386_, _34385_, _34131_);
  or (_34387_, _34386_, _34382_);
  or (_34388_, _34387_, _34381_);
  and (_34389_, _34388_, _33991_);
  or (_28685_, _34389_, _34370_);
  or (_34390_, _34287_, _34281_);
  or (_34391_, _34390_, _34276_);
  and (_34392_, _34391_, _30002_);
  and (_34393_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34394_, _34393_, _34298_);
  or (_34395_, _34394_, _34392_);
  and (_28687_, _34395_, _36029_);
  and (_34396_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34397_, _34396_, _34297_);
  and (_34398_, _34397_, _36029_);
  and (_34399_, _30310_, _30180_);
  or (_34400_, _34399_, _30229_);
  or (_34401_, _34400_, _34286_);
  or (_34402_, _34401_, _34203_);
  and (_34403_, _34402_, _33991_);
  or (_28689_, _34403_, _34398_);
  and (_34404_, _34270_, _30088_);
  and (_34405_, _30238_, _30215_);
  and (_34406_, _34251_, _30180_);
  or (_34407_, _34406_, _34405_);
  or (_34408_, _34407_, _34404_);
  or (_34409_, _34408_, _34203_);
  and (_34410_, _30221_, _30183_);
  or (_34411_, _34255_, _34410_);
  or (_34412_, _34129_, _30382_);
  and (_34413_, _34251_, _30181_);
  or (_34414_, _34413_, _34338_);
  or (_34415_, _34414_, _34412_);
  or (_34416_, _34415_, _34411_);
  or (_34417_, _34416_, _34409_);
  and (_34418_, _30380_, _30297_);
  or (_34419_, _34354_, _34418_);
  or (_34420_, _34419_, _34353_);
  and (_34421_, _34144_, _30295_);
  or (_34422_, _34421_, _34127_);
  or (_34423_, _34337_, _30381_);
  or (_34424_, _34423_, _34351_);
  or (_34425_, _34424_, _34422_);
  or (_34426_, _34284_, _34277_);
  or (_34427_, _34426_, _34357_);
  or (_34428_, _34237_, _30252_);
  or (_34429_, _34340_, _34383_);
  or (_34430_, _34429_, _34428_);
  or (_34431_, _34430_, _34427_);
  or (_34432_, _34431_, _34425_);
  or (_34433_, _34432_, _34420_);
  or (_34434_, _34433_, _34417_);
  and (_34435_, _34434_, _30002_);
  and (_34436_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_34437_, _30383_, _34204_);
  or (_34438_, _34198_, _34437_);
  or (_34439_, _34438_, _34436_);
  or (_34440_, _34439_, _34435_);
  and (_28691_, _34440_, _36029_);
  or (_34441_, _30311_, _30291_);
  and (_34442_, _34441_, _30245_);
  or (_34443_, _30382_, _30318_);
  and (_34444_, _30223_, _30183_);
  or (_34445_, _34444_, _34148_);
  or (_34446_, _34445_, _34443_);
  or (_34447_, _34446_, _34411_);
  or (_34448_, _34447_, _34442_);
  and (_34449_, _34175_, _30223_);
  or (_34450_, _34449_, _34270_);
  nor (_34451_, _34450_, _34357_);
  nand (_34452_, _34451_, _30255_);
  or (_34453_, _34452_, _30326_);
  or (_34454_, _34453_, _34425_);
  or (_34455_, _34454_, _34420_);
  or (_34456_, _34455_, _34448_);
  and (_34457_, _34456_, _30002_);
  and (_34458_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34459_, _34458_, _34438_);
  or (_34460_, _34459_, _34457_);
  and (_28693_, _34460_, _36029_);
  and (_34461_, _34114_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_34462_, _30246_, _30295_);
  and (_34463_, _30343_, _30351_);
  and (_34464_, _34253_, _30181_);
  or (_34465_, _34464_, _34463_);
  or (_34466_, _34465_, _34462_);
  or (_34467_, _34466_, _34216_);
  and (_34468_, _30246_, _30187_);
  and (_34469_, _34468_, _30181_);
  and (_34470_, _34121_, _30245_);
  or (_34471_, _34470_, _34469_);
  not (_34472_, _31840_);
  or (_34473_, _34259_, _34472_);
  or (_34474_, _34473_, _34471_);
  or (_34475_, _34474_, _34467_);
  or (_34476_, _34254_, _34141_);
  and (_34477_, _30380_, _30257_);
  or (_34478_, _34477_, _34169_);
  or (_34479_, _34478_, _34265_);
  or (_34480_, _34479_, _34476_);
  or (_34481_, _30313_, _34357_);
  and (_34482_, _30246_, _30343_);
  or (_34483_, _34482_, _34413_);
  or (_34484_, _34483_, _34481_);
  not (_34485_, _31839_);
  or (_34486_, _34221_, _34485_);
  or (_34487_, _34486_, _34484_);
  or (_34488_, _34487_, _34480_);
  or (_34489_, _34488_, _34475_);
  and (_34490_, _34489_, _33991_);
  or (_28695_, _34490_, _34461_);
  or (_34491_, _34406_, _34233_);
  or (_34492_, _34234_, _34145_);
  or (_34493_, _34492_, _34491_);
  or (_34494_, _34493_, _34238_);
  or (_34495_, _34494_, _34415_);
  or (_34496_, _34482_, _34477_);
  or (_34497_, _34469_, _34353_);
  or (_34498_, _34497_, _34496_);
  or (_34499_, _34140_, _30247_);
  or (_34500_, _30300_, _30252_);
  or (_34501_, _34500_, _34499_);
  or (_34502_, _30320_, _30241_);
  or (_34503_, _34502_, _34501_);
  or (_34504_, _34503_, _34498_);
  or (_34505_, _34504_, _34495_);
  and (_34506_, _34505_, _33991_);
  and (_34507_, _29998_, _36029_);
  and (_34508_, _34507_, _30382_);
  and (_34509_, _34114_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_34510_, _34509_, _34508_);
  or (_28697_, _34510_, _34506_);
  and (_34511_, _30246_, _30216_);
  or (_34512_, _34259_, _34180_);
  or (_34513_, _34512_, _34511_);
  or (_34514_, _34145_, _30301_);
  or (_34515_, _34514_, _30235_);
  or (_34516_, _34515_, _34513_);
  not (_34517_, _30317_);
  nor (_34518_, _34338_, _30318_);
  and (_34519_, _34518_, _34517_);
  not (_34520_, _34519_);
  or (_34521_, _34337_, _30296_);
  or (_34522_, _34521_, _34462_);
  or (_34523_, _34522_, _34520_);
  or (_34524_, _34523_, _34516_);
  or (_34525_, _34352_, _34410_);
  or (_34526_, _34476_, _34422_);
  or (_34527_, _34526_, _34525_);
  or (_34528_, _34527_, _34178_);
  or (_34529_, _34528_, _34171_);
  or (_34530_, _34529_, _34524_);
  and (_34531_, _34530_, _30002_);
  and (_34532_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34533_, _34532_, _30387_);
  or (_34534_, _34533_, _34531_);
  and (_28699_, _34534_, _36029_);
  or (_34535_, _34478_, _34220_);
  not (_34536_, _34518_);
  or (_34537_, _34525_, _34536_);
  or (_34538_, _34537_, _34535_);
  or (_34539_, _30229_, _30188_);
  nor (_34540_, _34539_, _34468_);
  nand (_34541_, _34540_, _31840_);
  or (_34542_, _34541_, _34177_);
  or (_34543_, _34522_, _34168_);
  or (_34544_, _34543_, _34542_);
  or (_34545_, _34544_, _34538_);
  and (_34546_, _34545_, _30002_);
  and (_34547_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34548_, _34547_, _30388_);
  or (_34549_, _34548_, _34546_);
  and (_28701_, _34549_, _36029_);
  and (_34550_, _34114_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_34551_, _34118_, _30333_);
  nand (_34552_, _34551_, _31839_);
  not (_34553_, _30213_);
  or (_34554_, _30246_, _34553_);
  and (_34555_, _34554_, _30295_);
  or (_34556_, _34555_, _34496_);
  or (_34557_, _34556_, _34552_);
  or (_34558_, _34471_, _34258_);
  or (_34559_, _34558_, _34473_);
  or (_34560_, _34559_, _34557_);
  and (_34561_, _34560_, _33991_);
  or (_28704_, _34561_, _34550_);
  nor (_30768_, _30083_, rst);
  nor (_30770_, _31993_, rst);
  nor (_34562_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_34563_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_34564_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_34565_, _34564_, _34563_);
  and (_34566_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_34567_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34568_, _34567_, _34566_);
  and (_34569_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_34570_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34571_, _34570_, _34569_);
  and (_34572_, _34571_, _34568_);
  and (_34573_, _34572_, _34565_);
  and (_34574_, _34573_, _30093_);
  nor (_34575_, _34574_, _34562_);
  nor (_34576_, _34575_, _31856_);
  nor (_34577_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nor (_34578_, _34577_, _34576_);
  and (_30771_, _34578_, _36029_);
  nor (_30783_, _30207_, rst);
  nor (_30784_, _30109_, rst);
  nor (_30785_, _30131_, rst);
  nor (_30786_, _30154_, rst);
  and (_30787_, _30176_, _36029_);
  nor (_30788_, _30037_, rst);
  nor (_30789_, _30061_, rst);
  nor (_30791_, _32050_, rst);
  nor (_30792_, _32166_, rst);
  nor (_30793_, _31872_, rst);
  nor (_30794_, _32075_, rst);
  nor (_30795_, _32205_, rst);
  nor (_30797_, _31932_, rst);
  nor (_30798_, _32137_, rst);
  nor (_34579_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_34580_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_34581_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_34582_, _34581_, _34580_);
  and (_34583_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_34584_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_34585_, _34584_, _34583_);
  and (_34586_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_34587_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_34588_, _34587_, _34586_);
  and (_34589_, _34588_, _34585_);
  and (_34590_, _34589_, _34582_);
  and (_34591_, _34590_, _30093_);
  nor (_34592_, _34591_, _34579_);
  nor (_34593_, _34592_, _31856_);
  nor (_34594_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_34595_, _34594_, _34593_);
  and (_30799_, _34595_, _36029_);
  nor (_34596_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_34597_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_34598_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_34599_, _34598_, _34597_);
  and (_34600_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_34601_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_34602_, _34601_, _34600_);
  and (_34603_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_34604_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34605_, _34604_, _34603_);
  and (_34606_, _34605_, _34602_);
  and (_34607_, _34606_, _34599_);
  and (_34608_, _34607_, _30093_);
  nor (_34609_, _34608_, _34596_);
  nor (_34610_, _34609_, _31856_);
  nor (_34611_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nor (_34612_, _34611_, _34610_);
  and (_30800_, _34612_, _36029_);
  nor (_34613_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_34614_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_34615_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_34616_, _34615_, _34614_);
  and (_34617_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_34618_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_34619_, _34618_, _34617_);
  and (_34620_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_34621_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_34622_, _34621_, _34620_);
  and (_34623_, _34622_, _34619_);
  and (_34624_, _34623_, _34616_);
  and (_34625_, _34624_, _30093_);
  nor (_34626_, _34625_, _34613_);
  nor (_34627_, _34626_, _31856_);
  nor (_34628_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nor (_34629_, _34628_, _34627_);
  and (_30801_, _34629_, _36029_);
  nor (_34630_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_34631_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_34632_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_34633_, _34632_, _34631_);
  and (_34634_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_34635_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_34636_, _34635_, _34634_);
  and (_34637_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_34638_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_34639_, _34638_, _34637_);
  and (_34640_, _34639_, _34636_);
  and (_34641_, _34640_, _34633_);
  and (_34642_, _34641_, _30093_);
  nor (_34643_, _34642_, _34630_);
  nor (_34644_, _34643_, _31856_);
  nor (_34645_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  nor (_34646_, _34645_, _34644_);
  and (_30803_, _34646_, _36029_);
  nor (_34647_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_34648_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_34649_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_34650_, _34649_, _34648_);
  and (_34651_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_34652_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_34653_, _34652_, _34651_);
  and (_34654_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_34655_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_34656_, _34655_, _34654_);
  and (_34657_, _34656_, _34653_);
  and (_34658_, _34657_, _34650_);
  and (_34659_, _34658_, _30093_);
  nor (_34660_, _34659_, _34647_);
  nor (_34661_, _34660_, _31856_);
  nor (_34662_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  nor (_34663_, _34662_, _34661_);
  and (_30804_, _34663_, _36029_);
  nor (_34664_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_34665_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_34666_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34667_, _34666_, _34665_);
  and (_34668_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34669_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34670_, _34669_, _34668_);
  and (_34671_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_34672_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_34673_, _34672_, _34671_);
  and (_34674_, _34673_, _34670_);
  and (_34675_, _34674_, _34667_);
  and (_34676_, _34675_, _30093_);
  nor (_34677_, _34676_, _34664_);
  nor (_34678_, _34677_, _31856_);
  nor (_34679_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  nor (_34680_, _34679_, _34678_);
  and (_30805_, _34680_, _36029_);
  nor (_34681_, _30093_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_34682_, _30024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_34683_, _30028_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_34684_, _34683_, _34682_);
  and (_34685_, _30017_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34686_, _30021_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_34687_, _34686_, _34685_);
  and (_34688_, _30011_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_34689_, _30013_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_34690_, _34689_, _34688_);
  and (_34691_, _34690_, _34687_);
  and (_34692_, _34691_, _34684_);
  and (_34693_, _34692_, _30093_);
  nor (_34694_, _34693_, _34681_);
  nor (_34695_, _34694_, _31856_);
  nor (_34696_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  nor (_34697_, _34696_, _34695_);
  and (_30806_, _34697_, _36029_);
  and (_34698_, _30003_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_34699_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_34700_, _34698_, _30578_);
  and (_34701_, _34700_, _36029_);
  and (_30832_, _34701_, _34699_);
  not (_34702_, _34698_);
  or (_34703_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _34698_, _36029_);
  and (_34704_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _36029_);
  or (_34705_, _34704_, _00000_);
  and (_30833_, _34705_, _34703_);
  nor (_30871_, _32013_, rst);
  and (_30873_, _32208_, _36029_);
  nor (_30874_, _32008_, rst);
  nor (_34706_, _32058_, _24056_);
  and (_34707_, _32058_, _24056_);
  nor (_34708_, _34707_, _34706_);
  and (_34709_, _32190_, _29704_);
  nor (_34710_, _31915_, _24319_);
  and (_34711_, _31915_, _24319_);
  nor (_34712_, _34711_, _34710_);
  or (_34713_, _34712_, _34709_);
  or (_34714_, _34713_, _34708_);
  nor (_34715_, _32013_, _23420_);
  and (_34716_, _32013_, _23420_);
  nor (_34717_, _34716_, _34715_);
  nor (_34718_, _32142_, _23287_);
  and (_34719_, _32142_, _23287_);
  nor (_34720_, _34719_, _34718_);
  nor (_34721_, _34720_, _34717_);
  nor (_34722_, _32230_, _23770_);
  and (_34723_, _32230_, _23770_);
  nor (_34724_, _34723_, _34722_);
  nor (_34725_, _31953_, _23924_);
  and (_34726_, _31953_, _23924_);
  nor (_34727_, _34726_, _34725_);
  nor (_34728_, _34727_, _34724_);
  nor (_34729_, _32095_, _23606_);
  and (_34730_, _32095_, _23606_);
  nor (_34731_, _34730_, _34729_);
  not (_34732_, _34731_);
  nor (_34733_, _32190_, _29704_);
  nor (_34734_, _34733_, _31507_);
  and (_34735_, _34734_, _34732_);
  and (_34736_, _34735_, _34728_);
  nand (_34737_, _34736_, _34721_);
  nor (_34738_, _34737_, _34714_);
  nor (_34739_, _23420_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_34740_, _34739_, _34738_);
  not (_34741_, _34740_);
  and (_34742_, _34732_, _34728_);
  and (_34743_, _34742_, _34721_);
  nor (_34744_, _30346_, _34154_);
  nor (_34745_, _27836_, _31093_);
  and (_34746_, _34745_, _34744_);
  and (_34747_, _34746_, _34743_);
  and (_34748_, _34192_, _30251_);
  nor (_34749_, _34748_, _34119_);
  and (_34750_, _29268_, _25083_);
  nand (_34751_, _34750_, _29719_);
  nor (_34752_, _34751_, _29785_);
  and (_34753_, _34752_, _29861_);
  and (_34754_, _34753_, _29935_);
  and (_34755_, _31956_, _31967_);
  nor (_34756_, _34755_, _34154_);
  or (_34757_, _34756_, _30364_);
  nor (_34758_, _34757_, _27988_);
  and (_34759_, _34758_, _34754_);
  and (_34760_, _34759_, _25699_);
  and (_34761_, _34744_, _25446_);
  or (_34762_, _34744_, _30041_);
  and (_34763_, _34762_, _30364_);
  and (_34764_, _34763_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_34765_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_34766_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_34767_, _34766_, _34765_);
  nor (_34768_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_34769_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_34770_, _34769_, _34768_);
  and (_34771_, _34770_, _34767_);
  and (_34772_, _34771_, _30276_);
  or (_34773_, _34772_, _34764_);
  or (_34774_, _34773_, _34761_);
  nor (_34775_, _34774_, _34760_);
  or (_34776_, _30251_, _30343_);
  nor (_34777_, _34776_, _30238_);
  or (_34778_, _34777_, _30342_);
  not (_34779_, _34212_);
  nor (_34780_, _34421_, _30288_);
  and (_34781_, _34780_, _34779_);
  and (_34782_, _34781_, _34377_);
  nand (_34783_, _34782_, _34778_);
  nand (_34784_, _34783_, _34775_);
  nand (_34785_, _30363_, _30180_);
  and (_34786_, _34785_, _30370_);
  or (_34787_, _34786_, _34775_);
  and (_34788_, _34787_, _34784_);
  and (_34789_, _34788_, _34749_);
  or (_34790_, _34789_, _30365_);
  nor (_34791_, _34202_, _29998_);
  nor (_34792_, _34791_, _30277_);
  and (_34793_, _34792_, _34790_);
  or (_34794_, _30990_, _30980_);
  or (_34795_, _34794_, _30958_);
  and (_34796_, _34795_, _34763_);
  nor (_34797_, _31104_, _31087_);
  nand (_34798_, _34797_, _31100_);
  and (_34799_, _34798_, _30276_);
  or (_34800_, _34799_, _34796_);
  nor (_34801_, _34800_, _34793_);
  not (_34802_, _34801_);
  nor (_34803_, _34802_, _34747_);
  and (_34804_, _34803_, _34741_);
  nor (_34805_, _30278_, rst);
  and (_30878_, _34805_, _34804_);
  and (_30879_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _36029_);
  and (_30880_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _36029_);
  nor (_34806_, _30016_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34807_, _34806_, _31856_);
  nor (_34808_, _34807_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_34809_, _34808_);
  and (_34810_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_34811_, _34810_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_34812_, _34811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_34813_, _34812_, _34809_);
  and (_34814_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_34815_, _34814_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_34816_, _34815_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_34817_, _34816_, _34813_);
  and (_34818_, _34817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_34819_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_34820_, _34819_, _34818_);
  and (_34821_, _34820_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_34822_, _34821_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_34823_, _34822_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_34824_, _34822_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_34825_, _34824_, _34823_);
  or (_34826_, _34825_, _34804_);
  and (_34827_, _34826_, _36029_);
  and (_34828_, _34377_, _34755_);
  and (_34829_, _34828_, _34780_);
  nor (_34830_, _34829_, _30365_);
  not (_34831_, _34830_);
  not (_34832_, _30278_);
  and (_34833_, _34201_, _34204_);
  and (_34834_, _30340_, _34204_);
  nor (_34835_, _34834_, _34833_);
  and (_34836_, _34835_, _34832_);
  and (_34837_, _34836_, _34831_);
  and (_34838_, _34837_, _31993_);
  nor (_34839_, _34837_, _34578_);
  nor (_34840_, _34839_, _34838_);
  not (_34841_, _34840_);
  and (_34842_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_34843_, _34842_);
  nor (_34844_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_34845_, _34844_, _34842_);
  and (_34846_, _34837_, _32137_);
  nor (_34847_, _34837_, _34697_);
  nor (_34848_, _34847_, _34846_);
  and (_34849_, _34848_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34850_, _34848_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34851_, _34850_, _34849_);
  and (_34852_, _34837_, _31932_);
  nor (_34853_, _34837_, _34680_);
  nor (_34854_, _34853_, _34852_);
  and (_34855_, _34854_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_34856_, _34854_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_34857_, _34837_, _32205_);
  nor (_34858_, _34837_, _34663_);
  nor (_34859_, _34858_, _34857_);
  nand (_34860_, _34859_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34861_, _34837_, _32075_);
  nor (_34862_, _34837_, _34646_);
  nor (_34863_, _34862_, _34861_);
  and (_34864_, _34863_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_34865_, _34863_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34866_, _34837_, _31872_);
  nor (_34867_, _34837_, _34629_);
  nor (_34868_, _34867_, _34866_);
  and (_34869_, _34868_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_34870_, _34837_, _32166_);
  nor (_34871_, _34837_, _34612_);
  nor (_34872_, _34871_, _34870_);
  and (_34873_, _34872_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34874_, _34837_, _32050_);
  nor (_34875_, _34837_, _34595_);
  nor (_34876_, _34875_, _34874_);
  and (_34877_, _34876_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_34878_, _34872_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_34879_, _34878_, _34873_);
  and (_34880_, _34879_, _34877_);
  nor (_34881_, _34880_, _34873_);
  not (_34882_, _34881_);
  nor (_34883_, _34868_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_34884_, _34883_, _34869_);
  and (_34885_, _34884_, _34882_);
  nor (_34886_, _34885_, _34869_);
  nor (_34887_, _34886_, _34865_);
  or (_34888_, _34887_, _34864_);
  or (_34889_, _34859_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34890_, _34889_, _34860_);
  nand (_34891_, _34890_, _34888_);
  and (_34892_, _34891_, _34860_);
  nor (_34893_, _34892_, _34856_);
  or (_34894_, _34893_, _34855_);
  and (_34895_, _34894_, _34851_);
  nor (_34896_, _34895_, _34849_);
  not (_34897_, _34896_);
  nand (_34898_, _34897_, _34845_);
  and (_34899_, _34898_, _34843_);
  nor (_34900_, _34899_, _30550_);
  and (_34901_, _34900_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_34902_, _34901_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34903_, _34902_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_34904_, _34903_, _34841_);
  and (_34905_, _34904_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34906_, _34899_, _30550_);
  and (_34907_, _34906_, _30556_);
  and (_34908_, _34907_, _30561_);
  and (_34909_, _34908_, _30546_);
  and (_34910_, _34909_, _30567_);
  and (_34911_, _34910_, _34840_);
  nor (_34912_, _34911_, _34905_);
  nor (_34913_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_34914_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_34915_, _34914_, _34913_);
  nor (_34916_, _34915_, _34912_);
  nor (_34917_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_34918_, _34840_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_34919_, _34918_, _34917_);
  nand (_34920_, _34919_, _34916_);
  or (_34921_, _34920_, _30578_);
  nand (_34922_, _34920_, _30578_);
  not (_34923_, _30363_);
  and (_34924_, _34828_, _34923_);
  and (_34925_, _34924_, _34749_);
  and (_34926_, _34925_, _34781_);
  nor (_34927_, _34926_, _30365_);
  nor (_34928_, _34927_, _34834_);
  and (_34929_, _30274_, _30252_);
  nor (_34930_, _34929_, _34791_);
  not (_34931_, _34930_);
  and (_34932_, _34931_, _34837_);
  nor (_34933_, _34932_, _34928_);
  and (_34934_, _34933_, _34922_);
  and (_34935_, _34934_, _34921_);
  nor (_34936_, _34832_, _27126_);
  not (_34937_, _34929_);
  nor (_34938_, _34937_, _30629_);
  and (_34939_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34940_, _34939_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34941_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34942_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34943_, _34942_, _34941_);
  and (_34944_, _34943_, _34940_);
  and (_34945_, _34944_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_34946_, _34945_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_34947_, _34946_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34948_, _34947_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_34949_, _34948_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34950_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_34951_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_34952_, _34951_, _30578_);
  or (_34953_, _34951_, _30578_);
  and (_34954_, _34953_, _34952_);
  and (_34955_, _34932_, _34928_);
  and (_34956_, _34955_, _34954_);
  not (_34957_, _34200_);
  and (_34958_, _30347_, _30215_);
  nor (_34959_, _34958_, _34272_);
  and (_34960_, _34959_, _34957_);
  or (_34961_, _34960_, _29998_);
  nor (_34962_, _30211_, _30113_);
  and (_34963_, _34962_, _30213_);
  nand (_34964_, _34963_, _30251_);
  or (_34965_, _30365_, _34964_);
  and (_34966_, _34965_, _34961_);
  not (_34967_, _31955_);
  and (_34968_, _34959_, _34967_);
  and (_34969_, _34968_, _31967_);
  or (_34970_, _34969_, _29998_);
  nor (_34971_, _34830_, _30361_);
  and (_34972_, _34971_, _34970_);
  nor (_34973_, _31955_, _30368_);
  nor (_34974_, _34973_, _29998_);
  nor (_34975_, _34974_, _34927_);
  and (_34976_, _34975_, _34972_);
  and (_34977_, _34976_, _34966_);
  and (_34978_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_34979_, _34833_, _31994_);
  or (_34980_, _34979_, _34978_);
  or (_34981_, _34980_, _34956_);
  nor (_34982_, _34981_, _34938_);
  nand (_34983_, _34982_, _34804_);
  or (_34984_, _34983_, _34936_);
  or (_34985_, _34984_, _34935_);
  and (_30881_, _34985_, _34827_);
  and (_34986_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _36029_);
  and (_34987_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_34988_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_34989_, _30002_, _34988_);
  not (_34990_, _34989_);
  not (_34991_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_34992_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_34993_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_34994_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_34995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_34996_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_34997_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_34998_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_34999_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_35000_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_35001_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_35002_, _35001_, _35000_);
  and (_35003_, _35002_, _34999_);
  and (_35004_, _35003_, _34998_);
  and (_35005_, _35004_, _34997_);
  and (_35006_, _35005_, _34996_);
  and (_35007_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_35008_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_35009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_35010_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_35011_, _35010_, _35008_);
  and (_35012_, _35011_, _35009_);
  nor (_35013_, _35012_, _35008_);
  nor (_35014_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_35015_, _35014_, _35007_);
  not (_35016_, _35015_);
  nor (_35017_, _35016_, _35013_);
  nor (_35018_, _35017_, _35007_);
  and (_35019_, _35018_, _35006_);
  and (_35020_, _35019_, _34995_);
  and (_35021_, _35020_, _34994_);
  and (_35022_, _35021_, _34993_);
  and (_35023_, _35022_, _34992_);
  and (_35024_, _35023_, _34991_);
  nor (_35025_, _35024_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_35026_, _35024_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_35027_, _35026_, _35025_);
  nor (_35028_, _35023_, _34991_);
  nor (_35029_, _35028_, _35024_);
  not (_35030_, _35029_);
  nor (_35031_, _35022_, _34992_);
  nor (_35032_, _35031_, _35023_);
  not (_35033_, _35032_);
  nor (_35034_, _35021_, _34993_);
  or (_35035_, _35034_, _35022_);
  nor (_35036_, _35020_, _34994_);
  nor (_35037_, _35036_, _35021_);
  not (_35038_, _35037_);
  nor (_35039_, _35019_, _34995_);
  or (_35040_, _35039_, _35020_);
  and (_35041_, _35018_, _35005_);
  nor (_35042_, _35041_, _34996_);
  nor (_35043_, _35042_, _35019_);
  not (_35044_, _35043_);
  and (_35045_, _35018_, _35003_);
  nor (_35046_, _35045_, _34998_);
  and (_35047_, _35018_, _35004_);
  nor (_35048_, _35047_, _35046_);
  not (_35049_, _35048_);
  and (_35050_, _35018_, _35002_);
  nor (_35051_, _35050_, _34999_);
  nor (_35052_, _35051_, _35045_);
  not (_35053_, _35052_);
  and (_35054_, _35018_, _35001_);
  nor (_35055_, _35054_, _35000_);
  nor (_35056_, _35055_, _35050_);
  not (_35057_, _35056_);
  not (_35058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_35059_, _35018_, _35058_);
  nor (_35060_, _35018_, _35058_);
  nor (_35061_, _35060_, _35059_);
  not (_35062_, _35061_);
  and (_35063_, _34036_, _34014_);
  or (_35064_, _34087_, _34055_);
  nor (_35065_, _35064_, _35063_);
  and (_35066_, _34065_, _34014_);
  nor (_35067_, _35066_, _34003_);
  not (_35068_, _34065_);
  nor (_35069_, _34081_, _34046_);
  and (_35070_, _35069_, _35068_);
  nor (_35071_, _35070_, _35067_);
  not (_35072_, _35071_);
  and (_35073_, _35072_, _34080_);
  and (_35074_, _35073_, _35065_);
  not (_35075_, _34027_);
  and (_35076_, _34007_, _34073_);
  and (_35077_, _34024_, _30037_);
  nor (_35078_, _35077_, _35076_);
  nor (_35079_, _35078_, _35075_);
  not (_35080_, _34084_);
  and (_35081_, _34044_, _34007_);
  nor (_35082_, _34075_, _35081_);
  nor (_35083_, _35082_, _35080_);
  nor (_35084_, _35083_, _35079_);
  and (_35085_, _34065_, _34018_);
  and (_35086_, _34053_, _34007_);
  and (_35087_, _35086_, _34003_);
  nor (_35088_, _35087_, _35085_);
  and (_35089_, _35088_, _35084_);
  or (_35090_, _34081_, _34056_);
  and (_35091_, _35090_, _34086_);
  nor (_35092_, _35091_, _34093_);
  nor (_35093_, _34081_, _35076_);
  nor (_35094_, _35093_, _30154_);
  not (_35095_, _34003_);
  and (_35096_, _34024_, _34051_);
  nor (_35097_, _35096_, _34036_);
  nor (_35098_, _35097_, _35095_);
  nor (_35099_, _35098_, _35094_);
  and (_35100_, _35099_, _35092_);
  and (_35101_, _35100_, _35089_);
  and (_35102_, _34056_, _34003_);
  not (_35103_, _35102_);
  and (_35104_, _35096_, _34086_);
  and (_35105_, _34081_, _34014_);
  nor (_35106_, _35105_, _35104_);
  and (_35107_, _35106_, _35103_);
  not (_35108_, _34086_);
  and (_35109_, _34024_, _34035_);
  nor (_35110_, _35109_, _34065_);
  nor (_35111_, _35110_, _35108_);
  and (_35112_, _34024_, _34073_);
  nor (_35113_, _35112_, _33996_);
  nor (_35114_, _35113_, _35108_);
  nor (_35115_, _35114_, _35111_);
  and (_35116_, _34027_, _35081_);
  and (_35117_, _34014_, _34068_);
  nor (_35118_, _35117_, _35116_);
  and (_35119_, _35118_, _35115_);
  and (_35120_, _35119_, _35107_);
  and (_35121_, _35120_, _35101_);
  and (_35122_, _34015_, _33998_);
  not (_35123_, _35122_);
  and (_35124_, _34086_, _34036_);
  and (_35125_, _34064_, _34044_);
  and (_35126_, _35125_, _34018_);
  nor (_35127_, _35126_, _35124_);
  not (_35128_, _35127_);
  nor (_35129_, _30131_, _30109_);
  not (_35130_, _35129_);
  and (_35131_, _34064_, _33995_);
  and (_35132_, _35131_, _34040_);
  and (_35133_, _34030_, _34007_);
  nor (_35134_, _35133_, _35132_);
  nor (_35135_, _35134_, _35130_);
  nor (_35136_, _35135_, _35128_);
  and (_35137_, _35136_, _35123_);
  nor (_35138_, _34091_, _34057_);
  and (_35139_, _34056_, _34010_);
  not (_35140_, _35139_);
  and (_35141_, _35131_, _34031_);
  nor (_35142_, _35141_, _34047_);
  and (_35143_, _35142_, _35140_);
  and (_35144_, _35143_, _35138_);
  not (_35145_, _35125_);
  nor (_35146_, _34084_, _34003_);
  nor (_35147_, _35146_, _35145_);
  nor (_35148_, _35129_, _34010_);
  and (_35149_, _35148_, _35075_);
  nor (_35150_, _35149_, _34038_);
  nor (_35151_, _35150_, _35147_);
  and (_35152_, _35151_, _35144_);
  and (_35153_, _35152_, _35137_);
  and (_35154_, _35153_, _35121_);
  and (_35158_, _35154_, _35074_);
  not (_35163_, _35158_);
  nor (_35171_, _35011_, _35009_);
  nor (_35177_, _35171_, _35012_);
  nand (_35181_, _35177_, _35163_);
  nor (_35192_, _35148_, _34038_);
  nor (_35203_, _35192_, _34069_);
  nand (_35207_, _35203_, _35092_);
  or (_35212_, _35207_, _35128_);
  and (_35220_, _34075_, _34018_);
  or (_35226_, _35116_, _35085_);
  nor (_35230_, _35226_, _35220_);
  nand (_35237_, _35230_, _35065_);
  or (_35238_, _35237_, _35212_);
  nor (_35248_, _35238_, _35158_);
  not (_35255_, _35248_);
  nor (_35263_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_35274_, _35263_, _35009_);
  and (_35285_, _35274_, _35255_);
  or (_35289_, _35177_, _35163_);
  and (_35300_, _35289_, _35181_);
  nand (_35311_, _35300_, _35285_);
  and (_35322_, _35311_, _35181_);
  not (_35333_, _35322_);
  and (_35341_, _35016_, _35013_);
  nor (_35348_, _35341_, _35017_);
  and (_35352_, _35348_, _35333_);
  and (_35358_, _35352_, _35062_);
  not (_35366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_35371_, _35059_, _35366_);
  or (_35375_, _35371_, _35054_);
  and (_35376_, _35375_, _35358_);
  and (_35377_, _35376_, _35057_);
  and (_35378_, _35377_, _35053_);
  and (_35379_, _35378_, _35049_);
  nor (_35380_, _35047_, _34997_);
  or (_35381_, _35380_, _35041_);
  and (_35382_, _35381_, _35379_);
  and (_35383_, _35382_, _35044_);
  and (_35384_, _35383_, _35040_);
  and (_35385_, _35384_, _35038_);
  and (_35386_, _35385_, _35035_);
  and (_35387_, _35386_, _35033_);
  and (_35388_, _35387_, _35030_);
  or (_35389_, _35388_, _35027_);
  nand (_35390_, _35388_, _35027_);
  and (_35391_, _35390_, _35389_);
  or (_35392_, _35391_, _34990_);
  or (_35393_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_35394_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_35395_, _35394_, _35393_);
  and (_35396_, _35395_, _35392_);
  or (_30883_, _35396_, _34987_);
  nor (_35397_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_30884_, _35397_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_30885_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _36029_);
  and (_35398_, \oc8051_top_1.oc8051_rom1.ea_int , _29999_);
  nand (_35399_, _35398_, _30002_);
  and (_30886_, _35399_, _30885_);
  and (_30888_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _36029_);
  nor (_35400_, _34808_, _31856_);
  or (_35401_, _35158_, _30026_);
  nor (_35402_, _35248_, _30019_);
  nand (_35403_, _35158_, _30026_);
  and (_35404_, _35403_, _35401_);
  nand (_35405_, _35404_, _35402_);
  and (_35406_, _35405_, _35401_);
  nor (_35407_, _35406_, _31856_);
  and (_35408_, _35407_, _30009_);
  nor (_35409_, _35407_, _30009_);
  nor (_35410_, _35409_, _35408_);
  nor (_35411_, _35410_, _35400_);
  and (_35412_, _30027_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_35413_, _35412_, _35400_);
  and (_35414_, _35413_, _35238_);
  or (_35415_, _35414_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_35416_, _35415_, _35411_);
  and (_30889_, _35416_, _36029_);
  not (_35417_, _30150_);
  and (_35418_, _30033_, _35417_);
  nor (_35419_, _30079_, _30057_);
  and (_35420_, _35419_, _35418_);
  not (_35421_, _30170_);
  and (_35422_, _30003_, _36029_);
  and (_35423_, _35422_, _30126_);
  and (_35424_, _35423_, _35421_);
  nor (_35425_, _30203_, _30105_);
  and (_35426_, _35425_, _35424_);
  and (_30892_, _35426_, _35420_);
  nor (_35427_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_35428_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_35429_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_30895_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _36029_);
  and (_35430_, _30895_, _35429_);
  or (_30893_, _35430_, _35428_);
  not (_35431_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_35432_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35433_, _35432_, _35431_);
  and (_35434_, _35432_, _35431_);
  nor (_35435_, _35434_, _35433_);
  not (_35436_, _35435_);
  and (_35437_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_35438_, _35437_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35439_, _35437_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_35440_, _35439_, _35438_);
  or (_35441_, _35440_, _35432_);
  and (_35442_, _35441_, _35436_);
  nor (_35443_, _35433_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_35444_, _35433_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_35445_, _35444_, _35443_);
  or (_35446_, _35438_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_30897_, _35446_, _36029_);
  and (_35447_, _30897_, _35445_);
  and (_30896_, _35447_, _35442_);
  not (_35448_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_35449_, _34808_, _35448_);
  and (_35450_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_35451_, _35449_);
  and (_35452_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_35453_, _35452_, _35450_);
  and (_30898_, _35453_, _36029_);
  and (_35454_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_35455_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_35456_, _35455_, _35454_);
  and (_30899_, _35456_, _36029_);
  and (_35457_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_35458_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35459_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _35458_);
  and (_35460_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_35461_, _35460_, _35457_);
  and (_30900_, _35461_, _36029_);
  and (_35462_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_35463_, _35462_, _35459_);
  and (_30901_, _35463_, _36029_);
  or (_35464_, _35458_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_30903_, _35464_, _36029_);
  not (_35465_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_35466_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_35467_, _35466_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_35468_, _35458_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_35469_, _35468_, _36029_);
  and (_30904_, _35469_, _35467_);
  or (_35470_, _35458_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_30905_, _35470_, _36029_);
  nor (_35471_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_35472_, _35471_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35473_, _35472_, _36029_);
  and (_35474_, _30895_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_30906_, _35474_, _35473_);
  and (_35475_, _35448_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_35476_, _35475_, _35472_);
  and (_30907_, _35476_, _36029_);
  nand (_35477_, _35472_, _30629_);
  or (_35478_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_35479_, _35478_, _36029_);
  and (_30908_, _35479_, _35477_);
  and (_30909_, _30395_, _31853_);
  or (_35480_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_35481_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_35482_, _34698_, _35481_);
  and (_35483_, _35482_, _36029_);
  and (_30941_, _35483_, _35480_);
  or (_35484_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_35485_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_35486_, _34698_, _35485_);
  and (_35487_, _35486_, _36029_);
  and (_30942_, _35487_, _35484_);
  or (_35488_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_35489_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _36029_);
  or (_35490_, _35489_, _00000_);
  and (_30943_, _35490_, _35488_);
  or (_35491_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_35492_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_35493_, _34698_, _35492_);
  and (_35494_, _35493_, _36029_);
  and (_30944_, _35494_, _35491_);
  or (_35495_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_35496_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_35497_, _34698_, _35496_);
  and (_35498_, _35497_, _36029_);
  and (_30945_, _35498_, _35495_);
  or (_35499_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_35500_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_35501_, _34698_, _35500_);
  and (_35502_, _35501_, _36029_);
  and (_30946_, _35502_, _35499_);
  or (_35503_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_35504_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_35505_, _34698_, _35504_);
  and (_35506_, _35505_, _36029_);
  and (_30947_, _35506_, _35503_);
  or (_35507_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_35508_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7], _36029_);
  or (_35509_, _35508_, _00000_);
  and (_30948_, _35509_, _35507_);
  or (_35510_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_35511_, _34698_, _30550_);
  and (_35512_, _35511_, _36029_);
  and (_30949_, _35512_, _35510_);
  or (_35513_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_35514_, _34698_, _30556_);
  and (_35515_, _35514_, _36029_);
  and (_30950_, _35515_, _35513_);
  or (_35516_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_35517_, _34698_, _30561_);
  and (_35518_, _35517_, _36029_);
  and (_30951_, _35518_, _35516_);
  or (_35519_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_35520_, _34698_, _30546_);
  and (_35521_, _35520_, _36029_);
  and (_30952_, _35521_, _35519_);
  or (_35522_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_35523_, _34698_, _30567_);
  and (_35524_, _35523_, _36029_);
  and (_30953_, _35524_, _35522_);
  or (_35525_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_35526_, _34698_, _30542_);
  and (_35527_, _35526_, _36029_);
  and (_30954_, _35527_, _35525_);
  or (_35528_, _34698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_35529_, _34698_, _30573_);
  and (_35530_, _35529_, _36029_);
  and (_30956_, _35530_, _35528_);
  or (_35531_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_35532_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _36029_);
  or (_35533_, _35532_, _00000_);
  and (_30960_, _35533_, _35531_);
  or (_35534_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_35535_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _36029_);
  or (_35536_, _35535_, _00000_);
  and (_30961_, _35536_, _35534_);
  or (_35537_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_35538_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _36029_);
  or (_35539_, _35538_, _00000_);
  and (_30962_, _35539_, _35537_);
  or (_35540_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_35541_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _36029_);
  or (_35542_, _35541_, _00000_);
  and (_30963_, _35542_, _35540_);
  or (_35543_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_35544_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _36029_);
  or (_35545_, _35544_, _00000_);
  and (_30964_, _35545_, _35543_);
  or (_35546_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_35547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _36029_);
  or (_35548_, _35547_, _00000_);
  and (_30965_, _35548_, _35546_);
  or (_35549_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_35550_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _36029_);
  or (_35551_, _35550_, _00000_);
  and (_30966_, _35551_, _35549_);
  or (_35552_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_35553_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _36029_);
  or (_35554_, _35553_, _00000_);
  and (_30967_, _35554_, _35552_);
  or (_35555_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_35556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _36029_);
  or (_35557_, _35556_, _00000_);
  and (_30968_, _35557_, _35555_);
  or (_35558_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_35559_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _36029_);
  or (_35560_, _35559_, _00000_);
  and (_30970_, _35560_, _35558_);
  or (_35561_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_35562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _36029_);
  or (_35563_, _35562_, _00000_);
  and (_30971_, _35563_, _35561_);
  or (_35564_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_35565_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _36029_);
  or (_35566_, _35565_, _00000_);
  and (_30972_, _35566_, _35564_);
  or (_35567_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_35568_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _36029_);
  or (_35569_, _35568_, _00000_);
  and (_30973_, _35569_, _35567_);
  or (_35570_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_35571_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _36029_);
  or (_35572_, _35571_, _00000_);
  and (_30974_, _35572_, _35570_);
  or (_35573_, _34702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_35574_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _36029_);
  or (_35575_, _35574_, _00000_);
  and (_30975_, _35575_, _35573_);
  and (_35576_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_35577_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_35578_, _35577_, _35576_);
  and (_31153_, _35578_, _36029_);
  and (_35579_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35580_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_35581_, _35580_, _35579_);
  and (_31154_, _35581_, _36029_);
  and (_35582_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_35583_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_35584_, _35583_, _35582_);
  and (_31155_, _35584_, _36029_);
  and (_35585_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_35586_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_35587_, _35586_, _35585_);
  and (_31156_, _35587_, _36029_);
  and (_35588_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_35589_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_35590_, _35589_, _35449_);
  or (_35591_, _35590_, _35588_);
  and (_31157_, _35591_, _36029_);
  and (_35592_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_35593_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_35594_, _35593_, _35592_);
  and (_31158_, _35594_, _36029_);
  and (_35595_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_35596_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_35597_, _35596_, _35595_);
  and (_31159_, _35597_, _36029_);
  and (_35598_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_35599_, _35449_, _35429_);
  or (_35600_, _35599_, _35598_);
  and (_31161_, _35600_, _36029_);
  and (_35601_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_35602_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_35603_, _35602_, _35601_);
  and (_31162_, _35603_, _36029_);
  and (_35604_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_35605_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_35606_, _35605_, _35604_);
  and (_31163_, _35606_, _36029_);
  and (_35607_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_35608_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_35609_, _35608_, _35607_);
  and (_31164_, _35609_, _36029_);
  and (_35610_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_35611_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_35612_, _35611_, _35610_);
  and (_31165_, _35612_, _36029_);
  and (_35613_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_35614_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_35615_, _35614_, _35613_);
  and (_31166_, _35615_, _36029_);
  and (_35616_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_35617_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_35618_, _35617_, _35616_);
  and (_31167_, _35618_, _36029_);
  and (_35619_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_35620_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_35621_, _35620_, _35619_);
  and (_31168_, _35621_, _36029_);
  and (_35622_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_35623_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_35624_, _35623_, _35622_);
  and (_31169_, _35624_, _36029_);
  and (_35625_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_35626_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_35627_, _35626_, _35625_);
  and (_31170_, _35627_, _36029_);
  and (_35628_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_35629_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_35630_, _35629_, _35628_);
  and (_31172_, _35630_, _36029_);
  and (_35631_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_35632_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_35633_, _35632_, _35631_);
  and (_31173_, _35633_, _36029_);
  and (_35634_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_35635_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_35636_, _35635_, _35634_);
  and (_31174_, _35636_, _36029_);
  and (_35637_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_35638_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_35639_, _35638_, _35637_);
  and (_31175_, _35639_, _36029_);
  and (_35640_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_35641_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_35642_, _35641_, _35640_);
  and (_31176_, _35642_, _36029_);
  and (_35643_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_35644_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_35645_, _35644_, _35643_);
  and (_31177_, _35645_, _36029_);
  and (_35646_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_35647_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_35648_, _35647_, _35646_);
  and (_31178_, _35648_, _36029_);
  and (_35649_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_35650_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_35651_, _35650_, _35649_);
  and (_31179_, _35651_, _36029_);
  and (_35652_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_35653_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_35654_, _35653_, _35652_);
  and (_31180_, _35654_, _36029_);
  and (_35655_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_35656_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_35657_, _35656_, _35655_);
  and (_31181_, _35657_, _36029_);
  and (_35658_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_35659_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_35660_, _35659_, _35658_);
  and (_31183_, _35660_, _36029_);
  and (_35661_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_35662_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_35663_, _35662_, _35661_);
  and (_31184_, _35663_, _36029_);
  and (_35664_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_35665_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_35666_, _35665_, _35664_);
  and (_31185_, _35666_, _36029_);
  and (_35667_, _35449_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_35668_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_35669_, _35668_, _35667_);
  and (_31186_, _35669_, _36029_);
  nor (_31187_, _30211_, rst);
  nor (_31188_, _30113_, rst);
  nor (_31189_, _30135_, rst);
  nor (_31190_, _31892_, rst);
  nor (_31191_, _32034_, rst);
  nor (_31193_, _32179_, rst);
  nor (_31194_, _31911_, rst);
  nor (_31195_, _32091_, rst);
  nor (_31196_, _32221_, rst);
  nor (_31197_, _31946_, rst);
  nor (_31199_, _32121_, rst);
  and (_31215_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _36029_);
  and (_31216_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36029_);
  and (_31217_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _36029_);
  and (_31218_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _36029_);
  and (_31220_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36029_);
  and (_31221_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _36029_);
  and (_31222_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _36029_);
  or (_35670_, _34804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_35671_, _35670_, _36029_);
  and (_35672_, _34930_, _34928_);
  and (_35673_, _35672_, _34837_);
  or (_35674_, _35673_, _34929_);
  and (_35675_, _35674_, _28305_);
  or (_35676_, _34876_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_35677_, _34877_);
  and (_35678_, _34933_, _35677_);
  and (_35679_, _35678_, _35676_);
  and (_35680_, _34955_, _32051_);
  and (_35681_, _34833_, _34595_);
  and (_35682_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_35683_, _35682_, _35681_);
  or (_35684_, _35683_, _35680_);
  nor (_35685_, _35684_, _35679_);
  nand (_35686_, _35685_, _34804_);
  or (_35687_, _35686_, _35675_);
  and (_31223_, _35687_, _35671_);
  or (_35688_, _34804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_35689_, _35688_, _36029_);
  and (_35690_, _35674_, _28950_);
  or (_35691_, _34879_, _34877_);
  not (_35692_, _34880_);
  and (_35693_, _34933_, _35692_);
  and (_35694_, _35693_, _35691_);
  and (_35695_, _34955_, _32167_);
  and (_35696_, _34833_, _34612_);
  and (_35697_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_35698_, _35697_, _35696_);
  or (_35699_, _35698_, _35695_);
  nor (_35700_, _35699_, _35694_);
  nand (_35701_, _35700_, _34804_);
  or (_35702_, _35701_, _35690_);
  and (_31224_, _35702_, _35689_);
  not (_35703_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_35704_, _34808_, _35703_);
  and (_35705_, _34808_, _35703_);
  nor (_35706_, _35705_, _35704_);
  or (_35707_, _35706_, _34804_);
  and (_35708_, _35707_, _36029_);
  and (_35709_, _35674_, _29595_);
  or (_35710_, _34884_, _34882_);
  not (_35711_, _34885_);
  and (_35712_, _34933_, _35711_);
  and (_35713_, _35712_, _35710_);
  and (_35714_, _34955_, _31873_);
  and (_35715_, _34833_, _34629_);
  and (_35716_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_35717_, _35716_, _35715_);
  or (_35718_, _35717_, _35714_);
  nor (_35719_, _35718_, _35713_);
  nand (_35720_, _35719_, _34804_);
  or (_35721_, _35720_, _35709_);
  and (_31225_, _35721_, _35708_);
  and (_35722_, _35704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35723_, _35704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35724_, _35723_, _35722_);
  or (_35725_, _35724_, _34804_);
  and (_35726_, _35725_, _36029_);
  and (_35727_, _35674_, _29761_);
  or (_35728_, _34865_, _34864_);
  or (_35729_, _35728_, _34886_);
  nand (_35730_, _35728_, _34886_);
  and (_35731_, _35730_, _34933_);
  and (_35732_, _35731_, _35729_);
  and (_35733_, _34955_, _32076_);
  and (_35734_, _34833_, _34646_);
  and (_35735_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_35736_, _35735_, _35734_);
  or (_35737_, _35736_, _35733_);
  nor (_35738_, _35737_, _35732_);
  nand (_35739_, _35738_, _34804_);
  or (_35740_, _35739_, _35727_);
  and (_31226_, _35740_, _35726_);
  and (_35741_, _34811_, _34809_);
  nor (_35742_, _35722_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_35743_, _35742_, _35741_);
  or (_35744_, _35743_, _34804_);
  and (_35745_, _35744_, _36029_);
  and (_35746_, _35674_, _29831_);
  or (_35747_, _34890_, _34888_);
  and (_35748_, _34933_, _34891_);
  and (_35749_, _35748_, _35747_);
  and (_35750_, _34955_, _32206_);
  and (_35751_, _34833_, _34663_);
  and (_35752_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_35753_, _35752_, _35751_);
  or (_35754_, _35753_, _35750_);
  nor (_35755_, _35754_, _35749_);
  nand (_35756_, _35755_, _34804_);
  or (_35757_, _35756_, _35746_);
  and (_31227_, _35757_, _35745_);
  nor (_35758_, _35741_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_35759_, _35758_, _34813_);
  or (_35760_, _35759_, _34804_);
  and (_35761_, _35760_, _36029_);
  and (_35762_, _35674_, _29904_);
  or (_35763_, _34855_, _34856_);
  nand (_35764_, _35763_, _34892_);
  or (_35765_, _35763_, _34892_);
  and (_35766_, _35765_, _34933_);
  and (_35767_, _35766_, _35764_);
  and (_35768_, _34955_, _31933_);
  and (_35769_, _34833_, _34680_);
  and (_35770_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_35771_, _35770_, _35769_);
  or (_35772_, _35771_, _35768_);
  nor (_35773_, _35772_, _35767_);
  nand (_35774_, _35773_, _34804_);
  or (_35775_, _35774_, _35762_);
  and (_31228_, _35775_, _35761_);
  nor (_35776_, _34813_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35777_, _34813_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_35778_, _35777_, _35776_);
  or (_35779_, _35778_, _34804_);
  and (_35780_, _35779_, _36029_);
  and (_35781_, _35674_, _29977_);
  or (_35782_, _34894_, _34851_);
  not (_35783_, _34895_);
  and (_35784_, _34933_, _35783_);
  and (_35785_, _35784_, _35782_);
  and (_35786_, _34833_, _34697_);
  and (_35787_, _34955_, _32138_);
  and (_35788_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_35789_, _35788_, _35787_);
  nor (_35790_, _35789_, _35786_);
  nand (_35791_, _35790_, _34804_);
  or (_35792_, _35791_, _35785_);
  or (_35793_, _35792_, _35781_);
  and (_31229_, _35793_, _35780_);
  nor (_35794_, _35777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35795_, _35777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_35796_, _35795_, _35794_);
  or (_35797_, _35796_, _34804_);
  and (_35798_, _35797_, _36029_);
  and (_35799_, _35674_, _27137_);
  or (_35800_, _34897_, _34845_);
  and (_35801_, _34933_, _34898_);
  and (_35802_, _35801_, _35800_);
  nand (_35803_, _34955_, _31994_);
  and (_35804_, _34833_, _34578_);
  and (_35805_, _30278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_35806_, _35805_, _35804_);
  and (_35807_, _35806_, _35803_);
  nand (_35808_, _35807_, _34804_);
  or (_35809_, _35808_, _35802_);
  or (_35810_, _35809_, _35799_);
  and (_31231_, _35810_, _35798_);
  or (_35811_, _35795_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_35812_, _34815_, _34813_);
  and (_35813_, _35812_, _35811_);
  or (_35814_, _35813_, _34804_);
  and (_35815_, _35814_, _36029_);
  nor (_35816_, _34832_, _28302_);
  nor (_35817_, _34937_, _30667_);
  nor (_35818_, _34899_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35819_, _34899_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_35820_, _35819_, _35818_);
  or (_35821_, _35820_, _34841_);
  nand (_35822_, _35820_, _34841_);
  and (_35823_, _35822_, _34933_);
  and (_35824_, _35823_, _35821_);
  nand (_35825_, _34955_, _33995_);
  and (_35826_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35827_, _34833_, _32051_);
  nor (_35828_, _35827_, _35826_);
  and (_35829_, _35828_, _35825_);
  nand (_35830_, _35829_, _34804_);
  or (_35831_, _35830_, _35824_);
  or (_35832_, _35831_, _35817_);
  or (_35833_, _35832_, _35816_);
  and (_31232_, _35833_, _35815_);
  nand (_35834_, _35812_, _34996_);
  or (_35835_, _35812_, _34996_);
  and (_35836_, _35835_, _35834_);
  or (_35837_, _35836_, _34804_);
  and (_35838_, _35837_, _36029_);
  nor (_35839_, _34832_, _28939_);
  and (_35840_, _34906_, _34840_);
  and (_35841_, _34900_, _34841_);
  nor (_35842_, _35841_, _35840_);
  and (_35843_, _35842_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_35844_, _35842_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_35845_, _35844_, _35843_);
  and (_35846_, _35845_, _34933_);
  not (_35847_, _34804_);
  nor (_35848_, _34937_, _30698_);
  and (_35849_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_35850_, _34833_, _32167_);
  and (_35851_, _34955_, _34063_);
  or (_35852_, _35851_, _35850_);
  or (_35853_, _35852_, _35849_);
  or (_35854_, _35853_, _35848_);
  or (_35855_, _35854_, _35847_);
  or (_35856_, _35855_, _35846_);
  or (_35857_, _35856_, _35839_);
  and (_31233_, _35857_, _35838_);
  and (_35858_, _34812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35859_, _35858_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35860_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35861_, _35860_, _35859_);
  and (_35862_, _35861_, _34809_);
  nor (_35863_, _35862_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35864_, _35862_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_35865_, _35864_, _35863_);
  or (_35866_, _35865_, _34804_);
  and (_35867_, _35866_, _36029_);
  nor (_35868_, _34832_, _29584_);
  and (_35869_, _34907_, _34840_);
  and (_35870_, _34901_, _34841_);
  nor (_35871_, _35870_, _35869_);
  nor (_35872_, _35871_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_35873_, _35871_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_35874_, _35873_, _35872_);
  and (_35875_, _35874_, _34933_);
  or (_35876_, _34937_, _30728_);
  and (_35877_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35878_, _34833_, _31873_);
  and (_35879_, _34955_, _34006_);
  or (_35880_, _35879_, _35878_);
  nor (_35881_, _35880_, _35877_);
  and (_35882_, _35881_, _35876_);
  nand (_35883_, _35882_, _34804_);
  or (_35884_, _35883_, _35875_);
  or (_35885_, _35884_, _35868_);
  and (_31234_, _35885_, _35867_);
  nor (_35886_, _35864_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35887_, _35864_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_35888_, _35887_, _35886_);
  or (_35889_, _35888_, _34804_);
  and (_35890_, _35889_, _36029_);
  nor (_35891_, _34832_, _29760_);
  and (_35892_, _34902_, _34841_);
  and (_35893_, _34908_, _34840_);
  nor (_35894_, _35893_, _35892_);
  nand (_35895_, _35894_, _30546_);
  or (_35896_, _35894_, _30546_);
  and (_35897_, _35896_, _34933_);
  and (_35898_, _35897_, _35895_);
  or (_35899_, _34937_, _30757_);
  and (_35900_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_35901_, _34947_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_35902_, _35901_, _34948_);
  and (_35903_, _35902_, _34955_);
  or (_35904_, _35903_, _35900_);
  and (_35905_, _34833_, _32076_);
  nor (_35906_, _35905_, _35904_);
  and (_35907_, _35906_, _35899_);
  nand (_35908_, _35907_, _34804_);
  or (_35909_, _35908_, _35898_);
  or (_35910_, _35909_, _35891_);
  and (_31235_, _35910_, _35890_);
  and (_35911_, _35887_, _34993_);
  nor (_35912_, _35887_, _34993_);
  nor (_35913_, _35912_, _35911_);
  nor (_35914_, _35913_, _34804_);
  and (_35915_, _34909_, _34840_);
  nor (_35916_, _35915_, _34904_);
  nor (_35917_, _35916_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_35918_, _35916_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_35919_, _35918_, _35917_);
  and (_35920_, _35919_, _34933_);
  nor (_35921_, _34937_, _30815_);
  and (_35922_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35923_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_35924_, _35923_, _35922_);
  and (_35925_, _34944_, _35924_);
  and (_35926_, _35925_, _30567_);
  nor (_35927_, _35925_, _30567_);
  or (_35928_, _35927_, _35926_);
  and (_35929_, _35928_, _34955_);
  and (_35930_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_35931_, _34833_, _32206_);
  or (_35932_, _35931_, _35930_);
  or (_35933_, _35932_, _35929_);
  or (_35934_, _35933_, _35921_);
  or (_35935_, _35934_, _35920_);
  nor (_35936_, _30362_, _29830_);
  or (_35937_, _35936_, _35935_);
  and (_35938_, _35937_, _34804_);
  or (_35939_, _35938_, _35914_);
  and (_31236_, _35939_, _36029_);
  nor (_35940_, _34820_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_35941_, _35940_, _34821_);
  or (_35942_, _35941_, _34804_);
  and (_35943_, _35942_, _36029_);
  nand (_35944_, _34912_, _30542_);
  or (_35945_, _34912_, _30542_);
  and (_35946_, _35945_, _34933_);
  and (_35947_, _35946_, _35944_);
  nor (_35948_, _34832_, _29903_);
  or (_35949_, _34937_, _30850_);
  and (_35950_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_35951_, _34833_, _31933_);
  nor (_35952_, _34949_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_35953_, _35952_, _34950_);
  and (_35954_, _35953_, _34955_);
  or (_35955_, _35954_, _35951_);
  nor (_35956_, _35955_, _35950_);
  and (_35957_, _35956_, _35949_);
  nand (_35958_, _35957_, _34804_);
  or (_35959_, _35958_, _35948_);
  or (_35960_, _35959_, _35947_);
  and (_31237_, _35960_, _35943_);
  nor (_35961_, _34821_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_35962_, _35961_, _34822_);
  or (_35963_, _35962_, _34804_);
  and (_35964_, _35963_, _36029_);
  nand (_35965_, _34916_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_35966_, _34916_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_35967_, _35966_, _34933_);
  and (_35968_, _35967_, _35965_);
  nor (_35969_, _34832_, _29976_);
  nor (_35970_, _34937_, _30914_);
  and (_35971_, _34977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_35972_, _34833_, _32138_);
  or (_35973_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_35974_, _35973_, _34951_);
  and (_35975_, _35974_, _34955_);
  or (_35976_, _35975_, _35972_);
  or (_35977_, _35976_, _35971_);
  nor (_35978_, _35977_, _35970_);
  nand (_35979_, _35978_, _34804_);
  or (_35980_, _35979_, _35969_);
  or (_35981_, _35980_, _35968_);
  and (_31238_, _35981_, _35964_);
  and (_35982_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_35983_, _35274_, _35255_);
  nor (_35984_, _35983_, _35285_);
  or (_35985_, _35984_, _34990_);
  or (_35986_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35987_, _35986_, _35394_);
  and (_35988_, _35987_, _35985_);
  or (_31239_, _35988_, _35982_);
  or (_35989_, _35300_, _35285_);
  and (_35990_, _35989_, _35311_);
  or (_35991_, _35990_, _34990_);
  or (_35992_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_35993_, _35992_, _35394_);
  and (_35994_, _35993_, _35991_);
  and (_35995_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_31240_, _35995_, _35994_);
  and (_35996_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_35997_, _35348_, _35333_);
  nor (_35998_, _35997_, _35352_);
  or (_35999_, _35998_, _34990_);
  or (_36000_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_36001_, _36000_, _35394_);
  and (_36002_, _36001_, _35999_);
  or (_31242_, _36002_, _35996_);
  and (_36003_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_36004_, _35352_, _35062_);
  nor (_36005_, _36004_, _35358_);
  or (_36006_, _36005_, _34990_);
  or (_36007_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_36009_, _36007_, _35394_);
  and (_36011_, _36009_, _36006_);
  or (_31243_, _36011_, _36003_);
  and (_36014_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_36016_, _35375_, _35358_);
  nor (_36018_, _36016_, _35376_);
  or (_36020_, _36018_, _34990_);
  or (_36021_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_36022_, _36021_, _35394_);
  and (_36023_, _36022_, _36020_);
  or (_31244_, _36023_, _36014_);
  and (_36024_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_36025_, _35376_, _35057_);
  nor (_36027_, _36025_, _35377_);
  or (_36028_, _36027_, _34990_);
  or (_36030_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_36031_, _36030_, _35394_);
  and (_36032_, _36031_, _36028_);
  or (_31245_, _36032_, _36024_);
  nor (_36034_, _35377_, _35053_);
  nor (_36035_, _36034_, _35378_);
  or (_36037_, _36035_, _34990_);
  or (_36038_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_36039_, _36038_, _35394_);
  and (_36041_, _36039_, _36037_);
  and (_36042_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_31246_, _36042_, _36041_);
  nor (_36044_, _35378_, _35049_);
  nor (_36045_, _36044_, _35379_);
  or (_36046_, _36045_, _34990_);
  or (_36048_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_36049_, _36048_, _35394_);
  and (_36050_, _36049_, _36046_);
  and (_36052_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_31247_, _36052_, _36050_);
  and (_36053_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_36055_, _35381_, _35379_);
  nor (_36056_, _36055_, _35382_);
  or (_36057_, _36056_, _34990_);
  or (_36058_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_36059_, _36058_, _35394_);
  and (_36060_, _36059_, _36057_);
  or (_31248_, _36060_, _36053_);
  and (_36061_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_36062_, _35382_, _35044_);
  nor (_36063_, _36062_, _35383_);
  or (_36064_, _36063_, _34990_);
  or (_36065_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_36066_, _36065_, _35394_);
  and (_36067_, _36066_, _36064_);
  or (_31249_, _36067_, _36061_);
  or (_36068_, _35383_, _35040_);
  nor (_36069_, _35384_, _34990_);
  and (_36070_, _36069_, _36068_);
  nor (_36071_, _34989_, _30561_);
  or (_36072_, _36071_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_36073_, _36072_, _36070_);
  or (_36075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _29999_);
  and (_36076_, _36075_, _36029_);
  and (_31250_, _36076_, _36073_);
  nor (_36078_, _35384_, _35038_);
  nor (_36079_, _36078_, _35385_);
  or (_36081_, _36079_, _34990_);
  or (_36082_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_36083_, _36082_, _35394_);
  and (_36085_, _36083_, _36081_);
  and (_36086_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_31251_, _36086_, _36085_);
  nor (_36088_, _35385_, _35035_);
  nor (_36089_, _36088_, _35386_);
  or (_36090_, _36089_, _34990_);
  or (_36092_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_36093_, _36092_, _35394_);
  and (_36094_, _36093_, _36090_);
  and (_36096_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_31253_, _36096_, _36094_);
  nor (_36097_, _35386_, _35033_);
  nor (_36099_, _36097_, _35387_);
  or (_36100_, _36099_, _34990_);
  or (_36101_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_36103_, _36101_, _35394_);
  and (_36104_, _36103_, _36100_);
  and (_36105_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_31254_, _36105_, _36104_);
  nor (_36106_, _35387_, _35030_);
  nor (_36107_, _36106_, _35388_);
  or (_36108_, _36107_, _34990_);
  or (_36109_, _34989_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_36110_, _36109_, _35394_);
  and (_36111_, _36110_, _36108_);
  and (_36112_, _34986_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_31255_, _36112_, _36111_);
  and (_31256_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _36029_);
  and (_31257_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _36029_);
  and (_31258_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _36029_);
  and (_31259_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _36029_);
  and (_31260_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _36029_);
  and (_31261_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _36029_);
  and (_31262_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _36029_);
  nor (_36113_, _35248_, _31856_);
  nand (_36114_, _36113_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_36116_, _36113_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_36117_, _36116_, _35394_);
  and (_31264_, _36117_, _36114_);
  or (_36119_, _35404_, _35402_);
  and (_36120_, _36119_, _35405_);
  or (_36122_, _36120_, _31856_);
  or (_36123_, _30002_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_36124_, _36123_, _35394_);
  and (_31265_, _36124_, _36122_);
  and (_36126_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_36127_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_36129_, _36127_, _30895_);
  or (_31281_, _36129_, _36126_);
  and (_00008_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00010_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00011_, _00010_, _30895_);
  or (_31282_, _00011_, _00008_);
  and (_00013_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00014_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00015_, _00014_, _30895_);
  or (_31283_, _00015_, _00013_);
  and (_00017_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00018_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00020_, _00018_, _30895_);
  or (_31284_, _00020_, _00017_);
  and (_00021_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00022_, _35589_, _30895_);
  or (_31286_, _00022_, _00021_);
  and (_00023_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00024_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00025_, _00024_, _30895_);
  or (_31287_, _00025_, _00023_);
  and (_00026_, _35427_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00027_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00028_, _00027_, _30895_);
  or (_31288_, _00028_, _00026_);
  and (_31289_, _35435_, _36029_);
  nor (_31290_, _35445_, rst);
  and (_31291_, _35441_, _36029_);
  and (_00029_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00030_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00031_, _00030_, _00029_);
  and (_31292_, _00031_, _36029_);
  and (_00032_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00034_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00035_, _00034_, _00032_);
  and (_31293_, _00035_, _36029_);
  and (_00037_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00038_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00040_, _00038_, _00037_);
  and (_31294_, _00040_, _36029_);
  and (_00041_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00043_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00044_, _00043_, _00041_);
  and (_31295_, _00044_, _36029_);
  and (_00046_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00047_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00048_, _00047_, _00046_);
  and (_31296_, _00048_, _36029_);
  and (_00050_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00051_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00053_, _00051_, _00050_);
  and (_31297_, _00053_, _36029_);
  and (_00054_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00056_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00057_, _00056_, _00054_);
  and (_31298_, _00057_, _36029_);
  and (_00059_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00060_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00061_, _00060_, _00059_);
  and (_31299_, _00061_, _36029_);
  and (_00062_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00063_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00064_, _00063_, _00062_);
  and (_31300_, _00064_, _36029_);
  and (_00065_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00066_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00067_, _00066_, _00065_);
  and (_31301_, _00067_, _36029_);
  and (_00068_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00069_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00070_, _00069_, _00068_);
  and (_31302_, _00070_, _36029_);
  and (_00071_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00072_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00073_, _00072_, _00071_);
  and (_31303_, _00073_, _36029_);
  and (_00074_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00076_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00077_, _00076_, _00074_);
  and (_31304_, _00077_, _36029_);
  and (_00079_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00080_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00082_, _00080_, _00079_);
  and (_31305_, _00082_, _36029_);
  and (_00083_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00085_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00086_, _00085_, _00083_);
  and (_31307_, _00086_, _36029_);
  and (_00088_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00089_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00090_, _00089_, _00088_);
  and (_31308_, _00090_, _36029_);
  and (_00092_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00093_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00095_, _00093_, _00092_);
  and (_31309_, _00095_, _36029_);
  and (_00096_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00098_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00099_, _00098_, _00096_);
  and (_31310_, _00099_, _36029_);
  and (_00101_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00102_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00103_, _00102_, _00101_);
  and (_31311_, _00103_, _36029_);
  and (_00104_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00105_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00106_, _00105_, _00104_);
  and (_31312_, _00106_, _36029_);
  and (_00107_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00108_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00109_, _00108_, _00107_);
  and (_31313_, _00109_, _36029_);
  and (_00110_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00111_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00112_, _00111_, _00110_);
  and (_31314_, _00112_, _36029_);
  and (_00113_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00114_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00115_, _00114_, _00113_);
  and (_31315_, _00115_, _36029_);
  and (_00116_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00118_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00119_, _00118_, _00116_);
  and (_31316_, _00119_, _36029_);
  and (_00121_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00122_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00124_, _00122_, _00121_);
  and (_31318_, _00124_, _36029_);
  and (_00125_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00127_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00128_, _00127_, _00125_);
  and (_31319_, _00128_, _36029_);
  and (_00130_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00131_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00132_, _00131_, _00130_);
  and (_31320_, _00132_, _36029_);
  and (_00134_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00135_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00137_, _00135_, _00134_);
  and (_31321_, _00137_, _36029_);
  and (_00138_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00140_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00141_, _00140_, _00138_);
  and (_31322_, _00141_, _36029_);
  and (_00143_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00144_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00145_, _00144_, _00143_);
  and (_31323_, _00145_, _36029_);
  and (_00146_, _35449_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00147_, _35451_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00148_, _00147_, _00146_);
  and (_31324_, _00148_, _36029_);
  and (_00149_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00150_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00151_, _00150_, _00149_);
  and (_31325_, _00151_, _36029_);
  and (_00152_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00153_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00154_, _00153_, _00152_);
  and (_31326_, _00154_, _36029_);
  and (_00155_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00156_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00157_, _00156_, _00155_);
  and (_31327_, _00157_, _36029_);
  and (_00158_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00160_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00161_, _00160_, _00158_);
  and (_31329_, _00161_, _36029_);
  and (_00163_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00164_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00166_, _00164_, _00163_);
  and (_31330_, _00166_, _36029_);
  and (_00167_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00169_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00170_, _00169_, _00167_);
  and (_31331_, _00170_, _36029_);
  and (_00172_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00173_, _35459_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00174_, _00173_, _00172_);
  and (_31332_, _00174_, _36029_);
  and (_00176_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00177_, _32034_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00179_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00180_, _00179_, _35458_);
  and (_00181_, _00180_, _00177_);
  or (_00183_, _00181_, _00176_);
  and (_31333_, _00183_, _36029_);
  and (_00184_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00186_, _32179_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00187_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00188_, _00187_, _35458_);
  and (_00189_, _00188_, _00186_);
  or (_00190_, _00189_, _00184_);
  and (_31334_, _00190_, _36029_);
  and (_00191_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00192_, _31911_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00193_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00194_, _00193_, _35458_);
  and (_00195_, _00194_, _00192_);
  or (_00196_, _00195_, _00191_);
  and (_31335_, _00196_, _36029_);
  and (_00197_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00198_, _32091_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00199_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00200_, _00199_, _35458_);
  and (_00201_, _00200_, _00198_);
  or (_00202_, _00201_, _00197_);
  and (_31336_, _00202_, _36029_);
  and (_00203_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00205_, _32221_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00206_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00208_, _00206_, _35458_);
  and (_00209_, _00208_, _00205_);
  or (_00210_, _00209_, _00203_);
  and (_31337_, _00210_, _36029_);
  and (_00212_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00213_, _31946_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00215_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00216_, _00215_, _35458_);
  and (_00217_, _00216_, _00213_);
  or (_00219_, _00217_, _00212_);
  and (_31338_, _00219_, _36029_);
  and (_00220_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00222_, _32121_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00223_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00224_, _00223_, _35458_);
  and (_00226_, _00224_, _00222_);
  or (_00227_, _00226_, _00220_);
  and (_31340_, _00227_, _36029_);
  and (_00229_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00230_, _32008_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00231_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00233_, _00231_, _35458_);
  and (_00234_, _00233_, _00230_);
  or (_00235_, _00234_, _00229_);
  and (_31341_, _00235_, _36029_);
  and (_00236_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00237_, _00236_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00238_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _35458_);
  and (_00239_, _00238_, _36029_);
  and (_31342_, _00239_, _00237_);
  and (_00240_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00241_, _00240_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00242_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _35458_);
  and (_00243_, _00242_, _36029_);
  and (_31343_, _00243_, _00241_);
  and (_00244_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00245_, _00244_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00246_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _35458_);
  and (_00247_, _00246_, _36029_);
  and (_31344_, _00247_, _00245_);
  and (_00248_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00249_, _00248_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00251_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _35458_);
  and (_00252_, _00251_, _36029_);
  and (_31345_, _00252_, _00249_);
  and (_00254_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00255_, _00254_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00257_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _35458_);
  and (_00258_, _00257_, _36029_);
  and (_31346_, _00258_, _00255_);
  and (_00260_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00261_, _00260_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00262_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _35458_);
  and (_00264_, _00262_, _36029_);
  and (_31347_, _00264_, _00261_);
  and (_00265_, _35465_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00267_, _00265_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00268_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _35458_);
  and (_00269_, _00268_, _36029_);
  and (_31348_, _00269_, _00267_);
  nand (_00271_, _35472_, _28302_);
  or (_00272_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00274_, _00272_, _36029_);
  and (_31349_, _00274_, _00271_);
  nand (_00275_, _35472_, _28939_);
  or (_00277_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00278_, _00277_, _36029_);
  and (_31351_, _00278_, _00275_);
  nand (_00279_, _35472_, _29584_);
  or (_00280_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00281_, _00280_, _36029_);
  and (_31352_, _00281_, _00279_);
  nand (_00282_, _35472_, _29760_);
  or (_00283_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00284_, _00283_, _36029_);
  and (_31353_, _00284_, _00282_);
  nand (_00285_, _35472_, _29830_);
  or (_00286_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00287_, _00286_, _36029_);
  and (_31354_, _00287_, _00285_);
  nand (_00288_, _35472_, _29903_);
  or (_00289_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00290_, _00289_, _36029_);
  and (_31355_, _00290_, _00288_);
  nand (_00291_, _35472_, _29976_);
  or (_00292_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00294_, _00292_, _36029_);
  and (_31356_, _00294_, _00291_);
  nand (_00296_, _35472_, _27126_);
  or (_00297_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00298_, _00297_, _36029_);
  and (_31357_, _00298_, _00296_);
  nand (_00300_, _35472_, _30667_);
  or (_00301_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00303_, _00301_, _36029_);
  and (_31358_, _00303_, _00300_);
  nand (_00304_, _35472_, _30698_);
  or (_00306_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00307_, _00306_, _36029_);
  and (_31359_, _00307_, _00304_);
  nand (_00309_, _35472_, _30728_);
  or (_00310_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00311_, _00310_, _36029_);
  and (_31360_, _00311_, _00309_);
  nand (_00313_, _35472_, _30757_);
  or (_00314_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00316_, _00314_, _36029_);
  and (_31362_, _00316_, _00313_);
  nand (_00317_, _35472_, _30815_);
  or (_00319_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00320_, _00319_, _36029_);
  and (_31363_, _00320_, _00317_);
  nand (_00321_, _35472_, _30850_);
  or (_00322_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00323_, _00322_, _36029_);
  and (_31364_, _00323_, _00321_);
  nand (_00324_, _35472_, _30914_);
  or (_00325_, _35472_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00326_, _00325_, _36029_);
  and (_31365_, _00326_, _00324_);
  nor (_31573_, _31848_, rst);
  nor (_00327_, _32096_, _32013_);
  and (_00328_, _00327_, _32230_);
  nor (_00329_, _32142_, _31953_);
  and (_00330_, _00329_, _00328_);
  and (_00331_, _00330_, _31091_);
  nand (_00332_, _00327_, _32142_);
  nor (_00333_, _32096_, _32230_);
  and (_00334_, _00333_, _31953_);
  nor (_00335_, _32142_, _32013_);
  and (_00337_, _00335_, _00334_);
  and (_00338_, _00329_, _00327_);
  nor (_00340_, _00338_, _00337_);
  and (_00341_, _00340_, _00332_);
  nand (_00342_, _34738_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  nor (_00344_, _00342_, _00341_);
  not (_00345_, _32058_);
  nor (_00346_, _00345_, _32190_);
  and (_00348_, _00346_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00349_, _00345_, _32190_);
  and (_00350_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00352_, _00350_, _00348_);
  and (_00353_, _32058_, _32190_);
  and (_00354_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_00356_, _32058_, _32190_);
  and (_00357_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00358_, _00357_, _00354_);
  or (_00360_, _00358_, _00352_);
  and (_00361_, _00360_, _31915_);
  not (_00362_, _31915_);
  and (_00364_, _00346_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00365_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00366_, _00365_, _00364_);
  and (_00368_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00369_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_00370_, _00369_, _00368_);
  or (_00371_, _00370_, _00366_);
  and (_00372_, _00371_, _00362_);
  or (_00373_, _00372_, _00361_);
  and (_00374_, _00330_, _00373_);
  nor (_00375_, _31136_, _31125_);
  and (_00376_, _31136_, _31125_);
  nor (_00377_, _00376_, _00375_);
  nor (_00378_, _31285_, _31151_);
  and (_00379_, _31285_, _31151_);
  nor (_00380_, _00379_, _00378_);
  nor (_00381_, _00380_, _00377_);
  and (_00382_, _00380_, _00377_);
  nor (_00383_, _00382_, _00381_);
  nor (_00384_, _31381_, _31370_);
  and (_00385_, _31381_, _31370_);
  nor (_00386_, _00385_, _00384_);
  not (_00387_, _31114_);
  nor (_00388_, _31392_, _00387_);
  and (_00390_, _31392_, _00387_);
  nor (_00391_, _00390_, _00388_);
  nor (_00393_, _00391_, _00386_);
  and (_00394_, _00391_, _00386_);
  or (_00395_, _00394_, _00393_);
  or (_00397_, _00395_, _00383_);
  nand (_00398_, _00395_, _00383_);
  and (_00399_, _00398_, _00397_);
  or (_00401_, _00399_, _00362_);
  or (_00402_, _31915_, _31058_);
  and (_00403_, _00402_, _00353_);
  and (_00405_, _00403_, _00401_);
  or (_00406_, _00362_, _31003_);
  or (_00407_, _31915_, _31068_);
  and (_00409_, _00407_, _00349_);
  and (_00410_, _00409_, _00406_);
  and (_00411_, _00356_, _00362_);
  and (_00413_, _00411_, _30994_);
  and (_00414_, _00356_, _31915_);
  and (_00415_, _00414_, _31047_);
  or (_00417_, _00415_, _00413_);
  or (_00418_, _00417_, _00410_);
  or (_00419_, _00362_, _31039_);
  or (_00421_, _31915_, _31085_);
  and (_00422_, _00421_, _00346_);
  and (_00423_, _00422_, _00419_);
  or (_00424_, _00423_, _00418_);
  or (_00425_, _00424_, _00405_);
  and (_00426_, _00425_, _00337_);
  and (_00427_, _30221_, _30351_);
  nor (_00428_, _00427_, _30335_);
  nor (_00429_, _30348_, _30332_);
  and (_00430_, _00429_, _00428_);
  nor (_00431_, _34242_, _34173_);
  and (_00432_, _00431_, _00430_);
  nor (_00433_, _34244_, _34176_);
  and (_00434_, _30220_, _30218_);
  nor (_00435_, _00434_, _34345_);
  and (_00436_, _00435_, _00433_);
  and (_00437_, _00436_, _34519_);
  and (_00438_, _00437_, _00432_);
  and (_00439_, _00438_, _30309_);
  nor (_00440_, _00439_, _29998_);
  and (_00441_, _34702_, p1in_reg[5]);
  and (_00443_, _34698_, p1_in[5]);
  or (_00444_, _00443_, _00441_);
  or (_00446_, _00444_, _00440_);
  not (_00447_, _00440_);
  or (_00448_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00450_, _00448_, _00446_);
  and (_00451_, _00450_, _00349_);
  or (_00452_, _00451_, _31915_);
  and (_00454_, _34702_, p1in_reg[7]);
  and (_00455_, _34698_, p1_in[7]);
  or (_00456_, _00455_, _00454_);
  or (_00458_, _00456_, _00440_);
  nand (_00459_, _00440_, _31417_);
  and (_00460_, _00459_, _00458_);
  and (_00462_, _00460_, _00356_);
  and (_00463_, _34702_, p1in_reg[6]);
  and (_00464_, _34698_, p1_in[6]);
  or (_00466_, _00464_, _00463_);
  or (_00467_, _00466_, _00440_);
  nand (_00468_, _00440_, _31635_);
  and (_00470_, _00468_, _00467_);
  and (_00471_, _00470_, _00346_);
  and (_00472_, _34702_, p1in_reg[4]);
  and (_00474_, _34698_, p1_in[4]);
  or (_00475_, _00474_, _00472_);
  or (_00476_, _00475_, _00440_);
  or (_00477_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00478_, _00477_, _00476_);
  and (_00479_, _00478_, _00353_);
  or (_00480_, _00479_, _00471_);
  or (_00481_, _00480_, _00462_);
  or (_00482_, _00481_, _00452_);
  and (_00483_, _32142_, _32014_);
  and (_00484_, _00483_, _00334_);
  and (_00485_, _34702_, p1in_reg[1]);
  and (_00486_, _34698_, p1_in[1]);
  or (_00487_, _00486_, _00485_);
  or (_00488_, _00487_, _00440_);
  nand (_00489_, _00440_, _31568_);
  and (_00490_, _00489_, _00488_);
  and (_00491_, _00490_, _00349_);
  or (_00492_, _00491_, _00362_);
  and (_00493_, _34702_, p1in_reg[3]);
  and (_00494_, _34698_, p1_in[3]);
  or (_00496_, _00494_, _00493_);
  or (_00497_, _00496_, _00440_);
  or (_00499_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00500_, _00499_, _00497_);
  and (_00501_, _00500_, _00356_);
  and (_00503_, _34702_, p1in_reg[2]);
  and (_00504_, _34698_, p1_in[2]);
  or (_00505_, _00504_, _00503_);
  or (_00507_, _00505_, _00440_);
  nand (_00508_, _00440_, _31582_);
  and (_00509_, _00508_, _00507_);
  and (_00511_, _00509_, _00346_);
  and (_00512_, _34702_, p1in_reg[0]);
  and (_00513_, _34698_, p1_in[0]);
  or (_00515_, _00513_, _00512_);
  or (_00516_, _00515_, _00440_);
  nand (_00517_, _00440_, _31555_);
  and (_00519_, _00517_, _00516_);
  and (_00520_, _00519_, _00353_);
  or (_00521_, _00520_, _00511_);
  or (_00523_, _00521_, _00501_);
  or (_00524_, _00523_, _00492_);
  and (_00525_, _00524_, _00484_);
  and (_00527_, _00525_, _00482_);
  and (_00528_, _34702_, p2in_reg[2]);
  and (_00529_, _34698_, p2_in[2]);
  or (_00530_, _00529_, _00528_);
  or (_00531_, _00530_, _00440_);
  nand (_00532_, _00440_, _31681_);
  and (_00533_, _00532_, _00531_);
  and (_00534_, _00533_, _00346_);
  and (_00535_, _34702_, p2in_reg[0]);
  and (_00536_, _34698_, p2_in[0]);
  or (_00537_, _00536_, _00535_);
  or (_00538_, _00537_, _00440_);
  nand (_00539_, _00440_, _31648_);
  and (_00540_, _00539_, _00538_);
  and (_00541_, _00540_, _00353_);
  or (_00542_, _00541_, _00534_);
  and (_00543_, _34702_, p2in_reg[1]);
  and (_00544_, _34698_, p2_in[1]);
  or (_00545_, _00544_, _00543_);
  or (_00546_, _00545_, _00440_);
  nand (_00547_, _00440_, _31661_);
  and (_00549_, _00547_, _00546_);
  and (_00550_, _00549_, _00349_);
  and (_00552_, _34702_, p2in_reg[3]);
  and (_00553_, _34698_, p2_in[3]);
  or (_00554_, _00553_, _00552_);
  or (_00556_, _00554_, _00440_);
  or (_00557_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00558_, _00557_, _00556_);
  and (_00560_, _00558_, _00356_);
  or (_00561_, _00560_, _00550_);
  or (_00562_, _00561_, _00542_);
  and (_00564_, _00562_, _31915_);
  and (_00565_, _34702_, p2in_reg[6]);
  and (_00566_, _34698_, p2_in[6]);
  or (_00568_, _00566_, _00565_);
  or (_00569_, _00568_, _00440_);
  nand (_00570_, _00440_, _31743_);
  and (_00572_, _00570_, _00569_);
  and (_00573_, _00572_, _00346_);
  and (_00574_, _34702_, p2in_reg[4]);
  and (_00576_, _34698_, p2_in[4]);
  or (_00577_, _00576_, _00574_);
  or (_00578_, _00577_, _00440_);
  or (_00580_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00581_, _00580_, _00578_);
  and (_00582_, _00581_, _00353_);
  or (_00583_, _00582_, _00573_);
  and (_00584_, _34702_, p2in_reg[5]);
  and (_00585_, _34698_, p2_in[5]);
  or (_00586_, _00585_, _00584_);
  or (_00587_, _00586_, _00440_);
  or (_00588_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00589_, _00588_, _00587_);
  and (_00590_, _00589_, _00349_);
  and (_00591_, _34702_, p2in_reg[7]);
  and (_00592_, _34698_, p2_in[7]);
  or (_00593_, _00592_, _00591_);
  or (_00594_, _00593_, _00440_);
  nand (_00595_, _00440_, _31435_);
  and (_00596_, _00595_, _00594_);
  and (_00597_, _00596_, _00356_);
  or (_00598_, _00597_, _00590_);
  or (_00599_, _00598_, _00583_);
  and (_00600_, _00599_, _00362_);
  or (_00602_, _00600_, _00564_);
  and (_00603_, _32142_, _31954_);
  and (_00605_, _00603_, _00328_);
  and (_00606_, _00605_, _00602_);
  or (_00607_, _00606_, _00527_);
  and (_00609_, _00603_, _00327_);
  and (_00610_, _34702_, p3in_reg[0]);
  and (_00611_, _34698_, p3_in[0]);
  or (_00613_, _00611_, _00610_);
  or (_00614_, _00613_, _00440_);
  nand (_00615_, _00440_, _31756_);
  and (_00617_, _00615_, _00614_);
  and (_00618_, _00617_, _00353_);
  and (_00619_, _34702_, p3in_reg[2]);
  and (_00621_, _34698_, p3_in[2]);
  or (_00622_, _00621_, _00619_);
  or (_00623_, _00622_, _00440_);
  nand (_00625_, _00440_, _31782_);
  and (_00626_, _00625_, _00623_);
  and (_00627_, _00626_, _00346_);
  or (_00629_, _00627_, _00618_);
  and (_00630_, _34702_, p3in_reg[1]);
  and (_00631_, _34698_, p3_in[1]);
  or (_00633_, _00631_, _00630_);
  or (_00634_, _00633_, _00440_);
  nand (_00635_, _00440_, _31769_);
  and (_00636_, _00635_, _00634_);
  and (_00637_, _00636_, _00349_);
  and (_00638_, _34702_, p3in_reg[3]);
  and (_00639_, _34698_, p3_in[3]);
  or (_00640_, _00639_, _00638_);
  or (_00641_, _00640_, _00440_);
  or (_00642_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00643_, _00642_, _00641_);
  and (_00644_, _00643_, _00356_);
  or (_00645_, _00644_, _00637_);
  or (_00646_, _00645_, _00629_);
  and (_00647_, _00646_, _31915_);
  and (_00648_, _34702_, p3in_reg[4]);
  and (_00649_, _34698_, p3_in[4]);
  or (_00650_, _00649_, _00648_);
  or (_00651_, _00650_, _00440_);
  or (_00652_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00653_, _00652_, _00651_);
  and (_00654_, _00653_, _00353_);
  and (_00655_, _34702_, p3in_reg[6]);
  and (_00656_, _34698_, p3_in[6]);
  or (_00657_, _00656_, _00655_);
  or (_00658_, _00657_, _00440_);
  nand (_00659_, _00440_, _31831_);
  and (_00660_, _00659_, _00658_);
  and (_00661_, _00660_, _00346_);
  or (_00662_, _00661_, _00654_);
  and (_00663_, _34702_, p3in_reg[5]);
  and (_00664_, _34698_, p3_in[5]);
  or (_00665_, _00664_, _00663_);
  or (_00666_, _00665_, _00440_);
  or (_00667_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00668_, _00667_, _00666_);
  and (_00669_, _00668_, _00349_);
  and (_00670_, _34702_, p3in_reg[7]);
  and (_00671_, _34698_, p3_in[7]);
  or (_00672_, _00671_, _00670_);
  or (_00673_, _00672_, _00440_);
  nand (_00674_, _00440_, _31451_);
  and (_00675_, _00674_, _00673_);
  and (_00676_, _00675_, _00356_);
  or (_00677_, _00676_, _00669_);
  or (_00678_, _00677_, _00662_);
  and (_00679_, _00678_, _00362_);
  or (_00680_, _00679_, _00647_);
  and (_00681_, _00680_, _00609_);
  and (_00682_, _00346_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00683_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00684_, _00683_, _00682_);
  and (_00685_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00686_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00687_, _00686_, _00685_);
  or (_00688_, _00687_, _00684_);
  and (_00689_, _00688_, _31915_);
  and (_00690_, _00346_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_00691_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_00692_, _00691_, _00690_);
  and (_00693_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00694_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00695_, _00694_, _00693_);
  or (_00696_, _00695_, _00692_);
  and (_00697_, _00696_, _00362_);
  or (_00698_, _00697_, _00689_);
  and (_00699_, _00698_, _00338_);
  or (_00700_, _00699_, _00681_);
  and (_00701_, _00700_, _32231_);
  and (_00702_, _34702_, p0in_reg[6]);
  and (_00703_, _34698_, p0_in[6]);
  or (_00704_, _00703_, _00702_);
  or (_00705_, _00704_, _00440_);
  nand (_00706_, _00440_, _31537_);
  and (_00707_, _00706_, _00705_);
  and (_00708_, _00707_, _00346_);
  or (_00709_, _00708_, _31915_);
  and (_00710_, _34702_, p0in_reg[7]);
  and (_00711_, _34698_, p0_in[7]);
  or (_00712_, _00711_, _00710_);
  or (_00713_, _00712_, _00440_);
  nand (_00714_, _00440_, _31403_);
  and (_00715_, _00714_, _00713_);
  and (_00716_, _00715_, _00356_);
  and (_00717_, _34702_, p0in_reg[5]);
  and (_00718_, _34698_, p0_in[5]);
  or (_00719_, _00718_, _00717_);
  or (_00720_, _00719_, _00440_);
  or (_00721_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_00722_, _00721_, _00720_);
  and (_00723_, _00722_, _00349_);
  and (_00724_, _34702_, p0in_reg[4]);
  and (_00725_, _34698_, p0_in[4]);
  or (_00726_, _00725_, _00724_);
  or (_00727_, _00726_, _00440_);
  or (_00728_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00729_, _00728_, _00727_);
  and (_00730_, _00729_, _00353_);
  or (_00731_, _00730_, _00723_);
  or (_00732_, _00731_, _00716_);
  or (_00733_, _00732_, _00709_);
  and (_00734_, _32230_, _31953_);
  and (_00735_, _00734_, _00483_);
  and (_00736_, _00735_, _32095_);
  and (_00737_, _34702_, p0in_reg[2]);
  and (_00738_, _34698_, p0_in[2]);
  or (_00739_, _00738_, _00737_);
  or (_00740_, _00739_, _00440_);
  nand (_00741_, _00440_, _31481_);
  and (_00742_, _00741_, _00740_);
  and (_00743_, _00742_, _00346_);
  or (_00744_, _00743_, _00362_);
  and (_00745_, _34702_, p0in_reg[3]);
  and (_00746_, _34698_, p0_in[3]);
  or (_00747_, _00746_, _00745_);
  or (_00748_, _00747_, _00440_);
  or (_00749_, _00447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00750_, _00749_, _00748_);
  and (_00751_, _00750_, _00356_);
  and (_00752_, _34702_, p0in_reg[1]);
  and (_00753_, _34698_, p0_in[1]);
  or (_00754_, _00753_, _00752_);
  or (_00755_, _00754_, _00440_);
  nand (_00756_, _00440_, _31477_);
  and (_00757_, _00756_, _00755_);
  and (_00758_, _00757_, _00349_);
  and (_00759_, _34702_, p0in_reg[0]);
  and (_00760_, _34698_, p0_in[0]);
  or (_00761_, _00760_, _00759_);
  or (_00762_, _00761_, _00440_);
  nand (_00763_, _00440_, _31458_);
  and (_00764_, _00763_, _00762_);
  and (_00765_, _00764_, _00353_);
  or (_00766_, _00765_, _00758_);
  or (_00767_, _00766_, _00751_);
  or (_00768_, _00767_, _00744_);
  and (_00769_, _00768_, _00736_);
  and (_00770_, _00769_, _00733_);
  or (_00771_, _00770_, _00701_);
  or (_00772_, _00771_, _00607_);
  or (_00773_, _00772_, _00426_);
  nor (_00774_, _00773_, _00374_);
  or (_00775_, _00774_, _00344_);
  nand (_00776_, _00344_, _28359_);
  and (_00777_, _00776_, _00775_);
  nor (_00778_, _00777_, _00331_);
  or (_00779_, _31915_, _31381_);
  or (_00780_, _00362_, _31136_);
  and (_00781_, _00780_, _00349_);
  and (_00782_, _00781_, _00779_);
  or (_00783_, _31915_, _31392_);
  nand (_00784_, _31915_, _31151_);
  and (_00785_, _00784_, _00346_);
  and (_00786_, _00785_, _00783_);
  or (_00787_, _00362_, _31125_);
  or (_00788_, _31915_, _31370_);
  and (_00789_, _00788_, _00353_);
  and (_00790_, _00789_, _00787_);
  or (_00791_, _00790_, _00786_);
  and (_00792_, _00411_, _31114_);
  not (_00793_, _00414_);
  nor (_00794_, _00793_, _31285_);
  or (_00795_, _00794_, _00792_);
  or (_00796_, _00795_, _00791_);
  or (_00797_, _00796_, _00782_);
  and (_00798_, _00797_, _00331_);
  or (_00799_, _00798_, _00778_);
  nor (_00800_, _00332_, _00440_);
  nand (_00801_, _34743_, _30989_);
  or (_00802_, _00801_, _00800_);
  or (_00803_, _00802_, _00341_);
  and (_00804_, _00803_, _00799_);
  or (_00805_, _31915_, _32111_);
  nand (_00806_, _31915_, _30455_);
  and (_00807_, _00806_, _00346_);
  and (_00808_, _00807_, _00805_);
  or (_00809_, _31915_, _32219_);
  nand (_00810_, _31915_, _30470_);
  and (_00811_, _00810_, _00353_);
  and (_00812_, _00811_, _00809_);
  or (_00813_, _00812_, _00808_);
  nand (_00814_, _31915_, _30462_);
  or (_00815_, _31915_, _31944_);
  and (_00816_, _00815_, _00349_);
  and (_00817_, _00816_, _00814_);
  and (_00818_, _00411_, _30413_);
  and (_00819_, _00414_, _32089_);
  or (_00820_, _00819_, _00818_);
  or (_00821_, _00820_, _00817_);
  nor (_00822_, _00821_, _00813_);
  nor (_00823_, _00803_, _00822_);
  or (_00824_, _00823_, _00804_);
  and (_31601_, _00824_, _36029_);
  and (_00825_, _00736_, _00414_);
  nand (_00826_, _00825_, _30537_);
  nor (_00827_, _32230_, _31954_);
  and (_00828_, _32095_, _31915_);
  and (_00829_, _00828_, _00353_);
  and (_00830_, _00829_, _00827_);
  and (_00831_, _00830_, _00335_);
  nand (_00832_, _00831_, _30980_);
  and (_00833_, _00832_, _00826_);
  nor (_00834_, _00833_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_00835_, _00834_);
  not (_00836_, _30985_);
  nor (_00837_, _00411_, _00836_);
  and (_00838_, _00837_, _34743_);
  or (_00839_, _31091_, _31087_);
  and (_00840_, _00829_, _32230_);
  and (_00841_, _00840_, _31954_);
  and (_00842_, _00841_, _00335_);
  and (_00843_, _00842_, _00839_);
  nor (_00844_, _00843_, _00838_);
  and (_00845_, _00844_, _34741_);
  and (_00846_, _00845_, _00835_);
  and (_00847_, _00828_, _00346_);
  and (_00848_, _00847_, _00735_);
  and (_00849_, _00848_, _30537_);
  or (_00850_, _00849_, rst);
  nor (_31603_, _00850_, _00846_);
  not (_00851_, _00849_);
  and (_00852_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00853_, _00829_, _32231_);
  and (_00854_, _00853_, _31954_);
  and (_00855_, _00854_, _00335_);
  and (_00856_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_00857_, _00828_, _00356_);
  and (_00858_, _00857_, _00735_);
  and (_00859_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_00860_, _00859_, _00856_);
  and (_00861_, _00828_, _00349_);
  and (_00862_, _00861_, _00735_);
  and (_00863_, _00862_, _31977_);
  nor (_00864_, _32230_, _31953_);
  and (_00865_, _00864_, _00483_);
  and (_00866_, _00865_, _00829_);
  and (_00867_, _00866_, _00675_);
  or (_00868_, _00867_, _00863_);
  or (_00869_, _00868_, _00860_);
  or (_00870_, _00869_, _00852_);
  and (_00871_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00872_, _00841_, _00483_);
  and (_00873_, _00872_, _00596_);
  and (_00874_, _00830_, _00483_);
  and (_00875_, _00874_, _00460_);
  or (_00876_, _00875_, _00873_);
  and (_00877_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_00878_, _00829_, _00735_);
  and (_00879_, _00878_, _00715_);
  or (_00880_, _00879_, _00877_);
  or (_00881_, _00880_, _00876_);
  or (_00882_, _00881_, _00871_);
  or (_00883_, _00882_, _00870_);
  and (_00884_, _00883_, _00846_);
  nor (_00885_, _00846_, _16547_);
  or (_00886_, _00885_, _00884_);
  and (_00887_, _00886_, _00851_);
  nor (_00888_, _00851_, _27126_);
  or (_00889_, _00888_, _00887_);
  and (_31604_, _00889_, _36029_);
  and (_00890_, _00831_, _00399_);
  and (_00891_, _00874_, _00519_);
  and (_00892_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_00893_, _00892_, _00891_);
  or (_00894_, _00893_, _00890_);
  nand (_00895_, _00842_, _31091_);
  nand (_00896_, _00858_, _30537_);
  nand (_00897_, _00842_, _31087_);
  and (_00898_, _00897_, _00832_);
  and (_00899_, _00898_, _00896_);
  or (_00900_, _00899_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00901_, _34738_, _27781_);
  and (_00902_, _00901_, _27158_);
  not (_00903_, _00411_);
  nand (_00904_, _00903_, _34743_);
  nor (_00905_, _00904_, _00836_);
  nor (_00906_, _00905_, _00902_);
  and (_00907_, _00906_, _00900_);
  and (_00908_, _00907_, _00895_);
  and (_00909_, _00854_, _00483_);
  and (_00910_, _00909_, _00617_);
  and (_00911_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_00912_, _00911_, _00910_);
  and (_00913_, _00862_, _32054_);
  and (_00914_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00915_, _00878_, _00764_);
  or (_00916_, _00915_, _00914_);
  nor (_00917_, _00916_, _00913_);
  and (_00918_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00919_, _00872_, _00540_);
  nor (_00920_, _00919_, _00918_);
  and (_00921_, _00920_, _00917_);
  and (_00922_, _00921_, _00912_);
  nand (_00923_, _00922_, _00908_);
  or (_00924_, _00923_, _00894_);
  or (_00925_, _00908_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_00926_, _00925_, _00924_);
  or (_00927_, _00926_, _00849_);
  nand (_00928_, _00849_, _28302_);
  and (_00929_, _00928_, _36029_);
  and (_31664_, _00929_, _00927_);
  and (_00930_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00931_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00932_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00933_, _00932_, _00931_);
  and (_00934_, _00862_, _32183_);
  and (_00935_, _00866_, _00636_);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00933_);
  or (_00938_, _00937_, _00930_);
  and (_00939_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00940_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_00941_, _00878_, _00757_);
  or (_00942_, _00941_, _00940_);
  and (_00943_, _00874_, _00490_);
  and (_00944_, _32230_, _31954_);
  and (_00945_, _00944_, _00483_);
  and (_00946_, _00945_, _00829_);
  and (_00947_, _00946_, _00549_);
  or (_00948_, _00947_, _00943_);
  or (_00949_, _00948_, _00942_);
  or (_00950_, _00949_, _00939_);
  or (_00951_, _00950_, _00938_);
  and (_00952_, _00951_, _00846_);
  nor (_00953_, _00846_, _16372_);
  or (_00954_, _00953_, _00952_);
  and (_00955_, _00954_, _00851_);
  nor (_00956_, _00851_, _28939_);
  or (_00957_, _00956_, _00955_);
  and (_31666_, _00957_, _36029_);
  and (_00958_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00959_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00960_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00961_, _00960_, _00959_);
  and (_00962_, _00862_, _31877_);
  and (_00963_, _00866_, _00626_);
  or (_00964_, _00963_, _00962_);
  or (_00965_, _00964_, _00961_);
  or (_00966_, _00965_, _00958_);
  and (_00967_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00968_, _00874_, _00509_);
  and (_00969_, _00946_, _00533_);
  or (_00970_, _00969_, _00968_);
  and (_00971_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_00972_, _00878_, _00742_);
  or (_00973_, _00972_, _00971_);
  or (_00974_, _00973_, _00970_);
  or (_00975_, _00974_, _00967_);
  or (_00976_, _00975_, _00966_);
  and (_00977_, _00976_, _00846_);
  nor (_00978_, _00846_, _15031_);
  or (_00979_, _00978_, _00977_);
  and (_00980_, _00979_, _00851_);
  nor (_00981_, _00851_, _29584_);
  or (_00982_, _00981_, _00980_);
  and (_31667_, _00982_, _36029_);
  and (_00983_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00984_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00985_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00986_, _00985_, _00984_);
  and (_00987_, _00862_, _32079_);
  and (_00988_, _00866_, _00643_);
  or (_00989_, _00988_, _00987_);
  or (_00990_, _00989_, _00986_);
  or (_00991_, _00990_, _00983_);
  and (_00992_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00993_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_00994_, _00878_, _00750_);
  or (_00995_, _00994_, _00993_);
  and (_00996_, _00872_, _00558_);
  and (_00997_, _00874_, _00500_);
  or (_00998_, _00997_, _00996_);
  or (_00999_, _00998_, _00995_);
  or (_01000_, _00999_, _00992_);
  or (_01001_, _01000_, _00991_);
  and (_01002_, _01001_, _00846_);
  nor (_01003_, _00846_, _16057_);
  or (_01004_, _01003_, _01002_);
  and (_01005_, _01004_, _00851_);
  nor (_01006_, _00851_, _29760_);
  or (_01007_, _01006_, _01005_);
  and (_31668_, _01007_, _36029_);
  and (_01008_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01009_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01010_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01011_, _01010_, _01009_);
  and (_01012_, _00862_, _32226_);
  and (_01013_, _00866_, _00653_);
  or (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _01011_);
  or (_01016_, _01015_, _01008_);
  and (_01017_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01018_, _00872_, _00581_);
  and (_01019_, _00874_, _00478_);
  or (_01020_, _01019_, _01018_);
  and (_01021_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01022_, _00878_, _00729_);
  or (_01023_, _01022_, _01021_);
  or (_01024_, _01023_, _01020_);
  or (_01025_, _01024_, _01017_);
  or (_01026_, _01025_, _01016_);
  and (_01027_, _01026_, _00846_);
  nor (_01028_, _00846_, _15228_);
  or (_01029_, _01028_, _01027_);
  and (_01030_, _01029_, _00851_);
  nor (_01031_, _00851_, _29830_);
  or (_01032_, _01031_, _01030_);
  and (_31669_, _01032_, _36029_);
  and (_01033_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01034_, _00862_, _31917_);
  and (_01035_, _00909_, _00668_);
  or (_01036_, _01035_, _01034_);
  and (_01037_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01038_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01039_, _01038_, _01037_);
  or (_01040_, _01039_, _01036_);
  or (_01041_, _01040_, _01033_);
  and (_01042_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01043_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01044_, _00878_, _00722_);
  or (_01045_, _01044_, _01043_);
  and (_01046_, _00872_, _00589_);
  and (_01047_, _00874_, _00450_);
  or (_01048_, _01047_, _01046_);
  or (_01049_, _01048_, _01045_);
  or (_01050_, _01049_, _01042_);
  or (_01051_, _01050_, _01041_);
  and (_01052_, _01051_, _00846_);
  nor (_01054_, _00846_, _16209_);
  or (_01055_, _01054_, _01052_);
  and (_01056_, _01055_, _00851_);
  nor (_01057_, _00851_, _29903_);
  or (_01058_, _01057_, _01056_);
  and (_31670_, _01058_, _36029_);
  and (_01059_, _00848_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01060_, _00855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01061_, _00858_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01062_, _01061_, _01060_);
  and (_01063_, _00862_, _32109_);
  and (_01064_, _00866_, _00660_);
  or (_01065_, _01064_, _01063_);
  or (_01066_, _01065_, _01062_);
  or (_01067_, _01066_, _01059_);
  and (_01068_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01069_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01070_, _00878_, _00707_);
  or (_01071_, _01070_, _01069_);
  and (_01072_, _00874_, _00470_);
  and (_01073_, _00946_, _00572_);
  or (_01074_, _01073_, _01072_);
  or (_01075_, _01074_, _01071_);
  or (_01076_, _01075_, _01068_);
  or (_01077_, _01076_, _01067_);
  and (_01078_, _01077_, _00846_);
  nor (_01079_, _00846_, _15567_);
  or (_01080_, _01079_, _01078_);
  and (_01081_, _01080_, _00851_);
  nor (_01082_, _00851_, _29976_);
  or (_01084_, _01082_, _01081_);
  and (_31671_, _01084_, _36029_);
  and (_31715_, _32246_, _36029_);
  and (_31716_, _32319_, _36029_);
  nor (_31718_, _31915_, rst);
  and (_31733_, _32337_, _36029_);
  and (_31734_, _32350_, _36029_);
  and (_31736_, _32363_, _36029_);
  and (_31737_, _32372_, _36029_);
  and (_31738_, _32382_, _36029_);
  and (_31739_, _32391_, _36029_);
  and (_31740_, _32402_, _36029_);
  nor (_31741_, _32058_, rst);
  nor (_31742_, _32190_, rst);
  not (_01085_, _33269_);
  nor (_01086_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01087_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01088_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01087_);
  nor (_01089_, _01088_, _01086_);
  nor (_01091_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01092_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01087_);
  nor (_01093_, _01092_, _01091_);
  not (_01094_, _01093_);
  nor (_01095_, _01094_, _01089_);
  nor (_01096_, _01093_, _01089_);
  not (_01097_, _01096_);
  nor (_01098_, _35706_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01099_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01087_);
  nor (_01100_, _01099_, _01098_);
  and (_01101_, _01100_, _01097_);
  nor (_01102_, _01100_, _01097_);
  nor (_01103_, _01102_, _01101_);
  not (_01104_, _01103_);
  nor (_01105_, _35724_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01106_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01087_);
  nor (_01107_, _01106_, _01105_);
  not (_01108_, _01107_);
  and (_01109_, _01108_, _01101_);
  nor (_01110_, _01108_, _01101_);
  nor (_01111_, _01110_, _01109_);
  and (_01112_, _01111_, _01104_);
  and (_01113_, _01112_, _01095_);
  and (_01114_, _01113_, _01085_);
  not (_01115_, _33627_);
  nor (_01116_, _01111_, _01103_);
  and (_01117_, _01116_, _01095_);
  and (_01118_, _01117_, _01115_);
  not (_01119_, _33586_);
  and (_01120_, _01094_, _01089_);
  and (_01121_, _01120_, _01116_);
  and (_01122_, _01121_, _01119_);
  or (_01123_, _01122_, _01118_);
  or (_01124_, _01123_, _01114_);
  not (_01125_, _33463_);
  and (_01126_, _01108_, _01103_);
  and (_01127_, _01126_, _01095_);
  and (_01128_, _01127_, _01125_);
  not (_01129_, _33504_);
  and (_01130_, _01093_, _01089_);
  and (_01131_, _01126_, _01130_);
  and (_01132_, _01131_, _01129_);
  or (_01133_, _01132_, _01128_);
  not (_01134_, _33420_);
  and (_01135_, _01126_, _01120_);
  and (_01136_, _01135_, _01134_);
  not (_01137_, _33713_);
  and (_01138_, _01107_, _01102_);
  and (_01139_, _01138_, _01137_);
  not (_01140_, _33545_);
  and (_01141_, _01100_, _01096_);
  and (_01142_, _01108_, _01141_);
  and (_01143_, _01142_, _01140_);
  or (_01144_, _01143_, _01139_);
  and (_01145_, _01107_, _01141_);
  and (_01146_, _01145_, _33937_);
  not (_01147_, _33379_);
  and (_01148_, _01108_, _01102_);
  and (_01149_, _01148_, _01147_);
  or (_01150_, _01149_, _01146_);
  or (_01151_, _01150_, _01144_);
  or (_01152_, _01151_, _01136_);
  or (_01153_, _01152_, _01133_);
  not (_01154_, _33228_);
  and (_01155_, _01120_, _01112_);
  and (_01156_, _01155_, _01154_);
  not (_01157_, _33310_);
  and (_01158_, _01112_, _01130_);
  and (_01159_, _01158_, _01157_);
  or (_01160_, _01159_, _01156_);
  not (_01161_, _33668_);
  and (_01162_, _01116_, _01130_);
  and (_01163_, _01162_, _01161_);
  not (_01164_, _33881_);
  and (_01165_, _01110_, _01130_);
  and (_01166_, _01165_, _01164_);
  not (_01167_, _33823_);
  and (_01168_, _01110_, _01095_);
  and (_01169_, _01168_, _01167_);
  not (_01170_, _33767_);
  and (_01171_, _01120_, _01110_);
  and (_01172_, _01171_, _01170_);
  or (_01173_, _01172_, _01169_);
  or (_01174_, _01173_, _01166_);
  or (_01175_, _01174_, _01163_);
  or (_01176_, _01175_, _01160_);
  or (_01177_, _01176_, _01153_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01177_, _01124_);
  and (_01178_, _01155_, _01164_);
  and (_01179_, _01165_, _01170_);
  and (_01180_, _01168_, _01137_);
  or (_01181_, _01180_, _01179_);
  or (_01182_, _01181_, _01178_);
  and (_01183_, _01113_, _33937_);
  and (_01184_, _01162_, _01119_);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01185_, _01182_);
  and (_01187_, _01131_, _01134_);
  and (_01188_, _01127_, _01147_);
  or (_01189_, _01188_, _01187_);
  and (_01190_, _01142_, _01125_);
  or (_01191_, _01190_, _01189_);
  and (_01192_, _01148_, _01085_);
  and (_01193_, _01121_, _01129_);
  or (_01194_, _01193_, _01192_);
  or (_01195_, _01194_, _01191_);
  or (_01196_, _01195_, _01186_);
  and (_01197_, _01145_, _01167_);
  and (_01198_, _01135_, _01157_);
  and (_01199_, _01158_, _01154_);
  or (_01200_, _01199_, _01198_);
  and (_01201_, _01117_, _01140_);
  and (_01202_, _01138_, _01115_);
  and (_01203_, _01171_, _01161_);
  or (_01204_, _01203_, _01202_);
  or (_01205_, _01204_, _01201_);
  or (_01206_, _01205_, _01200_);
  or (_01207_, _01206_, _01197_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01207_, _01196_);
  and (_01208_, _01162_, _01115_);
  and (_01209_, _01155_, _33937_);
  and (_01210_, _01113_, _01154_);
  or (_01211_, _01210_, _01209_);
  or (_01212_, _01211_, _01208_);
  and (_01213_, _01127_, _01134_);
  and (_01214_, _01142_, _01129_);
  and (_01215_, _01148_, _01157_);
  or (_01216_, _01215_, _01214_);
  and (_01217_, _01145_, _01164_);
  and (_01218_, _01138_, _01161_);
  or (_01219_, _01218_, _01217_);
  or (_01220_, _01219_, _01216_);
  or (_01221_, _01220_, _01213_);
  and (_01222_, _01131_, _01125_);
  and (_01223_, _01135_, _01147_);
  or (_01224_, _01223_, _01222_);
  or (_01225_, _01224_, _01221_);
  and (_01226_, _01117_, _01119_);
  and (_01227_, _01165_, _01167_);
  and (_01228_, _01168_, _01170_);
  and (_01229_, _01171_, _01137_);
  or (_01230_, _01229_, _01228_);
  or (_01231_, _01230_, _01227_);
  or (_01232_, _01231_, _01226_);
  and (_01233_, _01158_, _01085_);
  and (_01234_, _01121_, _01140_);
  or (_01235_, _01234_, _01233_);
  or (_01236_, _01235_, _01232_);
  or (_01237_, _01236_, _01225_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01237_, _01212_);
  and (_01238_, _01113_, _01164_);
  and (_01239_, _01162_, _01140_);
  and (_01240_, _01121_, _01125_);
  or (_01241_, _01240_, _01239_);
  or (_01242_, _01241_, _01238_);
  and (_01243_, _01127_, _01157_);
  and (_01244_, _01145_, _01170_);
  and (_01245_, _01142_, _01134_);
  or (_01246_, _01245_, _01244_);
  and (_01247_, _01138_, _01119_);
  and (_01248_, _01148_, _01154_);
  or (_01249_, _01248_, _01247_);
  or (_01250_, _01249_, _01246_);
  or (_01251_, _01250_, _01243_);
  and (_01252_, _01135_, _01085_);
  and (_01253_, _01131_, _01147_);
  or (_01254_, _01253_, _01252_);
  or (_01255_, _01254_, _01251_);
  and (_01256_, _01117_, _01129_);
  and (_01257_, _01171_, _01115_);
  and (_01258_, _01165_, _01137_);
  and (_01259_, _01168_, _01161_);
  or (_01260_, _01259_, _01258_);
  or (_01261_, _01260_, _01257_);
  or (_01262_, _01261_, _01256_);
  and (_01263_, _01158_, _33937_);
  and (_01264_, _01155_, _01167_);
  or (_01265_, _01264_, _01263_);
  or (_01266_, _01265_, _01262_);
  or (_01267_, _01266_, _01255_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01267_, _01242_);
  not (_01268_, _33274_);
  and (_01269_, _01113_, _01268_);
  not (_01270_, _33673_);
  and (_01271_, _01162_, _01270_);
  not (_01272_, _33632_);
  and (_01273_, _01117_, _01272_);
  or (_01274_, _01273_, _01271_);
  or (_01275_, _01274_, _01269_);
  not (_01276_, _33468_);
  and (_01277_, _01127_, _01276_);
  not (_01278_, _33509_);
  and (_01279_, _01131_, _01278_);
  or (_01280_, _01279_, _01277_);
  not (_01281_, _33425_);
  and (_01282_, _01135_, _01281_);
  not (_01283_, _33720_);
  and (_01284_, _01138_, _01283_);
  not (_01285_, _33550_);
  and (_01286_, _01142_, _01285_);
  or (_01287_, _01286_, _01284_);
  and (_01288_, _01145_, _33944_);
  not (_01289_, _33384_);
  and (_01290_, _01148_, _01289_);
  or (_01291_, _01290_, _01288_);
  or (_01292_, _01291_, _01287_);
  or (_01293_, _01292_, _01282_);
  or (_01294_, _01293_, _01280_);
  not (_01295_, _33233_);
  and (_01296_, _01155_, _01295_);
  not (_01297_, _33316_);
  and (_01298_, _01158_, _01297_);
  or (_01299_, _01298_, _01296_);
  not (_01300_, _33591_);
  and (_01301_, _01121_, _01300_);
  not (_01302_, _33830_);
  and (_01303_, _01168_, _01302_);
  not (_01304_, _33888_);
  and (_01305_, _01165_, _01304_);
  not (_01306_, _33774_);
  and (_01307_, _01171_, _01306_);
  or (_01308_, _01307_, _01305_);
  or (_01309_, _01308_, _01303_);
  or (_01310_, _01309_, _01301_);
  or (_01311_, _01310_, _01299_);
  or (_01312_, _01311_, _01294_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01312_, _01275_);
  not (_01313_, _33596_);
  and (_01314_, _01121_, _01313_);
  not (_01315_, _33678_);
  and (_01316_, _01162_, _01315_);
  not (_01317_, _33637_);
  and (_01318_, _01117_, _01317_);
  or (_01319_, _01318_, _01316_);
  or (_01320_, _01319_, _01314_);
  not (_01321_, _33514_);
  and (_01322_, _01131_, _01321_);
  not (_01323_, _33555_);
  and (_01324_, _01142_, _01323_);
  not (_01325_, _33389_);
  and (_01326_, _01148_, _01325_);
  or (_01327_, _01326_, _01324_);
  and (_01328_, _01145_, _33951_);
  not (_01329_, _33726_);
  and (_01330_, _01138_, _01329_);
  or (_01331_, _01330_, _01328_);
  or (_01332_, _01331_, _01327_);
  or (_01333_, _01332_, _01322_);
  not (_01334_, _33473_);
  and (_01335_, _01127_, _01334_);
  not (_01336_, _33430_);
  and (_01337_, _01135_, _01336_);
  or (_01338_, _01337_, _01335_);
  or (_01339_, _01338_, _01333_);
  not (_01340_, _33327_);
  and (_01341_, _01158_, _01340_);
  not (_01342_, _33895_);
  and (_01343_, _01165_, _01342_);
  not (_01344_, _33837_);
  and (_01345_, _01168_, _01344_);
  or (_01346_, _01345_, _01343_);
  not (_01347_, _33781_);
  and (_01348_, _01171_, _01347_);
  or (_01349_, _01348_, _01346_);
  or (_01350_, _01349_, _01341_);
  not (_01351_, _33238_);
  and (_01352_, _01155_, _01351_);
  not (_01353_, _33279_);
  and (_01354_, _01113_, _01353_);
  or (_01355_, _01354_, _01352_);
  or (_01356_, _01355_, _01350_);
  or (_01357_, _01356_, _01339_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01357_, _01320_);
  not (_01358_, _33642_);
  and (_01359_, _01117_, _01358_);
  not (_01360_, _33683_);
  and (_01361_, _01162_, _01360_);
  not (_01362_, _33601_);
  and (_01363_, _01121_, _01362_);
  or (_01364_, _01363_, _01361_);
  or (_01365_, _01364_, _01359_);
  not (_01366_, _33478_);
  and (_01367_, _01127_, _01366_);
  not (_01368_, _33519_);
  and (_01369_, _01131_, _01368_);
  or (_01370_, _01369_, _01367_);
  not (_01371_, _33435_);
  and (_01372_, _01135_, _01371_);
  not (_01373_, _33560_);
  and (_01374_, _01142_, _01373_);
  not (_01375_, _33394_);
  and (_01376_, _01148_, _01375_);
  or (_01377_, _01376_, _01374_);
  and (_01378_, _01145_, _33958_);
  not (_01379_, _33732_);
  and (_01380_, _01138_, _01379_);
  or (_01381_, _01380_, _01378_);
  or (_01382_, _01381_, _01377_);
  or (_01383_, _01382_, _01372_);
  or (_01384_, _01383_, _01370_);
  not (_01385_, _33789_);
  and (_01386_, _01171_, _01385_);
  not (_01387_, _33844_);
  and (_01388_, _01168_, _01387_);
  not (_01389_, _33902_);
  and (_01390_, _01165_, _01389_);
  or (_01391_, _01390_, _01388_);
  or (_01392_, _01391_, _01386_);
  not (_01393_, _33338_);
  and (_01394_, _01158_, _01393_);
  or (_01395_, _01394_, _01392_);
  not (_01396_, _33243_);
  and (_01397_, _01155_, _01396_);
  not (_01398_, _33284_);
  and (_01399_, _01113_, _01398_);
  or (_01400_, _01399_, _01397_);
  or (_01401_, _01400_, _01395_);
  or (_01402_, _01401_, _01384_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01402_, _01365_);
  not (_01403_, _33647_);
  and (_01404_, _01117_, _01403_);
  not (_01405_, _33688_);
  and (_01406_, _01162_, _01405_);
  not (_01407_, _33606_);
  and (_01408_, _01121_, _01407_);
  or (_01409_, _01408_, _01406_);
  or (_01410_, _01409_, _01404_);
  not (_01411_, _33524_);
  and (_01412_, _01131_, _01411_);
  not (_01413_, _33565_);
  and (_01414_, _01142_, _01413_);
  not (_01415_, _33399_);
  and (_01416_, _01148_, _01415_);
  or (_01417_, _01416_, _01414_);
  and (_01418_, _01145_, _33965_);
  not (_01419_, _33739_);
  and (_01420_, _01138_, _01419_);
  or (_01421_, _01420_, _01418_);
  or (_01422_, _01421_, _01417_);
  or (_01423_, _01422_, _01412_);
  not (_01424_, _33483_);
  and (_01425_, _01127_, _01424_);
  not (_01426_, _33441_);
  and (_01427_, _01135_, _01426_);
  or (_01428_, _01427_, _01425_);
  or (_01429_, _01428_, _01423_);
  not (_01430_, _33795_);
  and (_01431_, _01171_, _01430_);
  not (_01432_, _33851_);
  and (_01433_, _01168_, _01432_);
  not (_01434_, _33909_);
  and (_01435_, _01165_, _01434_);
  or (_01436_, _01435_, _01433_);
  or (_01437_, _01436_, _01431_);
  not (_01438_, _33349_);
  and (_01439_, _01158_, _01438_);
  or (_01440_, _01439_, _01437_);
  not (_01441_, _33248_);
  and (_01442_, _01155_, _01441_);
  not (_01443_, _33289_);
  and (_01444_, _01113_, _01443_);
  or (_01445_, _01444_, _01442_);
  or (_01446_, _01445_, _01440_);
  or (_01447_, _01446_, _01429_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01447_, _01410_);
  not (_01448_, _33611_);
  and (_01449_, _01121_, _01448_);
  not (_01450_, _33652_);
  and (_01451_, _01117_, _01450_);
  not (_01452_, _33694_);
  and (_01453_, _01162_, _01452_);
  or (_01454_, _01453_, _01451_);
  or (_01455_, _01454_, _01449_);
  not (_01456_, _33802_);
  and (_01457_, _01171_, _01456_);
  not (_01458_, _33858_);
  and (_01459_, _01168_, _01458_);
  not (_01460_, _33916_);
  and (_01461_, _01165_, _01460_);
  or (_01462_, _01461_, _01459_);
  or (_01463_, _01462_, _01457_);
  not (_01464_, _33570_);
  and (_01465_, _01142_, _01464_);
  not (_01466_, _33746_);
  and (_01467_, _01138_, _01466_);
  or (_01468_, _01467_, _01465_);
  or (_01469_, _01468_, _01463_);
  or (_01470_, _01469_, _01455_);
  not (_01471_, _33294_);
  and (_01472_, _01113_, _01471_);
  not (_01473_, _33529_);
  and (_01474_, _01131_, _01473_);
  not (_01475_, _33488_);
  and (_01476_, _01127_, _01475_);
  or (_01477_, _01476_, _01474_);
  not (_01478_, _33404_);
  and (_01479_, _01148_, _01478_);
  not (_01480_, _33446_);
  and (_01481_, _01135_, _01480_);
  or (_01482_, _01481_, _01479_);
  or (_01483_, _01482_, _01477_);
  or (_01484_, _01483_, _01472_);
  and (_01485_, _01145_, _33972_);
  not (_01486_, _33360_);
  and (_01487_, _01158_, _01486_);
  not (_01488_, _33253_);
  and (_01489_, _01155_, _01488_);
  or (_01490_, _01489_, _01487_);
  or (_01491_, _01490_, _01485_);
  or (_01492_, _01491_, _01484_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01492_, _01470_);
  not (_01493_, _33616_);
  and (_01494_, _01121_, _01493_);
  not (_01495_, _33657_);
  and (_01496_, _01117_, _01495_);
  not (_01497_, _33700_);
  and (_01498_, _01162_, _01497_);
  or (_01499_, _01498_, _01496_);
  or (_01500_, _01499_, _01494_);
  not (_01501_, _33753_);
  and (_01502_, _01138_, _01501_);
  not (_01503_, _33923_);
  and (_01504_, _01165_, _01503_);
  not (_01505_, _33865_);
  and (_01506_, _01168_, _01505_);
  or (_01507_, _01506_, _01504_);
  or (_01508_, _01507_, _01502_);
  not (_01509_, _33575_);
  and (_01510_, _01142_, _01509_);
  not (_01511_, _33809_);
  and (_01512_, _01171_, _01511_);
  or (_01513_, _01512_, _01510_);
  or (_01514_, _01513_, _01508_);
  or (_01515_, _01514_, _01500_);
  not (_01516_, _33299_);
  and (_01517_, _01113_, _01516_);
  not (_01518_, _33534_);
  and (_01519_, _01131_, _01518_);
  not (_01520_, _33493_);
  and (_01521_, _01127_, _01520_);
  or (_01522_, _01521_, _01519_);
  not (_01523_, _33409_);
  and (_01524_, _01148_, _01523_);
  not (_01525_, _33452_);
  and (_01526_, _01135_, _01525_);
  or (_01527_, _01526_, _01524_);
  or (_01528_, _01527_, _01522_);
  or (_01529_, _01528_, _01517_);
  and (_01530_, _01145_, _33979_);
  not (_01531_, _33368_);
  and (_01532_, _01158_, _01531_);
  not (_01533_, _33258_);
  and (_01534_, _01155_, _01533_);
  or (_01535_, _01534_, _01532_);
  or (_01536_, _01535_, _01530_);
  or (_01537_, _01536_, _01529_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01537_, _01515_);
  not (_01538_, _33621_);
  and (_01539_, _01121_, _01538_);
  not (_01540_, _33373_);
  and (_01541_, _01158_, _01540_);
  not (_01542_, _33706_);
  and (_01543_, _01162_, _01542_);
  or (_01544_, _01543_, _01541_);
  or (_01545_, _01544_, _01539_);
  not (_01546_, _33539_);
  and (_01547_, _01131_, _01546_);
  not (_01548_, _33414_);
  and (_01549_, _01148_, _01548_);
  not (_01550_, _33580_);
  and (_01551_, _01142_, _01550_);
  or (_01552_, _01551_, _01549_);
  and (_01553_, _01145_, _33986_);
  not (_01554_, _33760_);
  and (_01555_, _01138_, _01554_);
  or (_01556_, _01555_, _01553_);
  or (_01557_, _01556_, _01552_);
  or (_01558_, _01557_, _01547_);
  not (_01559_, _33498_);
  and (_01560_, _01127_, _01559_);
  not (_01561_, _33457_);
  and (_01562_, _01135_, _01561_);
  or (_01563_, _01562_, _01560_);
  or (_01564_, _01563_, _01558_);
  not (_01565_, _33662_);
  and (_01566_, _01117_, _01565_);
  not (_01567_, _33930_);
  and (_01568_, _01165_, _01567_);
  not (_01569_, _33872_);
  and (_01570_, _01168_, _01569_);
  not (_01571_, _33816_);
  and (_01572_, _01171_, _01571_);
  or (_01573_, _01572_, _01570_);
  or (_01574_, _01573_, _01568_);
  or (_01575_, _01574_, _01566_);
  not (_01576_, _33263_);
  and (_01577_, _01155_, _01576_);
  not (_01578_, _33304_);
  and (_01579_, _01113_, _01578_);
  or (_01580_, _01579_, _01577_);
  or (_01581_, _01580_, _01575_);
  or (_01582_, _01581_, _01564_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01582_, _01545_);
  and (_01583_, _01117_, _01285_);
  and (_01584_, _01113_, _33944_);
  and (_01585_, _01158_, _01295_);
  or (_01586_, _01585_, _01584_);
  or (_01587_, _01586_, _01583_);
  and (_01588_, _01127_, _01289_);
  and (_01589_, _01138_, _01272_);
  and (_01590_, _01145_, _01302_);
  or (_01591_, _01590_, _01589_);
  and (_01592_, _01142_, _01276_);
  and (_01593_, _01148_, _01268_);
  or (_01594_, _01593_, _01592_);
  or (_01595_, _01594_, _01591_);
  or (_01596_, _01595_, _01588_);
  and (_01597_, _01131_, _01281_);
  and (_01598_, _01135_, _01297_);
  or (_01599_, _01598_, _01597_);
  or (_01600_, _01599_, _01596_);
  and (_01601_, _01162_, _01300_);
  and (_01602_, _01171_, _01270_);
  and (_01603_, _01165_, _01306_);
  and (_01604_, _01168_, _01283_);
  or (_01605_, _01604_, _01603_);
  or (_01606_, _01605_, _01602_);
  or (_01607_, _01606_, _01601_);
  and (_01608_, _01155_, _01304_);
  and (_01609_, _01121_, _01278_);
  or (_01610_, _01609_, _01608_);
  or (_01611_, _01610_, _01607_);
  or (_01612_, _01611_, _01600_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01612_, _01587_);
  and (_01613_, _01117_, _01323_);
  and (_01614_, _01113_, _33951_);
  and (_01615_, _01158_, _01351_);
  or (_01616_, _01615_, _01614_);
  or (_01617_, _01616_, _01613_);
  and (_01618_, _01127_, _01325_);
  and (_01619_, _01142_, _01334_);
  and (_01620_, _01148_, _01353_);
  or (_01621_, _01620_, _01619_);
  and (_01622_, _01138_, _01317_);
  and (_01623_, _01145_, _01344_);
  or (_01624_, _01623_, _01622_);
  or (_01625_, _01624_, _01621_);
  or (_01626_, _01625_, _01618_);
  and (_01627_, _01131_, _01336_);
  and (_01628_, _01135_, _01340_);
  or (_01629_, _01628_, _01627_);
  or (_01630_, _01629_, _01626_);
  and (_01631_, _01162_, _01313_);
  and (_01632_, _01168_, _01329_);
  and (_01633_, _01171_, _01315_);
  and (_01634_, _01165_, _01347_);
  or (_01635_, _01634_, _01633_);
  or (_01636_, _01635_, _01632_);
  or (_01637_, _01636_, _01631_);
  and (_01638_, _01155_, _01342_);
  and (_01639_, _01121_, _01321_);
  or (_01640_, _01639_, _01638_);
  or (_01641_, _01640_, _01637_);
  or (_01642_, _01641_, _01630_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01642_, _01617_);
  and (_01643_, _01168_, _01379_);
  and (_01644_, _01165_, _01385_);
  or (_01645_, _01644_, _01643_);
  and (_01646_, _01155_, _01389_);
  or (_01647_, _01646_, _01645_);
  and (_01648_, _01162_, _01362_);
  and (_01649_, _01113_, _33958_);
  or (_01650_, _01649_, _01648_);
  or (_01651_, _01650_, _01647_);
  and (_01652_, _01142_, _01366_);
  and (_01653_, _01127_, _01375_);
  and (_01654_, _01131_, _01371_);
  or (_01655_, _01654_, _01653_);
  or (_01656_, _01655_, _01652_);
  and (_01657_, _01148_, _01398_);
  and (_01658_, _01121_, _01368_);
  or (_01659_, _01658_, _01657_);
  or (_01660_, _01659_, _01656_);
  or (_01661_, _01660_, _01651_);
  and (_01662_, _01145_, _01387_);
  and (_01663_, _01158_, _01396_);
  and (_01664_, _01135_, _01393_);
  or (_01665_, _01664_, _01663_);
  and (_01666_, _01117_, _01373_);
  and (_01667_, _01138_, _01358_);
  and (_01668_, _01171_, _01360_);
  or (_01669_, _01668_, _01667_);
  or (_01670_, _01669_, _01666_);
  or (_01671_, _01670_, _01665_);
  or (_01672_, _01671_, _01662_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01672_, _01661_);
  and (_01673_, _01162_, _01407_);
  and (_01674_, _01117_, _01413_);
  and (_01675_, _01158_, _01441_);
  or (_01676_, _01675_, _01674_);
  or (_01677_, _01676_, _01673_);
  and (_01678_, _01127_, _01415_);
  and (_01679_, _01131_, _01426_);
  or (_01680_, _01679_, _01678_);
  and (_01681_, _01135_, _01438_);
  and (_01682_, _01138_, _01403_);
  and (_01683_, _01145_, _01432_);
  or (_01684_, _01683_, _01682_);
  and (_01685_, _01148_, _01443_);
  and (_01686_, _01142_, _01424_);
  or (_01687_, _01686_, _01685_);
  or (_01688_, _01687_, _01684_);
  or (_01689_, _01688_, _01681_);
  or (_01690_, _01689_, _01680_);
  and (_01691_, _01121_, _01411_);
  and (_01692_, _01165_, _01430_);
  and (_01693_, _01171_, _01405_);
  and (_01694_, _01168_, _01419_);
  or (_01695_, _01694_, _01693_);
  or (_01696_, _01695_, _01692_);
  or (_01697_, _01696_, _01691_);
  and (_01698_, _01113_, _33965_);
  and (_01699_, _01155_, _01434_);
  or (_01700_, _01699_, _01698_);
  or (_01701_, _01700_, _01697_);
  or (_01702_, _01701_, _01690_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01702_, _01677_);
  and (_01703_, _01168_, _01466_);
  and (_01704_, _01165_, _01456_);
  or (_01705_, _01704_, _01703_);
  and (_01706_, _01155_, _01460_);
  or (_01707_, _01706_, _01705_);
  and (_01708_, _01162_, _01448_);
  and (_01709_, _01113_, _33972_);
  or (_01710_, _01709_, _01708_);
  or (_01711_, _01710_, _01707_);
  and (_01712_, _01142_, _01475_);
  and (_01713_, _01127_, _01478_);
  and (_01714_, _01131_, _01480_);
  or (_01715_, _01714_, _01713_);
  or (_01716_, _01715_, _01712_);
  and (_01717_, _01148_, _01471_);
  and (_01718_, _01121_, _01473_);
  or (_01719_, _01718_, _01717_);
  or (_01720_, _01719_, _01716_);
  or (_01721_, _01720_, _01711_);
  and (_01722_, _01145_, _01458_);
  and (_01723_, _01158_, _01488_);
  and (_01724_, _01135_, _01486_);
  or (_01725_, _01724_, _01723_);
  and (_01726_, _01117_, _01464_);
  and (_01727_, _01138_, _01450_);
  and (_01728_, _01171_, _01452_);
  or (_01729_, _01728_, _01727_);
  or (_01730_, _01729_, _01726_);
  or (_01731_, _01730_, _01725_);
  or (_01732_, _01731_, _01722_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01732_, _01721_);
  and (_01733_, _01168_, _01501_);
  and (_01734_, _01165_, _01511_);
  or (_01735_, _01734_, _01733_);
  and (_01736_, _01155_, _01503_);
  or (_01737_, _01736_, _01735_);
  and (_01738_, _01162_, _01493_);
  and (_01739_, _01113_, _33979_);
  or (_01740_, _01739_, _01738_);
  or (_01741_, _01740_, _01737_);
  and (_01742_, _01142_, _01520_);
  and (_01743_, _01127_, _01523_);
  and (_01744_, _01131_, _01525_);
  or (_01745_, _01744_, _01743_);
  or (_01746_, _01745_, _01742_);
  and (_01747_, _01148_, _01516_);
  and (_01748_, _01121_, _01518_);
  or (_01749_, _01748_, _01747_);
  or (_01750_, _01749_, _01746_);
  or (_01751_, _01750_, _01741_);
  and (_01752_, _01145_, _01505_);
  and (_01753_, _01158_, _01533_);
  and (_01754_, _01135_, _01531_);
  or (_01755_, _01754_, _01753_);
  and (_01756_, _01117_, _01509_);
  and (_01757_, _01138_, _01495_);
  and (_01758_, _01171_, _01497_);
  or (_01759_, _01758_, _01757_);
  or (_01760_, _01759_, _01756_);
  or (_01761_, _01760_, _01755_);
  or (_01762_, _01761_, _01752_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01762_, _01751_);
  and (_01763_, _01117_, _01550_);
  and (_01764_, _01155_, _01567_);
  and (_01765_, _01158_, _01576_);
  or (_01766_, _01765_, _01764_);
  or (_01767_, _01766_, _01763_);
  and (_01768_, _01127_, _01548_);
  and (_01769_, _01131_, _01561_);
  or (_01770_, _01769_, _01768_);
  and (_01771_, _01135_, _01540_);
  and (_01772_, _01145_, _01569_);
  and (_01773_, _01148_, _01578_);
  or (_01774_, _01773_, _01772_);
  and (_01775_, _01138_, _01565_);
  and (_01776_, _01142_, _01559_);
  or (_01777_, _01776_, _01775_);
  or (_01778_, _01777_, _01774_);
  or (_01779_, _01778_, _01771_);
  or (_01780_, _01779_, _01770_);
  and (_01781_, _01113_, _33986_);
  and (_01782_, _01162_, _01538_);
  or (_01783_, _01782_, _01781_);
  and (_01784_, _01121_, _01546_);
  and (_01785_, _01168_, _01554_);
  and (_01786_, _01165_, _01571_);
  and (_01787_, _01171_, _01542_);
  or (_01788_, _01787_, _01786_);
  or (_01789_, _01788_, _01785_);
  or (_01790_, _01789_, _01784_);
  or (_01791_, _01790_, _01783_);
  or (_01792_, _01791_, _01780_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01792_, _01767_);
  and (_01793_, _01155_, _33944_);
  and (_01794_, _01162_, _01272_);
  and (_01795_, _01117_, _01300_);
  or (_01796_, _01795_, _01794_);
  or (_01797_, _01796_, _01793_);
  and (_01798_, _01135_, _01289_);
  and (_01799_, _01138_, _01270_);
  and (_01800_, _01142_, _01278_);
  or (_01801_, _01800_, _01799_);
  and (_01802_, _01145_, _01304_);
  and (_01803_, _01148_, _01297_);
  or (_01804_, _01803_, _01802_);
  or (_01805_, _01804_, _01801_);
  or (_01806_, _01805_, _01798_);
  and (_01807_, _01131_, _01276_);
  and (_01808_, _01127_, _01281_);
  or (_01809_, _01808_, _01807_);
  or (_01810_, _01809_, _01806_);
  and (_01811_, _01113_, _01295_);
  and (_01812_, _01165_, _01302_);
  and (_01813_, _01171_, _01283_);
  and (_01814_, _01168_, _01306_);
  or (_01815_, _01814_, _01813_);
  or (_01816_, _01815_, _01812_);
  or (_01817_, _01816_, _01811_);
  and (_01818_, _01121_, _01285_);
  and (_01819_, _01158_, _01268_);
  or (_01820_, _01819_, _01818_);
  or (_01821_, _01820_, _01817_);
  or (_01822_, _01821_, _01810_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01822_, _01797_);
  and (_01823_, _01155_, _33951_);
  and (_01824_, _01162_, _01317_);
  and (_01825_, _01121_, _01323_);
  or (_01826_, _01825_, _01824_);
  or (_01827_, _01826_, _01823_);
  and (_01828_, _01135_, _01325_);
  and (_01829_, _01138_, _01315_);
  and (_01830_, _01142_, _01321_);
  or (_01831_, _01830_, _01829_);
  and (_01832_, _01145_, _01342_);
  and (_01833_, _01148_, _01340_);
  or (_01834_, _01833_, _01832_);
  or (_01835_, _01834_, _01831_);
  or (_01836_, _01835_, _01828_);
  and (_01837_, _01131_, _01334_);
  and (_01838_, _01127_, _01336_);
  or (_01839_, _01838_, _01837_);
  or (_01840_, _01839_, _01836_);
  and (_01841_, _01113_, _01351_);
  and (_01842_, _01165_, _01344_);
  and (_01843_, _01171_, _01329_);
  and (_01844_, _01168_, _01347_);
  or (_01845_, _01844_, _01843_);
  or (_01846_, _01845_, _01842_);
  or (_01847_, _01846_, _01841_);
  and (_01848_, _01117_, _01313_);
  and (_01849_, _01158_, _01353_);
  or (_01850_, _01849_, _01848_);
  or (_01851_, _01850_, _01847_);
  or (_01852_, _01851_, _01840_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01852_, _01827_);
  and (_01853_, _01162_, _01358_);
  and (_01854_, _01155_, _33958_);
  and (_01855_, _01113_, _01396_);
  or (_01856_, _01855_, _01854_);
  or (_01857_, _01856_, _01853_);
  and (_01858_, _01127_, _01371_);
  and (_01859_, _01142_, _01368_);
  and (_01860_, _01148_, _01393_);
  or (_01861_, _01860_, _01859_);
  and (_01862_, _01145_, _01389_);
  and (_01863_, _01138_, _01360_);
  or (_01864_, _01863_, _01862_);
  or (_01865_, _01864_, _01861_);
  or (_01866_, _01865_, _01858_);
  and (_01867_, _01131_, _01366_);
  and (_01868_, _01135_, _01375_);
  or (_01869_, _01868_, _01867_);
  or (_01870_, _01869_, _01866_);
  and (_01871_, _01117_, _01362_);
  and (_01872_, _01165_, _01387_);
  and (_01873_, _01168_, _01385_);
  and (_01874_, _01171_, _01379_);
  or (_01875_, _01874_, _01873_);
  or (_01876_, _01875_, _01872_);
  or (_01877_, _01876_, _01871_);
  and (_01878_, _01158_, _01398_);
  and (_01879_, _01121_, _01373_);
  or (_01880_, _01879_, _01878_);
  or (_01881_, _01880_, _01877_);
  or (_01882_, _01881_, _01870_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01882_, _01857_);
  and (_01883_, _01162_, _01403_);
  and (_01884_, _01155_, _33965_);
  and (_01885_, _01113_, _01441_);
  or (_01886_, _01885_, _01884_);
  or (_01887_, _01886_, _01883_);
  and (_01888_, _01127_, _01426_);
  and (_01889_, _01142_, _01411_);
  and (_01890_, _01148_, _01438_);
  or (_01891_, _01890_, _01889_);
  and (_01892_, _01145_, _01434_);
  and (_01893_, _01138_, _01405_);
  or (_01894_, _01893_, _01892_);
  or (_01895_, _01894_, _01891_);
  or (_01896_, _01895_, _01888_);
  and (_01897_, _01131_, _01424_);
  and (_01898_, _01135_, _01415_);
  or (_01899_, _01898_, _01897_);
  or (_01900_, _01899_, _01896_);
  and (_01901_, _01117_, _01407_);
  and (_01902_, _01165_, _01432_);
  and (_01903_, _01168_, _01430_);
  and (_01904_, _01171_, _01419_);
  or (_01905_, _01904_, _01903_);
  or (_01906_, _01905_, _01902_);
  or (_01907_, _01906_, _01901_);
  and (_01908_, _01158_, _01443_);
  and (_01909_, _01121_, _01413_);
  or (_01910_, _01909_, _01908_);
  or (_01911_, _01910_, _01907_);
  or (_01912_, _01911_, _01900_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01912_, _01887_);
  and (_01913_, _01162_, _01450_);
  and (_01914_, _01113_, _01488_);
  and (_01915_, _01117_, _01448_);
  or (_01916_, _01915_, _01914_);
  or (_01917_, _01916_, _01913_);
  and (_01918_, _01127_, _01480_);
  and (_01919_, _01142_, _01473_);
  and (_01920_, _01148_, _01486_);
  or (_01921_, _01920_, _01919_);
  and (_01922_, _01138_, _01452_);
  and (_01923_, _01145_, _01460_);
  or (_01924_, _01923_, _01922_);
  or (_01925_, _01924_, _01921_);
  or (_01926_, _01925_, _01918_);
  and (_01927_, _01131_, _01475_);
  and (_01928_, _01135_, _01478_);
  or (_01929_, _01928_, _01927_);
  or (_01930_, _01929_, _01926_);
  and (_01931_, _01121_, _01464_);
  and (_01932_, _01165_, _01458_);
  and (_01933_, _01168_, _01456_);
  and (_01934_, _01171_, _01466_);
  or (_01935_, _01934_, _01933_);
  or (_01936_, _01935_, _01932_);
  or (_01937_, _01936_, _01931_);
  and (_01938_, _01155_, _33972_);
  and (_01939_, _01158_, _01471_);
  or (_01940_, _01939_, _01938_);
  or (_01941_, _01940_, _01937_);
  or (_01942_, _01941_, _01930_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01942_, _01917_);
  and (_01943_, _01162_, _01495_);
  and (_01944_, _01155_, _33979_);
  and (_01945_, _01113_, _01533_);
  or (_01946_, _01945_, _01944_);
  or (_01947_, _01946_, _01943_);
  and (_01948_, _01127_, _01525_);
  and (_01949_, _01142_, _01518_);
  and (_01950_, _01148_, _01531_);
  or (_01951_, _01950_, _01949_);
  and (_01952_, _01145_, _01503_);
  and (_01953_, _01138_, _01497_);
  or (_01954_, _01953_, _01952_);
  or (_01955_, _01954_, _01951_);
  or (_01956_, _01955_, _01948_);
  and (_01957_, _01131_, _01520_);
  and (_01958_, _01135_, _01523_);
  or (_01959_, _01958_, _01957_);
  or (_01960_, _01959_, _01956_);
  and (_01961_, _01117_, _01493_);
  and (_01962_, _01165_, _01505_);
  and (_01963_, _01168_, _01511_);
  and (_01964_, _01171_, _01501_);
  or (_01965_, _01964_, _01963_);
  or (_01966_, _01965_, _01962_);
  or (_01967_, _01966_, _01961_);
  and (_01968_, _01158_, _01516_);
  and (_01969_, _01121_, _01509_);
  or (_01970_, _01969_, _01968_);
  or (_01971_, _01970_, _01967_);
  or (_01972_, _01971_, _01960_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01972_, _01947_);
  and (_01973_, _01162_, _01565_);
  and (_01974_, _01113_, _01576_);
  and (_01975_, _01117_, _01538_);
  or (_01976_, _01975_, _01974_);
  or (_01977_, _01976_, _01973_);
  and (_01978_, _01127_, _01561_);
  and (_01979_, _01142_, _01546_);
  and (_01980_, _01148_, _01540_);
  or (_01981_, _01980_, _01979_);
  and (_01982_, _01138_, _01542_);
  and (_01983_, _01145_, _01567_);
  or (_01984_, _01983_, _01982_);
  or (_01985_, _01984_, _01981_);
  or (_01986_, _01985_, _01978_);
  and (_01987_, _01131_, _01559_);
  and (_01988_, _01135_, _01548_);
  or (_01989_, _01988_, _01987_);
  or (_01990_, _01989_, _01986_);
  and (_01991_, _01121_, _01550_);
  and (_01992_, _01165_, _01569_);
  and (_01993_, _01168_, _01571_);
  and (_01994_, _01171_, _01554_);
  or (_01995_, _01994_, _01993_);
  or (_01996_, _01995_, _01992_);
  or (_01997_, _01996_, _01991_);
  and (_01998_, _01155_, _33986_);
  and (_01999_, _01158_, _01578_);
  or (_02000_, _01999_, _01998_);
  or (_02001_, _02000_, _01997_);
  or (_02002_, _02001_, _01990_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02002_, _01977_);
  and (_02003_, _01113_, _01304_);
  and (_02004_, _01117_, _01278_);
  and (_02005_, _01121_, _01276_);
  or (_02006_, _02005_, _02004_);
  or (_02007_, _02006_, _02003_);
  and (_02008_, _01127_, _01297_);
  and (_02009_, _01145_, _01306_);
  and (_02010_, _01142_, _01281_);
  or (_02011_, _02010_, _02009_);
  and (_02012_, _01138_, _01300_);
  and (_02013_, _01148_, _01295_);
  or (_02014_, _02013_, _02012_);
  or (_02015_, _02014_, _02011_);
  or (_02016_, _02015_, _02008_);
  and (_02017_, _01135_, _01268_);
  and (_02018_, _01131_, _01289_);
  or (_02019_, _02018_, _02017_);
  or (_02020_, _02019_, _02016_);
  and (_02021_, _01162_, _01285_);
  and (_02022_, _01171_, _01272_);
  and (_02023_, _01165_, _01283_);
  and (_02024_, _01168_, _01270_);
  or (_02025_, _02024_, _02023_);
  or (_02026_, _02025_, _02022_);
  or (_02027_, _02026_, _02021_);
  and (_02028_, _01158_, _33944_);
  and (_02029_, _01155_, _01302_);
  or (_02030_, _02029_, _02028_);
  or (_02031_, _02030_, _02027_);
  or (_02032_, _02031_, _02020_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02032_, _02007_);
  and (_02033_, _01162_, _01323_);
  and (_02034_, _01121_, _01334_);
  and (_02035_, _01155_, _01344_);
  or (_02036_, _02035_, _02034_);
  or (_02037_, _02036_, _02033_);
  and (_02038_, _01127_, _01340_);
  and (_02039_, _01135_, _01353_);
  or (_02040_, _02039_, _02038_);
  and (_02041_, _01131_, _01325_);
  and (_02042_, _01148_, _01351_);
  and (_02043_, _01142_, _01336_);
  or (_02044_, _02043_, _02042_);
  and (_02045_, _01138_, _01313_);
  and (_02046_, _01145_, _01347_);
  or (_02047_, _02046_, _02045_);
  or (_02048_, _02047_, _02044_);
  or (_02049_, _02048_, _02041_);
  or (_02050_, _02049_, _02040_);
  and (_02051_, _01158_, _33951_);
  and (_02052_, _01168_, _01315_);
  and (_02053_, _01171_, _01317_);
  or (_02054_, _02053_, _02052_);
  and (_02055_, _01165_, _01329_);
  or (_02056_, _02055_, _02054_);
  or (_02057_, _02056_, _02051_);
  and (_02058_, _01117_, _01321_);
  and (_02059_, _01113_, _01342_);
  or (_02060_, _02059_, _02058_);
  or (_02061_, _02060_, _02057_);
  or (_02062_, _02061_, _02050_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02062_, _02037_);
  and (_02063_, _01155_, _01387_);
  and (_02064_, _01162_, _01373_);
  and (_02065_, _01121_, _01366_);
  or (_02066_, _02065_, _02064_);
  or (_02067_, _02066_, _02063_);
  and (_02068_, _01135_, _01398_);
  and (_02069_, _01145_, _01385_);
  and (_02070_, _01142_, _01371_);
  or (_02071_, _02070_, _02069_);
  and (_02072_, _01138_, _01362_);
  and (_02073_, _01148_, _01396_);
  or (_02074_, _02073_, _02072_);
  or (_02075_, _02074_, _02071_);
  or (_02076_, _02075_, _02068_);
  and (_02077_, _01127_, _01393_);
  and (_02078_, _01131_, _01375_);
  or (_02079_, _02078_, _02077_);
  or (_02080_, _02079_, _02076_);
  and (_02081_, _01158_, _33958_);
  and (_02082_, _01113_, _01389_);
  or (_02083_, _02082_, _02081_);
  and (_02084_, _01117_, _01368_);
  and (_02085_, _01168_, _01360_);
  and (_02086_, _01165_, _01379_);
  and (_02087_, _01171_, _01358_);
  or (_02088_, _02087_, _02086_);
  or (_02089_, _02088_, _02085_);
  or (_02090_, _02089_, _02084_);
  or (_02091_, _02090_, _02083_);
  or (_02092_, _02091_, _02080_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02092_, _02067_);
  and (_02093_, _01162_, _01413_);
  and (_02094_, _01155_, _01432_);
  and (_02095_, _01121_, _01424_);
  or (_02096_, _02095_, _02094_);
  or (_02097_, _02096_, _02093_);
  and (_02098_, _01127_, _01438_);
  and (_02099_, _01145_, _01430_);
  and (_02100_, _01142_, _01426_);
  or (_02101_, _02100_, _02099_);
  and (_02102_, _01138_, _01407_);
  and (_02103_, _01148_, _01441_);
  or (_02104_, _02103_, _02102_);
  or (_02105_, _02104_, _02101_);
  or (_02106_, _02105_, _02098_);
  and (_02107_, _01135_, _01443_);
  and (_02108_, _01131_, _01415_);
  or (_02109_, _02108_, _02107_);
  or (_02110_, _02109_, _02106_);
  and (_02111_, _01158_, _33965_);
  and (_02112_, _01113_, _01434_);
  or (_02113_, _02112_, _02111_);
  and (_02114_, _01117_, _01411_);
  and (_02115_, _01168_, _01405_);
  and (_02116_, _01165_, _01419_);
  and (_02117_, _01171_, _01403_);
  or (_02118_, _02117_, _02116_);
  or (_02119_, _02118_, _02115_);
  or (_02120_, _02119_, _02114_);
  or (_02121_, _02120_, _02113_);
  or (_02122_, _02121_, _02110_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02122_, _02097_);
  and (_02123_, _01113_, _01460_);
  and (_02124_, _01162_, _01464_);
  and (_02125_, _01121_, _01475_);
  or (_02126_, _02125_, _02124_);
  or (_02127_, _02126_, _02123_);
  and (_02128_, _01127_, _01486_);
  and (_02129_, _01145_, _01456_);
  and (_02130_, _01142_, _01480_);
  or (_02131_, _02130_, _02129_);
  and (_02132_, _01138_, _01448_);
  and (_02133_, _01148_, _01488_);
  or (_02134_, _02133_, _02132_);
  or (_02135_, _02134_, _02131_);
  or (_02136_, _02135_, _02128_);
  and (_02137_, _01135_, _01471_);
  and (_02138_, _01131_, _01478_);
  or (_02139_, _02138_, _02137_);
  or (_02140_, _02139_, _02136_);
  and (_02141_, _01117_, _01473_);
  and (_02142_, _01171_, _01450_);
  and (_02143_, _01165_, _01466_);
  and (_02144_, _01168_, _01452_);
  or (_02145_, _02144_, _02143_);
  or (_02146_, _02145_, _02142_);
  or (_02147_, _02146_, _02141_);
  and (_02148_, _01158_, _33972_);
  and (_02149_, _01155_, _01458_);
  or (_02150_, _02149_, _02148_);
  or (_02151_, _02150_, _02147_);
  or (_02152_, _02151_, _02140_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02152_, _02127_);
  and (_02153_, _01162_, _01509_);
  and (_02154_, _01155_, _01505_);
  and (_02155_, _01121_, _01520_);
  or (_02156_, _02155_, _02154_);
  or (_02157_, _02156_, _02153_);
  and (_02158_, _01127_, _01531_);
  and (_02159_, _01145_, _01511_);
  and (_02160_, _01142_, _01525_);
  or (_02161_, _02160_, _02159_);
  and (_02162_, _01138_, _01493_);
  and (_02163_, _01148_, _01533_);
  or (_02164_, _02163_, _02162_);
  or (_02165_, _02164_, _02161_);
  or (_02166_, _02165_, _02158_);
  and (_02167_, _01135_, _01516_);
  and (_02168_, _01131_, _01523_);
  or (_02169_, _02168_, _02167_);
  or (_02170_, _02169_, _02166_);
  and (_02171_, _01158_, _33979_);
  and (_02172_, _01113_, _01503_);
  or (_02173_, _02172_, _02171_);
  and (_02174_, _01117_, _01518_);
  and (_02175_, _01168_, _01497_);
  and (_02176_, _01165_, _01501_);
  and (_02177_, _01171_, _01495_);
  or (_02178_, _02177_, _02176_);
  or (_02179_, _02178_, _02175_);
  or (_02180_, _02179_, _02174_);
  or (_02181_, _02180_, _02173_);
  or (_02182_, _02181_, _02170_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02182_, _02157_);
  and (_02183_, _01162_, _01550_);
  and (_02184_, _01158_, _33986_);
  and (_02185_, _01121_, _01559_);
  or (_02186_, _02185_, _02184_);
  or (_02187_, _02186_, _02183_);
  and (_02188_, _01127_, _01540_);
  and (_02189_, _01148_, _01576_);
  and (_02190_, _01138_, _01538_);
  or (_02191_, _02190_, _02189_);
  and (_02192_, _01142_, _01561_);
  and (_02193_, _01145_, _01571_);
  or (_02194_, _02193_, _02192_);
  or (_02195_, _02194_, _02191_);
  or (_02196_, _02195_, _02188_);
  and (_02197_, _01135_, _01578_);
  and (_02198_, _01131_, _01548_);
  or (_02199_, _02198_, _02197_);
  or (_02200_, _02199_, _02196_);
  and (_02201_, _01113_, _01567_);
  and (_02202_, _01171_, _01565_);
  and (_02203_, _01168_, _01542_);
  and (_02204_, _01165_, _01554_);
  or (_02205_, _02204_, _02203_);
  or (_02206_, _02205_, _02202_);
  or (_02207_, _02206_, _02201_);
  and (_02208_, _01117_, _01546_);
  and (_02209_, _01155_, _01569_);
  or (_02210_, _02209_, _02208_);
  or (_02211_, _02210_, _02207_);
  or (_02212_, _02211_, _02200_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02212_, _02187_);
  nand (_02213_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02214_, \oc8051_golden_model_1.PC [3]);
  or (_02215_, \oc8051_golden_model_1.PC [2], _02214_);
  or (_02216_, _02215_, _02213_);
  or (_02217_, _02216_, _33760_);
  not (_02218_, \oc8051_golden_model_1.PC [1]);
  or (_02219_, _02218_, \oc8051_golden_model_1.PC [0]);
  or (_02220_, _02219_, _02215_);
  or (_02221_, _02220_, _33706_);
  and (_02222_, _02221_, _02217_);
  not (_02223_, \oc8051_golden_model_1.PC [2]);
  or (_02224_, _02223_, \oc8051_golden_model_1.PC [3]);
  or (_02225_, _02224_, _02213_);
  or (_02226_, _02225_, _33580_);
  or (_02227_, _02224_, _02219_);
  or (_02228_, _02227_, _33539_);
  and (_02229_, _02228_, _02226_);
  and (_02230_, _02229_, _02222_);
  and (_02231_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_02232_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_02233_, _02232_, _02231_);
  nand (_02234_, _02233_, _33986_);
  nand (_02235_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02236_, _02235_, _02219_);
  or (_02237_, _02236_, _33930_);
  and (_02238_, _02237_, _02234_);
  or (_02239_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02240_, _02239_, _02213_);
  or (_02241_, _02240_, _33414_);
  or (_02242_, _02239_, _02219_);
  or (_02243_, _02242_, _33373_);
  and (_02244_, _02243_, _02241_);
  and (_02245_, _02244_, _02238_);
  and (_02246_, _02245_, _02230_);
  not (_02247_, \oc8051_golden_model_1.PC [0]);
  or (_02248_, \oc8051_golden_model_1.PC [1], _02247_);
  or (_02249_, _02248_, _02235_);
  or (_02250_, _02249_, _33872_);
  or (_02251_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02252_, _02251_, _02235_);
  or (_02253_, _02252_, _33816_);
  and (_02254_, _02253_, _02250_);
  or (_02255_, _02239_, _02251_);
  or (_02256_, _02255_, _33263_);
  or (_02257_, _02239_, _02248_);
  or (_02258_, _02257_, _33304_);
  and (_02259_, _02258_, _02256_);
  and (_02260_, _02259_, _02254_);
  or (_02261_, _02248_, _02215_);
  or (_02262_, _02261_, _33662_);
  or (_02263_, _02251_, _02215_);
  or (_02264_, _02263_, _33621_);
  and (_02265_, _02264_, _02262_);
  or (_02266_, _02248_, _02224_);
  or (_02267_, _02266_, _33498_);
  or (_02268_, _02251_, _02224_);
  or (_02269_, _02268_, _33457_);
  and (_02270_, _02269_, _02267_);
  and (_02271_, _02270_, _02265_);
  and (_02272_, _02271_, _02260_);
  and (_02273_, _02272_, _02246_);
  or (_02274_, _02216_, _33713_);
  or (_02275_, _02220_, _33668_);
  and (_02276_, _02275_, _02274_);
  or (_02277_, _02225_, _33545_);
  or (_02278_, _02227_, _33504_);
  and (_02279_, _02278_, _02277_);
  and (_02280_, _02279_, _02276_);
  nand (_02281_, _02233_, _33937_);
  or (_02282_, _02236_, _33881_);
  and (_02283_, _02282_, _02281_);
  or (_02284_, _02240_, _33379_);
  or (_02285_, _02242_, _33310_);
  and (_02286_, _02285_, _02284_);
  and (_02287_, _02286_, _02283_);
  and (_02288_, _02287_, _02280_);
  or (_02289_, _02249_, _33823_);
  or (_02290_, _02252_, _33767_);
  and (_02291_, _02290_, _02289_);
  or (_02292_, _02255_, _33228_);
  or (_02293_, _02257_, _33269_);
  and (_02294_, _02293_, _02292_);
  and (_02295_, _02294_, _02291_);
  or (_02296_, _02261_, _33627_);
  or (_02297_, _02263_, _33586_);
  and (_02298_, _02297_, _02296_);
  or (_02299_, _02266_, _33463_);
  or (_02300_, _02268_, _33420_);
  and (_02301_, _02300_, _02299_);
  and (_02302_, _02301_, _02298_);
  and (_02303_, _02302_, _02295_);
  and (_02304_, _02303_, _02288_);
  and (_02305_, _02304_, _02273_);
  or (_02306_, _02216_, _33746_);
  or (_02307_, _02220_, _33694_);
  and (_02308_, _02307_, _02306_);
  or (_02309_, _02225_, _33570_);
  or (_02310_, _02227_, _33529_);
  and (_02311_, _02310_, _02309_);
  and (_02312_, _02311_, _02308_);
  nand (_02313_, _02233_, _33972_);
  or (_02314_, _02236_, _33916_);
  and (_02315_, _02314_, _02313_);
  or (_02316_, _02240_, _33404_);
  or (_02317_, _02242_, _33360_);
  and (_02318_, _02317_, _02316_);
  and (_02319_, _02318_, _02315_);
  and (_02320_, _02319_, _02312_);
  or (_02321_, _02249_, _33858_);
  or (_02322_, _02252_, _33802_);
  and (_02323_, _02322_, _02321_);
  or (_02324_, _02255_, _33253_);
  or (_02325_, _02257_, _33294_);
  and (_02326_, _02325_, _02324_);
  and (_02327_, _02326_, _02323_);
  or (_02328_, _02261_, _33652_);
  or (_02329_, _02263_, _33611_);
  and (_02330_, _02329_, _02328_);
  or (_02331_, _02266_, _33488_);
  or (_02332_, _02268_, _33446_);
  and (_02333_, _02332_, _02331_);
  and (_02334_, _02333_, _02330_);
  and (_02335_, _02334_, _02327_);
  and (_02336_, _02335_, _02320_);
  or (_02337_, _02216_, _33753_);
  or (_02338_, _02220_, _33700_);
  and (_02339_, _02338_, _02337_);
  or (_02340_, _02225_, _33575_);
  or (_02341_, _02227_, _33534_);
  and (_02342_, _02341_, _02340_);
  and (_02343_, _02342_, _02339_);
  nand (_02344_, _02233_, _33979_);
  or (_02345_, _02236_, _33923_);
  and (_02346_, _02345_, _02344_);
  or (_02347_, _02240_, _33409_);
  or (_02348_, _02242_, _33368_);
  and (_02349_, _02348_, _02347_);
  and (_02350_, _02349_, _02346_);
  and (_02351_, _02350_, _02343_);
  or (_02352_, _02249_, _33865_);
  or (_02353_, _02252_, _33809_);
  and (_02354_, _02353_, _02352_);
  or (_02355_, _02255_, _33258_);
  or (_02356_, _02257_, _33299_);
  and (_02357_, _02356_, _02355_);
  and (_02358_, _02357_, _02354_);
  or (_02359_, _02261_, _33657_);
  or (_02360_, _02263_, _33616_);
  and (_02361_, _02360_, _02359_);
  or (_02362_, _02266_, _33493_);
  or (_02363_, _02268_, _33452_);
  and (_02364_, _02363_, _02362_);
  and (_02365_, _02364_, _02361_);
  and (_02366_, _02365_, _02358_);
  nand (_02367_, _02366_, _02351_);
  or (_02368_, _02367_, _02336_);
  not (_02369_, _02368_);
  and (_02370_, _02369_, _02305_);
  or (_02371_, _02216_, _33732_);
  or (_02372_, _02220_, _33683_);
  and (_02373_, _02372_, _02371_);
  or (_02374_, _02225_, _33560_);
  or (_02375_, _02227_, _33519_);
  and (_02376_, _02375_, _02374_);
  and (_02377_, _02376_, _02373_);
  nand (_02378_, _02233_, _33958_);
  or (_02379_, _02236_, _33902_);
  and (_02380_, _02379_, _02378_);
  or (_02381_, _02240_, _33394_);
  or (_02382_, _02242_, _33338_);
  and (_02383_, _02382_, _02381_);
  and (_02384_, _02383_, _02380_);
  and (_02385_, _02384_, _02377_);
  or (_02386_, _02249_, _33844_);
  or (_02387_, _02252_, _33789_);
  and (_02388_, _02387_, _02386_);
  or (_02389_, _02255_, _33243_);
  or (_02390_, _02257_, _33284_);
  and (_02391_, _02390_, _02389_);
  and (_02392_, _02391_, _02388_);
  or (_02393_, _02261_, _33642_);
  or (_02394_, _02263_, _33601_);
  and (_02395_, _02394_, _02393_);
  or (_02396_, _02266_, _33478_);
  or (_02397_, _02268_, _33435_);
  and (_02398_, _02397_, _02396_);
  and (_02399_, _02398_, _02395_);
  and (_02400_, _02399_, _02392_);
  nand (_02401_, _02400_, _02385_);
  or (_02402_, _02216_, _33739_);
  or (_02403_, _02220_, _33688_);
  and (_02404_, _02403_, _02402_);
  or (_02405_, _02225_, _33565_);
  or (_02406_, _02227_, _33524_);
  and (_02407_, _02406_, _02405_);
  and (_02408_, _02407_, _02404_);
  nand (_02409_, _02233_, _33965_);
  or (_02410_, _02236_, _33909_);
  and (_02411_, _02410_, _02409_);
  or (_02412_, _02240_, _33399_);
  or (_02413_, _02242_, _33349_);
  and (_02414_, _02413_, _02412_);
  and (_02415_, _02414_, _02411_);
  and (_02416_, _02415_, _02408_);
  or (_02417_, _02249_, _33851_);
  or (_02418_, _02252_, _33795_);
  and (_02419_, _02418_, _02417_);
  or (_02420_, _02255_, _33248_);
  or (_02421_, _02257_, _33289_);
  and (_02422_, _02421_, _02420_);
  and (_02423_, _02422_, _02419_);
  or (_02424_, _02261_, _33647_);
  or (_02425_, _02263_, _33606_);
  and (_02426_, _02425_, _02424_);
  or (_02427_, _02266_, _33483_);
  or (_02428_, _02268_, _33441_);
  and (_02429_, _02428_, _02427_);
  and (_02430_, _02429_, _02426_);
  and (_02431_, _02430_, _02423_);
  nand (_02432_, _02431_, _02416_);
  or (_02433_, _02432_, _02401_);
  not (_02434_, _02433_);
  or (_02435_, _02216_, _33720_);
  or (_02436_, _02220_, _33673_);
  and (_02437_, _02436_, _02435_);
  or (_02438_, _02225_, _33550_);
  or (_02439_, _02227_, _33509_);
  and (_02440_, _02439_, _02438_);
  and (_02441_, _02440_, _02437_);
  nand (_02442_, _02233_, _33944_);
  or (_02443_, _02236_, _33888_);
  and (_02444_, _02443_, _02442_);
  or (_02445_, _02240_, _33384_);
  or (_02446_, _02242_, _33316_);
  and (_02447_, _02446_, _02445_);
  and (_02448_, _02447_, _02444_);
  and (_02449_, _02448_, _02441_);
  or (_02450_, _02249_, _33830_);
  or (_02451_, _02252_, _33774_);
  and (_02452_, _02451_, _02450_);
  or (_02453_, _02255_, _33233_);
  or (_02454_, _02257_, _33274_);
  and (_02455_, _02454_, _02453_);
  and (_02456_, _02455_, _02452_);
  or (_02457_, _02261_, _33632_);
  or (_02458_, _02263_, _33591_);
  and (_02459_, _02458_, _02457_);
  or (_02460_, _02266_, _33468_);
  or (_02461_, _02268_, _33425_);
  and (_02462_, _02461_, _02460_);
  and (_02463_, _02462_, _02459_);
  and (_02464_, _02463_, _02456_);
  and (_02465_, _02464_, _02449_);
  or (_02466_, _02216_, _33726_);
  or (_02467_, _02220_, _33678_);
  and (_02468_, _02467_, _02466_);
  or (_02469_, _02225_, _33555_);
  or (_02470_, _02227_, _33514_);
  and (_02471_, _02470_, _02469_);
  and (_02472_, _02471_, _02468_);
  nand (_02473_, _02233_, _33951_);
  or (_02474_, _02236_, _33895_);
  and (_02475_, _02474_, _02473_);
  or (_02476_, _02240_, _33389_);
  or (_02477_, _02242_, _33327_);
  and (_02478_, _02477_, _02476_);
  and (_02479_, _02478_, _02475_);
  and (_02480_, _02479_, _02472_);
  or (_02481_, _02249_, _33837_);
  or (_02482_, _02252_, _33781_);
  and (_02483_, _02482_, _02481_);
  or (_02484_, _02255_, _33238_);
  or (_02485_, _02257_, _33279_);
  and (_02486_, _02485_, _02484_);
  and (_02487_, _02486_, _02483_);
  or (_02488_, _02261_, _33637_);
  or (_02489_, _02263_, _33596_);
  and (_02490_, _02489_, _02488_);
  or (_02491_, _02266_, _33473_);
  or (_02492_, _02268_, _33430_);
  and (_02493_, _02492_, _02491_);
  and (_02494_, _02493_, _02490_);
  and (_02495_, _02494_, _02487_);
  nand (_02496_, _02495_, _02480_);
  not (_02497_, _02496_);
  and (_02498_, _02497_, _02465_);
  and (_02499_, _02498_, _02434_);
  and (_02500_, _02499_, _02370_);
  not (_02501_, _02500_);
  or (_02502_, _02496_, _02465_);
  or (_02503_, _02502_, _02433_);
  not (_02504_, _02503_);
  nand (_02505_, _02335_, _02320_);
  and (_02506_, _02366_, _02351_);
  or (_02507_, _02506_, _02505_);
  not (_02508_, _02507_);
  nand (_02509_, _02272_, _02246_);
  and (_02510_, _02304_, _02509_);
  and (_02511_, _02510_, _02508_);
  and (_02512_, _02511_, _02504_);
  not (_02513_, _02512_);
  or (_02514_, _02506_, _02336_);
  not (_02515_, _02514_);
  and (_02516_, _02515_, _02510_);
  and (_02517_, _02516_, _02504_);
  or (_02518_, _02367_, _02505_);
  or (_02519_, _02304_, _02509_);
  nor (_02520_, _02519_, _02518_);
  and (_02521_, _02520_, _02504_);
  nor (_02522_, _02521_, _02517_);
  and (_02523_, _02522_, _02513_);
  not (_02524_, _02518_);
  and (_02525_, _02524_, _02305_);
  and (_02526_, _02525_, _02504_);
  not (_02527_, _02526_);
  and (_02528_, _02504_, _02370_);
  not (_02529_, _02528_);
  and (_02530_, _02515_, _02305_);
  and (_02531_, _02530_, _02504_);
  and (_02532_, _02510_, _02369_);
  and (_02533_, _02532_, _02504_);
  nor (_02534_, _02533_, _02531_);
  and (_02535_, _02508_, _02305_);
  and (_02536_, _02535_, _02504_);
  and (_02537_, _02524_, _02510_);
  and (_02538_, _02537_, _02504_);
  nor (_02539_, _02538_, _02536_);
  and (_02540_, _02539_, _02534_);
  and (_02541_, _02540_, _02529_);
  and (_02542_, _02541_, _02527_);
  and (_02543_, _02542_, _02523_);
  or (_02544_, _02543_, \oc8051_golden_model_1.PC [0]);
  not (_02545_, _02465_);
  and (_02546_, _02496_, _02545_);
  and (_02547_, _02546_, _02434_);
  and (_02548_, _02547_, _02520_);
  not (_02549_, \oc8051_golden_model_1.ACC [0]);
  and (_02550_, _02549_, \oc8051_golden_model_1.PC [0]);
  and (_02551_, \oc8051_golden_model_1.ACC [0], _02247_);
  nor (_02552_, _02551_, _02550_);
  and (_02553_, _02552_, _02548_);
  or (_02554_, _02304_, _02273_);
  or (_02555_, _02554_, _02368_);
  or (_02556_, _02555_, _02503_);
  or (_02557_, _02554_, _02514_);
  or (_02558_, _02557_, _02503_);
  and (_02559_, _02558_, _02556_);
  or (_02560_, _02519_, _02514_);
  or (_02561_, _02560_, _02503_);
  or (_02562_, _02554_, _02507_);
  or (_02563_, _02562_, _02503_);
  and (_02564_, _02563_, _02561_);
  or (_02565_, _02519_, _02507_);
  or (_02566_, _02565_, _02503_);
  or (_02567_, _02554_, _02518_);
  or (_02568_, _02567_, _02503_);
  and (_02569_, _02568_, _02566_);
  and (_02570_, _02569_, _02564_);
  nand (_02571_, _02570_, _02559_);
  not (_02572_, _02502_);
  not (_02573_, _02401_);
  nor (_02574_, _02432_, _02573_);
  and (_02575_, _02574_, _02572_);
  and (_02576_, _02575_, _02520_);
  nor (_02577_, _02519_, _02368_);
  and (_02578_, _02577_, _02504_);
  nor (_02579_, _02578_, _02576_);
  not (_02580_, _02579_);
  or (_02581_, _02580_, _02571_);
  nand (_02582_, _02581_, _02247_);
  not (_02583_, _02543_);
  not (_02584_, _02548_);
  and (_02585_, _02577_, _02547_);
  not (_02586_, _02585_);
  or (_02587_, _02571_, _02247_);
  and (_02588_, _02587_, _02586_);
  and (_02589_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02590_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02591_, _02590_, _02589_);
  nand (_02592_, _02591_, _02585_);
  nand (_02593_, _02592_, _02579_);
  or (_02594_, _02593_, _02588_);
  and (_02595_, _02594_, _02584_);
  or (_02596_, _02595_, _02583_);
  and (_02597_, _02596_, _02582_);
  or (_02598_, _02597_, _02553_);
  nand (_02599_, _02598_, _02544_);
  and (_02600_, _02570_, _02559_);
  or (_02601_, _02600_, \oc8051_golden_model_1.PC [1]);
  and (_02602_, _02248_, _02219_);
  or (_02603_, _02602_, _02571_);
  nand (_02604_, _02603_, _02601_);
  nand (_02605_, _02604_, _02586_);
  and (_02606_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02607_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02608_, _02607_, _02606_);
  and (_02609_, _02608_, _02589_);
  nor (_02610_, _02608_, _02589_);
  nor (_02611_, _02610_, _02609_);
  nand (_02612_, _02611_, _02585_);
  and (_02613_, _02612_, _02579_);
  nand (_02614_, _02613_, _02605_);
  or (_02615_, _02579_, _02218_);
  and (_02616_, _02615_, _02584_);
  and (_02617_, _02616_, _02614_);
  not (_02618_, \oc8051_golden_model_1.ACC [1]);
  nor (_02619_, _02602_, _02618_);
  and (_02620_, _02602_, _02618_);
  nor (_02621_, _02620_, _02619_);
  and (_02622_, _02621_, _02551_);
  nor (_02623_, _02621_, _02551_);
  nor (_02624_, _02623_, _02622_);
  and (_02625_, _02624_, _02548_);
  or (_02626_, _02625_, _02617_);
  and (_02627_, _02626_, _02543_);
  nor (_02628_, _02543_, \oc8051_golden_model_1.PC [1]);
  or (_02629_, _02628_, _02627_);
  and (_02630_, _02629_, _02599_);
  and (_02631_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02632_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02633_, _02632_, _02631_);
  not (_02634_, _02633_);
  and (_02635_, _02634_, _02581_);
  and (_02636_, _02231_, \oc8051_golden_model_1.PC [2]);
  and (_02637_, _02213_, _02223_);
  nor (_02638_, _02637_, _02636_);
  nor (_02639_, _02638_, _02585_);
  and (_02640_, _02639_, _02600_);
  nor (_02641_, _02609_, _02606_);
  and (_02642_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02643_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02644_, _02643_, _02642_);
  not (_02645_, _02644_);
  nor (_02646_, _02645_, _02641_);
  and (_02647_, _02645_, _02641_);
  nor (_02648_, _02647_, _02646_);
  not (_02649_, _02648_);
  and (_02650_, _02649_, _02585_);
  or (_02651_, _02650_, _02640_);
  and (_02652_, _02651_, _02579_);
  or (_02653_, _02652_, _02548_);
  or (_02654_, _02653_, _02635_);
  nor (_02655_, _02622_, _02619_);
  and (_02656_, _02638_, \oc8051_golden_model_1.ACC [2]);
  nor (_02657_, _02638_, \oc8051_golden_model_1.ACC [2]);
  nor (_02658_, _02657_, _02656_);
  not (_02659_, _02658_);
  and (_02660_, _02659_, _02655_);
  nor (_02661_, _02659_, _02655_);
  nor (_02662_, _02661_, _02660_);
  and (_02663_, _02662_, _02548_);
  not (_02664_, _02663_);
  and (_02665_, _02664_, _02523_);
  nand (_02666_, _02665_, _02654_);
  not (_02667_, _02542_);
  nor (_02668_, _02633_, _02523_);
  nor (_02669_, _02668_, _02667_);
  nand (_02670_, _02669_, _02666_);
  nor (_02671_, _02634_, _02542_);
  not (_02672_, _02671_);
  and (_02673_, _02672_, _02670_);
  and (_02674_, _02232_, \oc8051_golden_model_1.PC [1]);
  nor (_02675_, _02631_, \oc8051_golden_model_1.PC [3]);
  nor (_02676_, _02675_, _02674_);
  not (_02677_, _02676_);
  or (_02678_, _02581_, _02583_);
  and (_02679_, _02678_, _02677_);
  nor (_02680_, _02646_, _02642_);
  and (_02681_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02682_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02683_, _02682_, _02681_);
  not (_02684_, _02683_);
  nor (_02685_, _02684_, _02680_);
  and (_02686_, _02684_, _02680_);
  nor (_02687_, _02686_, _02685_);
  not (_02688_, _02687_);
  and (_02689_, _02688_, _02585_);
  not (_02690_, _02225_);
  nor (_02691_, _02636_, _02214_);
  nor (_02692_, _02691_, _02690_);
  not (_02693_, _02692_);
  nor (_02694_, _02585_, _02693_);
  and (_02695_, _02694_, _02600_);
  or (_02696_, _02695_, _02689_);
  and (_02697_, _02579_, _02584_);
  and (_02698_, _02697_, _02696_);
  nor (_02700_, _02661_, _02656_);
  not (_02701_, \oc8051_golden_model_1.ACC [3]);
  nor (_02702_, _02692_, _02701_);
  and (_02703_, _02692_, _02701_);
  nor (_02704_, _02703_, _02702_);
  or (_02705_, _02704_, _02700_);
  nand (_02706_, _02704_, _02700_);
  and (_02707_, _02706_, _02705_);
  and (_02708_, _02707_, _02548_);
  or (_02709_, _02708_, _02698_);
  and (_02710_, _02709_, _02543_);
  or (_02711_, _02710_, _02679_);
  nor (_02712_, _02711_, _02673_);
  and (_02713_, _02712_, _02630_);
  nand (_02714_, _02713_, _01164_);
  and (_02715_, _02598_, _02544_);
  nor (_02716_, _02628_, _02627_);
  and (_02717_, _02716_, _02715_);
  and (_02718_, _02717_, _02712_);
  nand (_02719_, _02718_, _01167_);
  and (_02720_, _02719_, _02714_);
  and (_02721_, _02716_, _02599_);
  nand (_02722_, _02672_, _02670_);
  and (_02723_, _02711_, _02722_);
  and (_02724_, _02723_, _02721_);
  nand (_02725_, _02724_, _01134_);
  and (_02726_, _02629_, _02715_);
  and (_02727_, _02711_, _02673_);
  and (_02728_, _02727_, _02726_);
  nand (_02729_, _02728_, _01147_);
  and (_02730_, _02729_, _02725_);
  and (_02731_, _02730_, _02720_);
  and (_02732_, _02723_, _02630_);
  nand (_02733_, _02732_, _01129_);
  and (_02734_, _02723_, _02717_);
  nand (_02735_, _02734_, _01125_);
  and (_02736_, _02735_, _02733_);
  and (_02737_, _02727_, _02630_);
  nand (_02738_, _02737_, _01157_);
  and (_02739_, _02727_, _02717_);
  nand (_02740_, _02739_, _01085_);
  and (_02741_, _02740_, _02738_);
  and (_02742_, _02741_, _02736_);
  and (_02743_, _02742_, _02731_);
  nor (_02744_, _02711_, _02722_);
  and (_02745_, _02744_, _02630_);
  nand (_02746_, _02745_, _01161_);
  and (_02747_, _02744_, _02721_);
  nand (_02748_, _02747_, _01119_);
  and (_02749_, _02748_, _02746_);
  and (_02750_, _02726_, _02712_);
  nand (_02751_, _02750_, _33937_);
  and (_02752_, _02721_, _02712_);
  nand (_02753_, _02752_, _01170_);
  and (_02754_, _02753_, _02751_);
  and (_02755_, _02754_, _02749_);
  and (_02756_, _02726_, _02723_);
  nand (_02757_, _02756_, _01140_);
  and (_02758_, _02727_, _02721_);
  nand (_02759_, _02758_, _01154_);
  and (_02760_, _02759_, _02757_);
  and (_02761_, _02744_, _02726_);
  nand (_02762_, _02761_, _01137_);
  and (_02763_, _02744_, _02717_);
  nand (_02764_, _02763_, _01115_);
  and (_02765_, _02764_, _02762_);
  and (_02766_, _02765_, _02760_);
  and (_02767_, _02766_, _02755_);
  nand (_02768_, _02767_, _02743_);
  nand (_02769_, _02752_, _01430_);
  nand (_02770_, _02758_, _01441_);
  and (_02771_, _02770_, _02769_);
  nand (_02772_, _02718_, _01432_);
  nand (_02773_, _02756_, _01413_);
  and (_02774_, _02773_, _02772_);
  and (_02775_, _02774_, _02771_);
  nand (_02776_, _02713_, _01434_);
  nand (_02777_, _02745_, _01405_);
  and (_02778_, _02777_, _02776_);
  nand (_02779_, _02728_, _01415_);
  nand (_02780_, _02739_, _01443_);
  and (_02781_, _02780_, _02779_);
  and (_02782_, _02781_, _02778_);
  and (_02783_, _02782_, _02775_);
  nand (_02784_, _02763_, _01403_);
  nand (_02785_, _02724_, _01426_);
  and (_02786_, _02785_, _02784_);
  nand (_02787_, _02750_, _33965_);
  nand (_02788_, _02761_, _01419_);
  and (_02789_, _02788_, _02787_);
  and (_02790_, _02789_, _02786_);
  nand (_02791_, _02747_, _01407_);
  nand (_02792_, _02732_, _01411_);
  and (_02793_, _02792_, _02791_);
  nand (_02794_, _02734_, _01424_);
  nand (_02795_, _02737_, _01438_);
  and (_02796_, _02795_, _02794_);
  and (_02797_, _02796_, _02793_);
  and (_02798_, _02797_, _02790_);
  and (_02799_, _02798_, _02783_);
  or (_02800_, _02799_, _02768_);
  nor (_02801_, _02800_, _02501_);
  nand (_02802_, _02761_, _01283_);
  nand (_02803_, _02745_, _01270_);
  and (_02804_, _02803_, _02802_);
  nand (_02805_, _02756_, _01285_);
  nand (_02806_, _02732_, _01278_);
  and (_02807_, _02806_, _02805_);
  and (_02808_, _02807_, _02804_);
  nand (_02809_, _02750_, _33944_);
  nand (_02810_, _02713_, _01304_);
  and (_02811_, _02810_, _02809_);
  nand (_02812_, _02728_, _01289_);
  nand (_02813_, _02737_, _01297_);
  and (_02814_, _02813_, _02812_);
  and (_02815_, _02814_, _02811_);
  and (_02816_, _02815_, _02808_);
  nand (_02817_, _02718_, _01302_);
  nand (_02818_, _02752_, _01306_);
  and (_02819_, _02818_, _02817_);
  nand (_02820_, _02758_, _01295_);
  nand (_02821_, _02739_, _01268_);
  and (_02822_, _02821_, _02820_);
  and (_02823_, _02822_, _02819_);
  nand (_02824_, _02763_, _01272_);
  nand (_02825_, _02747_, _01300_);
  and (_02826_, _02825_, _02824_);
  nand (_02827_, _02734_, _01276_);
  nand (_02828_, _02724_, _01281_);
  and (_02829_, _02828_, _02827_);
  and (_02830_, _02829_, _02826_);
  and (_02831_, _02830_, _02823_);
  and (_02832_, _02831_, _02816_);
  not (_02833_, _02832_);
  and (_02834_, _02432_, _02401_);
  and (_02835_, _02834_, _02572_);
  and (_02836_, _02835_, _02520_);
  and (_02837_, _02834_, _02496_);
  and (_02838_, _02837_, _02520_);
  nor (_02839_, _02838_, _02836_);
  nor (_02840_, _02839_, _02768_);
  and (_02841_, _02496_, _02465_);
  and (_02842_, _02432_, _02573_);
  and (_02843_, _02842_, _02841_);
  and (_02844_, _02843_, _02520_);
  and (_02845_, _02842_, _02546_);
  and (_02846_, _02845_, _02520_);
  nor (_02847_, _02846_, _02844_);
  nor (_02848_, _02847_, _02768_);
  or (_02849_, _02848_, _02840_);
  not (_02850_, _02849_);
  not (_02851_, _02576_);
  nor (_02852_, _02768_, _02851_);
  not (_02853_, _02852_);
  and (_02854_, _02574_, _02496_);
  and (_02855_, _02854_, _02520_);
  not (_02856_, _02855_);
  nor (_02857_, _02856_, _02768_);
  not (_02858_, _02768_);
  and (_02859_, _02834_, _02498_);
  and (_02860_, _02859_, _02520_);
  not (_02861_, _02860_);
  and (_02862_, _02842_, _02498_);
  and (_02863_, _02862_, _02520_);
  and (_02864_, _02842_, _02572_);
  and (_02865_, _02864_, _02520_);
  nor (_02866_, _02865_, _02863_);
  nand (_02867_, _02866_, _02861_);
  and (_02868_, _02867_, _02858_);
  nor (_02869_, _02868_, _02857_);
  and (_02870_, _02869_, _02853_);
  and (_02871_, _02870_, _02850_);
  nor (_02872_, _02871_, _02833_);
  and (_02873_, _02841_, _02434_);
  and (_02874_, _02873_, _02577_);
  not (_02875_, _02874_);
  nor (_02876_, _02875_, _02800_);
  not (_02877_, \oc8051_golden_model_1.SP [0]);
  nor (_02878_, _02561_, _02877_);
  not (_02879_, _02560_);
  and (_02880_, _02873_, _02879_);
  not (_02881_, _02880_);
  nor (_02882_, _02881_, _02800_);
  nor (_02883_, _02881_, _02768_);
  not (_02884_, _02883_);
  not (_02885_, _02567_);
  and (_02886_, _02885_, _02499_);
  and (_02887_, _02873_, _02885_);
  not (_02888_, _02887_);
  nor (_02889_, _02888_, _02800_);
  not (_02890_, _02555_);
  and (_02891_, _02873_, _02890_);
  not (_02892_, _02891_);
  or (_02893_, _02892_, _02800_);
  nor (_02894_, _02892_, _02768_);
  and (_02895_, _02535_, _02499_);
  not (_02896_, _02895_);
  and (_02897_, _02873_, _02535_);
  not (_02898_, _02897_);
  and (_02899_, _02575_, _02535_);
  not (_02901_, _02899_);
  and (_02902_, _02750_, _33986_);
  and (_02903_, _02761_, _01554_);
  nor (_02904_, _02903_, _02902_);
  and (_02905_, _02724_, _01561_);
  and (_02906_, _02758_, _01576_);
  nor (_02907_, _02906_, _02905_);
  and (_02908_, _02907_, _02904_);
  and (_02909_, _02713_, _01567_);
  and (_02910_, _02718_, _01569_);
  nor (_02911_, _02910_, _02909_);
  and (_02912_, _02745_, _01542_);
  and (_02913_, _02763_, _01565_);
  nor (_02914_, _02913_, _02912_);
  and (_02915_, _02914_, _02911_);
  and (_02916_, _02915_, _02908_);
  and (_02917_, _02756_, _01550_);
  and (_02918_, _02732_, _01546_);
  nor (_02919_, _02918_, _02917_);
  and (_02920_, _02734_, _01559_);
  and (_02921_, _02728_, _01548_);
  nor (_02922_, _02921_, _02920_);
  and (_02923_, _02922_, _02919_);
  and (_02924_, _02737_, _01540_);
  and (_02925_, _02739_, _01578_);
  nor (_02926_, _02925_, _02924_);
  and (_02927_, _02752_, _01571_);
  and (_02928_, _02747_, _01538_);
  nor (_02929_, _02928_, _02927_);
  and (_02930_, _02929_, _02926_);
  and (_02931_, _02930_, _02923_);
  and (_02932_, _02931_, _02916_);
  nor (_02933_, _02932_, _02768_);
  not (_02934_, _02799_);
  and (_02935_, _02934_, _02768_);
  nor (_02936_, _02935_, _02933_);
  and (_02937_, _02873_, _02516_);
  and (_02938_, _02873_, _02520_);
  nor (_02939_, _02938_, _02937_);
  not (_02940_, _02939_);
  and (_02941_, _02940_, _02936_);
  and (_02942_, _02879_, _02499_);
  nor (_02943_, _02880_, _02942_);
  or (_02944_, _02943_, _02936_);
  and (_02945_, _02936_, _02891_);
  not (_02946_, \oc8051_golden_model_1.SP [3]);
  and (_02947_, _02890_, _02499_);
  and (_02948_, _02947_, _02946_);
  or (_02949_, _02948_, _02945_);
  and (_02950_, _02575_, _02885_);
  nor (_02951_, _02947_, _02891_);
  and (_02952_, _02575_, _02890_);
  not (_02953_, _02562_);
  and (_02954_, _02575_, _02953_);
  nor (_02955_, _02954_, _02952_);
  nand (_02956_, _02955_, \oc8051_golden_model_1.PSW [3]);
  and (_02957_, _02956_, _02951_);
  or (_02958_, _02957_, _02950_);
  not (_02959_, _02950_);
  nand (_02960_, _02955_, _02959_);
  nand (_02961_, _02960_, _02934_);
  and (_02962_, _02961_, _02958_);
  or (_02963_, _02962_, _02887_);
  or (_02964_, _02963_, _02949_);
  or (_02965_, _02936_, _02888_);
  and (_02966_, _02575_, _02879_);
  nor (_02967_, _02966_, _02886_);
  and (_02968_, _02967_, _02965_);
  and (_02969_, _02968_, _02964_);
  not (_02970_, _02943_);
  nor (_02971_, _02967_, _02934_);
  or (_02972_, _02971_, _02970_);
  or (_02973_, _02972_, _02969_);
  and (_02974_, _02973_, _02944_);
  nor (_02975_, _02837_, _02835_);
  nor (_02976_, _02859_, _02845_);
  and (_02977_, _02976_, _02975_);
  nor (_02978_, _02977_, _02565_);
  not (_02979_, _02546_);
  not (_02980_, _02565_);
  and (_02981_, _02842_, _02980_);
  and (_02982_, _02981_, _02979_);
  nor (_02983_, _02982_, _02978_);
  not (_02984_, _02983_);
  or (_02985_, _02984_, _02974_);
  and (_02986_, _02980_, _02499_);
  and (_02987_, _02873_, _02980_);
  nor (_02988_, _02987_, _02986_);
  or (_02989_, _02983_, _02799_);
  and (_02990_, _02989_, _02988_);
  and (_02991_, _02990_, _02985_);
  and (_02992_, _02577_, _02575_);
  not (_02993_, _02988_);
  and (_02994_, _02993_, _02936_);
  or (_02995_, _02994_, _02992_);
  or (_02996_, _02995_, _02991_);
  not (_02997_, _02992_);
  or (_02998_, _02997_, _02799_);
  and (_02999_, _02998_, _02875_);
  and (_03000_, _02999_, _02996_);
  and (_03001_, _02936_, _02874_);
  or (_03002_, _03001_, _02576_);
  or (_03003_, _03002_, _03000_);
  and (_03004_, _02873_, _02370_);
  nor (_03005_, _03004_, _02895_);
  and (_03006_, _02873_, _02525_);
  nor (_03007_, _03006_, _02500_);
  and (_03008_, _03007_, _03005_);
  and (_03009_, _02864_, _02879_);
  and (_03010_, _02842_, _02496_);
  nor (_03011_, _02859_, _03010_);
  nor (_03012_, _03011_, _02560_);
  nor (_03013_, _03012_, _03009_);
  and (_03014_, _02575_, _02516_);
  nor (_03015_, _03014_, _02966_);
  and (_03016_, _03015_, _03013_);
  and (_03017_, _02834_, _02841_);
  and (_03018_, _03017_, _02879_);
  not (_03019_, _03018_);
  and (_03020_, _02547_, _02532_);
  and (_03021_, _02547_, _02511_);
  nor (_03022_, _03021_, _03020_);
  and (_03023_, _02577_, _02499_);
  and (_03024_, _02574_, _02498_);
  and (_03025_, _03024_, _02879_);
  nor (_03026_, _03025_, _03023_);
  and (_03027_, _03026_, _03022_);
  and (_03028_, _03027_, _03019_);
  and (_03029_, _02834_, _02546_);
  nor (_03030_, _03029_, _02835_);
  not (_03031_, _02862_);
  and (_03032_, _03031_, _03030_);
  nor (_03033_, _03032_, _02560_);
  not (_03034_, _03033_);
  and (_03035_, _02530_, _02499_);
  and (_03036_, _02547_, _02537_);
  nor (_03037_, _03036_, _03035_);
  and (_03038_, _02854_, _02879_);
  nor (_03039_, _03038_, _02952_);
  and (_03040_, _03039_, _03037_);
  and (_03041_, _03040_, _03034_);
  and (_03042_, _03041_, _03028_);
  and (_03043_, _03042_, _03016_);
  and (_03044_, _03043_, _03008_);
  nor (_03045_, _03044_, _02247_);
  and (_03046_, _03044_, _02247_);
  nor (_03047_, _03046_, _03045_);
  not (_03048_, _03047_);
  nor (_03049_, _03046_, _02218_);
  and (_03050_, _03046_, _02218_);
  nor (_03051_, _03050_, _03049_);
  and (_03052_, _03051_, _03048_);
  nor (_03053_, _03044_, _02633_);
  not (_03054_, _02638_);
  and (_03055_, _03008_, _03054_);
  and (_03056_, _03055_, _03043_);
  nor (_03057_, _03056_, _03053_);
  nor (_03058_, _03044_, _02677_);
  and (_03059_, _03044_, _02693_);
  nor (_03060_, _03059_, _03058_);
  and (_03062_, _03060_, _03057_);
  and (_03063_, _03062_, _03052_);
  and (_03064_, _03063_, _01413_);
  nor (_03065_, _03051_, _03048_);
  not (_03066_, _03060_);
  nor (_03067_, _03066_, _03057_);
  and (_03068_, _03067_, _03065_);
  and (_03069_, _03068_, _01441_);
  nor (_03070_, _03069_, _03064_);
  and (_03071_, _03066_, _03057_);
  and (_03073_, _03051_, _03047_);
  and (_03074_, _03073_, _03071_);
  and (_03075_, _03074_, _01434_);
  and (_03076_, _03067_, _03052_);
  and (_03077_, _03076_, _01415_);
  nor (_03078_, _03077_, _03075_);
  and (_03079_, _03078_, _03070_);
  nor (_03080_, _03051_, _03047_);
  and (_03081_, _03080_, _03071_);
  and (_03082_, _03081_, _01432_);
  and (_03083_, _03071_, _03065_);
  and (_03084_, _03083_, _01430_);
  nor (_03085_, _03084_, _03082_);
  and (_03086_, _03080_, _03062_);
  and (_03087_, _03086_, _01424_);
  and (_03088_, _03065_, _03062_);
  and (_03089_, _03088_, _01426_);
  nor (_03090_, _03089_, _03087_);
  and (_03091_, _03090_, _03085_);
  and (_03092_, _03091_, _03079_);
  and (_03094_, _03073_, _03067_);
  and (_03095_, _03094_, _01438_);
  and (_03096_, _03080_, _03067_);
  and (_03097_, _03096_, _01443_);
  nor (_03098_, _03097_, _03095_);
  nor (_03099_, _03060_, _03057_);
  and (_03100_, _03099_, _03073_);
  and (_03101_, _03100_, _01405_);
  and (_03102_, _03099_, _03065_);
  and (_03103_, _03102_, _01407_);
  nor (_03105_, _03103_, _03101_);
  and (_03106_, _03105_, _03098_);
  and (_03107_, _03071_, _03052_);
  and (_03108_, _03107_, _33965_);
  and (_03109_, _03073_, _03062_);
  and (_03110_, _03109_, _01411_);
  nor (_03111_, _03110_, _03108_);
  and (_03112_, _03099_, _03052_);
  and (_03113_, _03112_, _01419_);
  and (_03114_, _03099_, _03080_);
  and (_03116_, _03114_, _01403_);
  nor (_03117_, _03116_, _03113_);
  and (_03118_, _03117_, _03111_);
  and (_03119_, _03118_, _03106_);
  and (_03120_, _03119_, _03092_);
  or (_03121_, _03120_, _02851_);
  and (_03122_, _03121_, _02939_);
  and (_03123_, _03122_, _03003_);
  or (_03124_, _03123_, _02941_);
  and (_03125_, _02575_, _02537_);
  not (_03126_, _03125_);
  and (_03127_, _02873_, _02537_);
  nor (_03128_, _03127_, _03036_);
  and (_03129_, _03128_, _03126_);
  and (_03130_, _02873_, _02511_);
  not (_03131_, _03130_);
  and (_03132_, _02575_, _02511_);
  nor (_03133_, _03132_, _03021_);
  and (_03134_, _03133_, _03131_);
  and (_03135_, _03134_, _03129_);
  and (_03137_, _02575_, _02530_);
  not (_03138_, _03137_);
  and (_03139_, _02873_, _02532_);
  not (_03140_, _03139_);
  and (_03141_, _02575_, _02532_);
  nor (_03142_, _03141_, _03020_);
  and (_03143_, _03142_, _03140_);
  and (_03144_, _03143_, _03138_);
  and (_03145_, _03144_, _03135_);
  and (_03146_, _03145_, _03124_);
  and (_03148_, _02873_, _02530_);
  nor (_03149_, _03145_, _02934_);
  or (_03150_, _03149_, _03148_);
  or (_03151_, _03150_, _03146_);
  not (_03152_, _03035_);
  nand (_03153_, _03148_, \oc8051_golden_model_1.SP [3]);
  and (_03154_, _03153_, _03152_);
  and (_03155_, _03154_, _03151_);
  and (_03156_, _03035_, _02936_);
  or (_03157_, _03156_, _03155_);
  and (_03159_, _03157_, _02901_);
  and (_03160_, _02899_, _02799_);
  nor (_03161_, _03160_, _03159_);
  and (_03162_, _03161_, _02898_);
  and (_03163_, _02897_, \oc8051_golden_model_1.SP [3]);
  or (_03164_, _03163_, _03162_);
  and (_03165_, _03164_, _02896_);
  and (_03166_, _02575_, _02370_);
  nor (_03167_, _02936_, _02896_);
  or (_03168_, _03167_, _03166_);
  or (_03170_, _03168_, _03165_);
  nand (_03171_, _03166_, _02799_);
  and (_03172_, _03171_, _03170_);
  nor (_03173_, _03172_, _02500_);
  and (_03174_, _02575_, _02525_);
  and (_03175_, _02936_, _02500_);
  or (_03176_, _03175_, _03174_);
  nor (_03177_, _03176_, _03173_);
  not (_03178_, _03174_);
  nor (_03179_, _03178_, _02799_);
  nor (_03181_, _03179_, _03177_);
  and (_03182_, _02756_, _01509_);
  and (_03183_, _02728_, _01523_);
  nor (_03184_, _03183_, _03182_);
  and (_03185_, _02713_, _01503_);
  and (_03186_, _02747_, _01493_);
  nor (_03187_, _03186_, _03185_);
  and (_03188_, _03187_, _03184_);
  and (_03189_, _02737_, _01531_);
  and (_03190_, _02739_, _01516_);
  nor (_03192_, _03190_, _03189_);
  and (_03193_, _02732_, _01518_);
  and (_03194_, _02724_, _01525_);
  nor (_03195_, _03194_, _03193_);
  and (_03196_, _03195_, _03192_);
  and (_03197_, _03196_, _03188_);
  and (_03198_, _02752_, _01511_);
  and (_03199_, _02761_, _01501_);
  nor (_03200_, _03199_, _03198_);
  and (_03201_, _02750_, _33979_);
  and (_03203_, _02718_, _01505_);
  nor (_03204_, _03203_, _03201_);
  and (_03205_, _03204_, _03200_);
  and (_03206_, _02745_, _01497_);
  and (_03207_, _02763_, _01495_);
  nor (_03208_, _03207_, _03206_);
  and (_03209_, _02734_, _01520_);
  and (_03210_, _02758_, _01533_);
  nor (_03211_, _03210_, _03209_);
  and (_03212_, _03211_, _03208_);
  and (_03214_, _03212_, _03205_);
  and (_03215_, _03214_, _03197_);
  nor (_03216_, _03215_, _02768_);
  and (_03217_, _03216_, _02891_);
  not (_03218_, _03217_);
  not (_03219_, _03216_);
  and (_03220_, _02988_, _02943_);
  nor (_03221_, _03035_, _02874_);
  and (_03222_, _03221_, _02888_);
  nor (_03223_, _02895_, _02500_);
  and (_03225_, _03223_, _02939_);
  and (_03226_, _03225_, _03222_);
  and (_03227_, _03226_, _03220_);
  nor (_03228_, _03227_, _03219_);
  not (_03229_, _03228_);
  and (_03230_, _02750_, _33958_);
  and (_03231_, _02761_, _01379_);
  nor (_03232_, _03231_, _03230_);
  and (_03233_, _02756_, _01373_);
  and (_03234_, _02734_, _01366_);
  nor (_03235_, _03234_, _03233_);
  and (_03236_, _03235_, _03232_);
  and (_03237_, _02713_, _01389_);
  and (_03238_, _02718_, _01387_);
  nor (_03239_, _03238_, _03237_);
  and (_03240_, _02745_, _01360_);
  and (_03241_, _02763_, _01358_);
  nor (_03242_, _03241_, _03240_);
  and (_03243_, _03242_, _03239_);
  and (_03244_, _03243_, _03236_);
  and (_03245_, _02758_, _01396_);
  and (_03246_, _02737_, _01393_);
  nor (_03247_, _03246_, _03245_);
  and (_03248_, _02732_, _01368_);
  and (_03249_, _02724_, _01371_);
  nor (_03250_, _03249_, _03248_);
  and (_03251_, _03250_, _03247_);
  and (_03252_, _02752_, _01385_);
  and (_03253_, _02747_, _01362_);
  nor (_03254_, _03253_, _03252_);
  and (_03255_, _02728_, _01375_);
  and (_03256_, _02739_, _01398_);
  nor (_03257_, _03256_, _03255_);
  and (_03258_, _03257_, _03254_);
  and (_03259_, _03258_, _03251_);
  and (_03260_, _03259_, _03244_);
  not (_03261_, _03260_);
  nand (_03262_, _02997_, _02967_);
  nor (_03263_, _03262_, _02960_);
  nand (_03264_, _03263_, _02983_);
  nor (_03265_, _03174_, _03166_);
  and (_03266_, _03265_, _02901_);
  and (_03267_, _03266_, _03135_);
  nand (_03268_, _03267_, _03144_);
  or (_03269_, _03268_, _03264_);
  and (_03270_, _03269_, _03261_);
  not (_03271_, _03270_);
  and (_03272_, _03076_, _01375_);
  and (_03273_, _03094_, _01393_);
  nor (_03274_, _03273_, _03272_);
  and (_03275_, _03086_, _01366_);
  and (_03276_, _03096_, _01398_);
  nor (_03277_, _03276_, _03275_);
  and (_03278_, _03277_, _03274_);
  and (_03279_, _03083_, _01385_);
  and (_03280_, _03100_, _01360_);
  nor (_03281_, _03280_, _03279_);
  and (_03282_, _03107_, _33958_);
  and (_03283_, _03081_, _01387_);
  nor (_03284_, _03283_, _03282_);
  and (_03285_, _03284_, _03281_);
  and (_03286_, _03285_, _03278_);
  and (_03287_, _03114_, _01358_);
  and (_03288_, _03088_, _01371_);
  nor (_03289_, _03288_, _03287_);
  and (_03290_, _03112_, _01379_);
  and (_03291_, _03068_, _01396_);
  nor (_03292_, _03291_, _03290_);
  and (_03293_, _03292_, _03289_);
  and (_03294_, _03102_, _01362_);
  and (_03295_, _03063_, _01373_);
  nor (_03296_, _03295_, _03294_);
  and (_03297_, _03074_, _01389_);
  and (_03298_, _03109_, _01368_);
  nor (_03299_, _03298_, _03297_);
  and (_03300_, _03299_, _03296_);
  and (_03301_, _03300_, _03293_);
  and (_03302_, _03301_, _03286_);
  nor (_03303_, _03302_, _02851_);
  and (_03304_, _02837_, _02890_);
  not (_03305_, _03304_);
  and (_03306_, _02859_, _02890_);
  and (_03307_, _02835_, _02890_);
  nor (_03308_, _03307_, _03306_);
  and (_03309_, _03308_, _03305_);
  and (_03310_, _02859_, _02530_);
  and (_03311_, _02835_, _02530_);
  nor (_03312_, _03311_, _03310_);
  and (_03313_, _02834_, _02497_);
  not (_03314_, _03313_);
  not (_03316_, _02577_);
  and (_03317_, _03316_, _02560_);
  nor (_03318_, _03317_, _03314_);
  nor (_03319_, _03318_, _02836_);
  and (_03320_, _03319_, _03312_);
  and (_03321_, _03320_, _03309_);
  nor (_03322_, _02975_, _02562_);
  and (_03323_, _02859_, _02953_);
  nor (_03324_, _03323_, _03322_);
  not (_03325_, _03324_);
  not (_03326_, \oc8051_golden_model_1.SP [2]);
  not (_03327_, _02947_);
  nor (_03328_, _03148_, _02897_);
  and (_03329_, _03328_, _03327_);
  nor (_03330_, _03329_, _03326_);
  nor (_03331_, _03330_, _03325_);
  and (_03332_, _03331_, _03321_);
  and (_03333_, _03313_, _02532_);
  and (_03334_, _03313_, _02511_);
  nor (_03335_, _03334_, _03333_);
  and (_03336_, _02837_, _02885_);
  and (_03337_, _03313_, _02370_);
  nor (_03338_, _03337_, _03336_);
  and (_03339_, _03313_, _02535_);
  not (_03340_, _03339_);
  and (_03341_, _03340_, _03338_);
  and (_03342_, _03341_, _03335_);
  and (_03343_, _02837_, _02525_);
  and (_03344_, _02837_, _02535_);
  nor (_03345_, _03344_, _03343_);
  not (_03346_, _02837_);
  nor (_03347_, _02577_, _02511_);
  nor (_03348_, _03347_, _03346_);
  not (_03349_, _03348_);
  and (_03350_, _03349_, _03345_);
  and (_03351_, _02837_, _02370_);
  nor (_03352_, _02860_, _03351_);
  and (_03353_, _03352_, _03350_);
  and (_03354_, _02837_, _02530_);
  not (_03355_, _03354_);
  and (_03356_, _02837_, _02532_);
  nor (_03357_, _02838_, _03356_);
  and (_03358_, _03357_, _03355_);
  and (_03359_, _02837_, _02879_);
  and (_03360_, _02834_, _02537_);
  nor (_03361_, _03360_, _03359_);
  and (_03362_, _03313_, _02885_);
  and (_03363_, _03313_, _02525_);
  nor (_03364_, _03363_, _03362_);
  and (_03365_, _03364_, _03361_);
  and (_03366_, _03365_, _03358_);
  and (_03367_, _03366_, _03353_);
  and (_03368_, _03367_, _03342_);
  and (_03369_, _03368_, _03332_);
  not (_03370_, _03369_);
  nor (_03371_, _03370_, _03303_);
  and (_03372_, _03371_, _03271_);
  and (_03373_, _03372_, _03229_);
  and (_03374_, _03373_, _03218_);
  not (_03375_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_03376_, _02988_, _02800_);
  not (_03377_, _02966_);
  nor (_03378_, _02832_, _03377_);
  or (_03379_, _02832_, _02959_);
  nor (_03380_, _02832_, _02955_);
  nor (_03381_, _02854_, _02862_);
  nor (_03382_, _03381_, _02562_);
  not (_03383_, _02557_);
  and (_03384_, _02854_, _03383_);
  nor (_03385_, _03384_, _03382_);
  nor (_03386_, _03385_, _02545_);
  not (_03387_, _03386_);
  and (_03388_, _02841_, _02574_);
  and (_03389_, _03388_, _02890_);
  not (_03390_, _03389_);
  and (_03391_, _02873_, _02953_);
  not (_03392_, _03391_);
  and (_03393_, _02465_, _02432_);
  and (_03394_, _03393_, _02890_);
  nor (_03395_, _03394_, _02952_);
  and (_03396_, _03395_, _03392_);
  and (_03397_, _03396_, _03390_);
  and (_03398_, _02834_, _02465_);
  nor (_03399_, _02843_, _03398_);
  nor (_03400_, _03399_, _02562_);
  not (_03401_, _03400_);
  and (_03402_, _02873_, _03383_);
  nor (_03403_, _03402_, _02954_);
  and (_03404_, _03403_, _03401_);
  and (_03405_, _03404_, _03397_);
  and (_03406_, _03405_, _03387_);
  or (_03407_, _03406_, _03380_);
  nand (_03408_, _03407_, _02892_);
  nand (_03409_, _02893_, _03408_);
  and (_03410_, _02947_, _02877_);
  nor (_03411_, _03410_, _02950_);
  and (_03412_, _03393_, _02885_);
  and (_03413_, _02854_, _02885_);
  and (_03414_, _03413_, _02465_);
  nor (_03415_, _03414_, _03412_);
  and (_03416_, _03415_, _03411_);
  nand (_03417_, _03416_, _03409_);
  nand (_03418_, _03417_, _03379_);
  and (_03419_, _03418_, _02888_);
  or (_03420_, _02889_, _03419_);
  and (_03421_, _02832_, _02886_);
  not (_03422_, _02574_);
  nor (_03423_, _02841_, _02572_);
  nor (_03424_, _03423_, _03422_);
  nor (_03425_, _03424_, _03393_);
  nor (_03426_, _03425_, _02560_);
  nor (_03427_, _03426_, _03421_);
  and (_03428_, _03427_, _03420_);
  or (_03429_, _03428_, _03378_);
  and (_03430_, _03429_, _02943_);
  nor (_03431_, _02943_, _02800_);
  or (_03432_, _03431_, _03430_);
  and (_03433_, _02832_, _02984_);
  and (_03434_, _03388_, _02980_);
  nor (_03435_, _03434_, _02993_);
  not (_03436_, _03435_);
  nor (_03437_, _03436_, _03433_);
  and (_03438_, _03437_, _03432_);
  or (_03439_, _03438_, _03376_);
  nand (_03440_, _03398_, _02577_);
  and (_03441_, _02854_, _02577_);
  and (_03442_, _03441_, _02465_);
  and (_03443_, _02843_, _02577_);
  and (_03444_, _02862_, _02577_);
  or (_03445_, _03444_, _02992_);
  or (_03446_, _03445_, _03443_);
  nor (_03447_, _03446_, _03442_);
  and (_03448_, _03447_, _03440_);
  and (_03449_, _03448_, _03439_);
  nor (_03450_, _02832_, _02997_);
  or (_03451_, _03450_, _03449_);
  and (_03452_, _03451_, _02875_);
  or (_03453_, _03452_, _02876_);
  nor (_03454_, _02860_, _02576_);
  and (_03455_, _03017_, _02520_);
  and (_03456_, _03388_, _02520_);
  or (_03457_, _03456_, _02863_);
  or (_03458_, _03457_, _02844_);
  nor (_03459_, _03458_, _03455_);
  and (_03460_, _03459_, _03454_);
  and (_03461_, _03460_, _03453_);
  and (_03462_, _03076_, _01289_);
  and (_03463_, _03094_, _01297_);
  nor (_03464_, _03463_, _03462_);
  and (_03465_, _03086_, _01276_);
  and (_03466_, _03096_, _01268_);
  nor (_03467_, _03466_, _03465_);
  and (_03468_, _03467_, _03464_);
  and (_03469_, _03107_, _33944_);
  and (_03470_, _03074_, _01304_);
  nor (_03471_, _03470_, _03469_);
  and (_03472_, _03081_, _01302_);
  and (_03473_, _03100_, _01270_);
  nor (_03474_, _03473_, _03472_);
  and (_03475_, _03474_, _03471_);
  and (_03476_, _03475_, _03468_);
  and (_03477_, _03102_, _01300_);
  and (_03478_, _03088_, _01281_);
  nor (_03479_, _03478_, _03477_);
  and (_03480_, _03112_, _01283_);
  and (_03481_, _03068_, _01295_);
  nor (_03482_, _03481_, _03480_);
  and (_03483_, _03482_, _03479_);
  and (_03484_, _03114_, _01272_);
  and (_03485_, _03063_, _01285_);
  nor (_03486_, _03485_, _03484_);
  and (_03487_, _03083_, _01306_);
  and (_03488_, _03109_, _01278_);
  nor (_03489_, _03488_, _03487_);
  and (_03490_, _03489_, _03486_);
  and (_03491_, _03490_, _03483_);
  and (_03492_, _03491_, _03476_);
  nor (_03493_, _03492_, _02851_);
  or (_03494_, _03493_, _03461_);
  and (_03495_, _02938_, _02800_);
  and (_03496_, _03388_, _02516_);
  nor (_03497_, _03496_, _02937_);
  not (_03498_, _03497_);
  nor (_03499_, _03498_, _03495_);
  and (_03500_, _03499_, _03494_);
  not (_03501_, _02800_);
  and (_03502_, _02937_, _03501_);
  or (_03503_, _03502_, _03500_);
  and (_03504_, _03388_, _02511_);
  and (_03505_, _03393_, _02511_);
  nor (_03506_, _03505_, _03504_);
  and (_03507_, _03506_, _03503_);
  nor (_03508_, _02833_, _03134_);
  not (_03509_, _02532_);
  nor (_03510_, _03399_, _03509_);
  not (_03511_, _03510_);
  and (_03512_, _02862_, _02532_);
  and (_03513_, _02854_, _02532_);
  and (_03514_, _03513_, _02465_);
  nor (_03515_, _03514_, _03512_);
  and (_03517_, _03515_, _03511_);
  not (_03518_, _03517_);
  nor (_03519_, _03518_, _03508_);
  and (_03520_, _03519_, _03507_);
  nor (_03521_, _02833_, _03143_);
  and (_03522_, _03398_, _02537_);
  and (_03523_, _02843_, _02537_);
  and (_03524_, _03388_, _02537_);
  and (_03525_, _02862_, _02537_);
  or (_03526_, _03525_, _03524_);
  or (_03527_, _03526_, _03523_);
  nor (_03528_, _03527_, _03522_);
  not (_03529_, _03528_);
  nor (_03530_, _03529_, _03521_);
  and (_03531_, _03530_, _03520_);
  nor (_03532_, _02833_, _03129_);
  and (_03533_, _03388_, _02530_);
  not (_03534_, _03533_);
  and (_03535_, _02843_, _02530_);
  nor (_03536_, _03535_, _03310_);
  not (_03537_, _02530_);
  nor (_03538_, _03017_, _02575_);
  and (_03539_, _03538_, _03031_);
  or (_03540_, _03539_, _03537_);
  and (_03541_, _03540_, _03536_);
  and (_03542_, _03541_, _03534_);
  not (_03543_, _03542_);
  nor (_03544_, _03543_, _03532_);
  and (_03545_, _03544_, _03531_);
  nor (_03546_, _02832_, _03138_);
  or (_03547_, _03546_, _03545_);
  and (_03548_, _03148_, _02877_);
  nor (_03549_, _03548_, _03035_);
  and (_03550_, _03549_, _03547_);
  nor (_03551_, _03152_, _02800_);
  nor (_03552_, _03551_, _03550_);
  not (_03553_, _02535_);
  nor (_03554_, _03425_, _03553_);
  nor (_03555_, _03554_, _03552_);
  nor (_03556_, _02832_, _02901_);
  or (_03557_, _03556_, _03555_);
  and (_03558_, _02897_, _02877_);
  nor (_03559_, _03558_, _02895_);
  and (_03560_, _03559_, _03557_);
  nor (_03561_, _02896_, _02800_);
  or (_03562_, _03561_, _03560_);
  not (_03563_, _03166_);
  and (_03564_, _03017_, _02370_);
  not (_03565_, _03564_);
  and (_03566_, _02859_, _02370_);
  and (_03567_, _02843_, _02370_);
  nor (_03568_, _03567_, _03566_);
  and (_03569_, _03568_, _03565_);
  and (_03570_, _02862_, _02370_);
  and (_03571_, _03388_, _02370_);
  nor (_03572_, _03571_, _03570_);
  and (_03573_, _03572_, _03569_);
  and (_03574_, _03573_, _03563_);
  and (_03575_, _03574_, _03562_);
  nor (_03576_, _02832_, _03563_);
  or (_03577_, _03576_, _03575_);
  and (_03578_, _03577_, _02501_);
  or (_03579_, _03578_, _02801_);
  and (_03580_, _02842_, _02525_);
  nor (_03581_, _03580_, _03343_);
  nor (_03582_, _03581_, _02545_);
  not (_03583_, _03582_);
  and (_03584_, _02859_, _02525_);
  not (_03585_, _03584_);
  and (_03586_, _03388_, _02525_);
  nor (_03587_, _03586_, _03174_);
  and (_03588_, _03587_, _03585_);
  and (_03589_, _03588_, _03583_);
  nand (_03590_, _03589_, _03579_);
  nor (_03591_, _02832_, _03178_);
  not (_03592_, _03591_);
  nand (_03593_, _03592_, _03590_);
  or (_03594_, _03593_, _03375_);
  and (_03595_, _02747_, _01448_);
  and (_03596_, _02724_, _01480_);
  nor (_03597_, _03596_, _03595_);
  and (_03598_, _02750_, _33972_);
  and (_03599_, _02756_, _01464_);
  nor (_03600_, _03599_, _03598_);
  and (_03601_, _03600_, _03597_);
  and (_03602_, _02763_, _01450_);
  and (_03603_, _02734_, _01475_);
  nor (_03604_, _03603_, _03602_);
  and (_03605_, _02728_, _01478_);
  and (_03606_, _02758_, _01488_);
  nor (_03607_, _03606_, _03605_);
  and (_03608_, _03607_, _03604_);
  and (_03609_, _03608_, _03601_);
  and (_03610_, _02718_, _01458_);
  and (_03611_, _02761_, _01466_);
  nor (_03612_, _03611_, _03610_);
  and (_03613_, _02732_, _01473_);
  and (_03614_, _02737_, _01486_);
  nor (_03615_, _03614_, _03613_);
  and (_03616_, _03615_, _03612_);
  and (_03617_, _02752_, _01456_);
  and (_03618_, _02745_, _01452_);
  nor (_03619_, _03618_, _03617_);
  and (_03620_, _02713_, _01460_);
  and (_03621_, _02739_, _01471_);
  nor (_03622_, _03621_, _03620_);
  and (_03623_, _03622_, _03619_);
  and (_03624_, _03623_, _03616_);
  and (_03625_, _03624_, _03609_);
  nor (_03626_, _02875_, _02768_);
  nor (_03627_, _02768_, _02501_);
  nor (_03628_, _03627_, _03626_);
  nor (_03629_, _03628_, _03625_);
  not (_03630_, _03629_);
  nor (_03631_, _03625_, _02768_);
  and (_03632_, _03631_, _02891_);
  not (_03633_, _03632_);
  nor (_03634_, _03035_, _02895_);
  and (_03635_, _03634_, _02888_);
  and (_03636_, _03635_, _02939_);
  and (_03637_, _03636_, _03220_);
  not (_03638_, _03637_);
  and (_03639_, _03638_, _03631_);
  not (_03640_, _03639_);
  and (_03641_, _02745_, _01315_);
  and (_03642_, _02763_, _01317_);
  nor (_03643_, _03642_, _03641_);
  and (_03644_, _02756_, _01323_);
  and (_03645_, _02728_, _01325_);
  nor (_03646_, _03645_, _03644_);
  and (_03647_, _03646_, _03643_);
  and (_03648_, _02737_, _01340_);
  and (_03649_, _02739_, _01353_);
  nor (_03650_, _03649_, _03648_);
  and (_03651_, _02734_, _01334_);
  and (_03652_, _02724_, _01336_);
  nor (_03653_, _03652_, _03651_);
  and (_03654_, _03653_, _03650_);
  and (_03655_, _03654_, _03647_);
  and (_03656_, _02750_, _33951_);
  and (_03657_, _02747_, _01313_);
  nor (_03658_, _03657_, _03656_);
  and (_03659_, _02718_, _01344_);
  and (_03660_, _02761_, _01329_);
  nor (_03661_, _03660_, _03659_);
  and (_03662_, _03661_, _03658_);
  and (_03663_, _02732_, _01321_);
  and (_03664_, _02758_, _01351_);
  nor (_03665_, _03664_, _03663_);
  and (_03666_, _02713_, _01342_);
  and (_03667_, _02752_, _01347_);
  nor (_03668_, _03667_, _03666_);
  and (_03669_, _03668_, _03665_);
  and (_03670_, _03669_, _03662_);
  and (_03671_, _03670_, _03655_);
  not (_03672_, _03671_);
  and (_03673_, _03672_, _03269_);
  not (_03674_, _03673_);
  and (_03675_, _03112_, _01329_);
  and (_03676_, _03068_, _01351_);
  nor (_03677_, _03676_, _03675_);
  and (_03678_, _03107_, _33951_);
  and (_03679_, _03088_, _01336_);
  nor (_03680_, _03679_, _03678_);
  and (_03681_, _03680_, _03677_);
  and (_03682_, _03100_, _01315_);
  and (_03683_, _03114_, _01317_);
  nor (_03684_, _03683_, _03682_);
  and (_03685_, _03074_, _01342_);
  and (_03686_, _03076_, _01325_);
  nor (_03687_, _03686_, _03685_);
  and (_03688_, _03687_, _03684_);
  and (_03689_, _03688_, _03681_);
  and (_03690_, _03063_, _01323_);
  and (_03691_, _03109_, _01321_);
  nor (_03692_, _03691_, _03690_);
  and (_03693_, _03086_, _01334_);
  and (_03694_, _03096_, _01353_);
  nor (_03695_, _03694_, _03693_);
  and (_03696_, _03695_, _03692_);
  and (_03697_, _03102_, _01313_);
  and (_03698_, _03094_, _01340_);
  nor (_03699_, _03698_, _03697_);
  and (_03700_, _03081_, _01344_);
  and (_03701_, _03083_, _01347_);
  nor (_03702_, _03701_, _03700_);
  and (_03703_, _03702_, _03699_);
  and (_03704_, _03703_, _03696_);
  and (_03705_, _03704_, _03689_);
  nor (_03706_, _03705_, _02851_);
  nor (_03707_, _02838_, _03359_);
  and (_03708_, _03707_, _03345_);
  nor (_03709_, _03351_, _03348_);
  and (_03710_, _03709_, _03708_);
  and (_03711_, _03010_, _02370_);
  and (_03712_, _03010_, _02953_);
  nor (_03713_, _03712_, _03711_);
  and (_03714_, _03010_, _02885_);
  and (_03715_, _03010_, _02537_);
  nor (_03716_, _03715_, _03714_);
  and (_03718_, _03716_, _03713_);
  and (_03719_, _02837_, _02953_);
  nor (_03720_, _03336_, _03719_);
  nor (_03721_, _03356_, _03354_);
  and (_03722_, _03721_, _03720_);
  and (_03723_, _03722_, _03718_);
  and (_03724_, _03723_, _03710_);
  nor (_03725_, _03304_, _03010_);
  and (_03726_, _02560_, _02555_);
  nand (_03727_, _02336_, _02305_);
  and (_03728_, _03727_, _03726_);
  and (_03729_, _02577_, _02545_);
  not (_03730_, _03729_);
  nor (_03731_, _02532_, _02530_);
  and (_03732_, _03731_, _03730_);
  and (_03733_, _03732_, _03728_);
  nor (_03734_, _03733_, _03725_);
  not (_03735_, _03734_);
  and (_03736_, _02837_, _02537_);
  and (_03737_, _03148_, \oc8051_golden_model_1.SP [1]);
  nor (_03738_, _03737_, _03736_);
  and (_03739_, _02897_, \oc8051_golden_model_1.SP [1]);
  and (_03740_, _02947_, \oc8051_golden_model_1.SP [1]);
  nor (_03741_, _03740_, _03739_);
  and (_03742_, _03741_, _03738_);
  nor (_03743_, _02844_, _03443_);
  and (_03744_, _02843_, _02511_);
  not (_03745_, _02845_);
  nor (_03746_, _02520_, _02511_);
  nor (_03747_, _03746_, _03745_);
  nor (_03748_, _03747_, _03744_);
  and (_03749_, _03748_, _03743_);
  and (_03750_, _03749_, _03742_);
  and (_03751_, _03750_, _03735_);
  and (_03752_, _03751_, _03724_);
  not (_03753_, _03752_);
  nor (_03754_, _03753_, _03706_);
  and (_03755_, _03754_, _03674_);
  and (_03756_, _03755_, _03640_);
  and (_03757_, _03756_, _03633_);
  and (_03758_, _03757_, _03630_);
  not (_03759_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_03760_, _03592_, _03590_);
  or (_03761_, _03760_, _03759_);
  and (_03762_, _03761_, _03758_);
  nand (_03763_, _03762_, _03594_);
  not (_03764_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_03765_, _03760_, _03764_);
  not (_03766_, _03758_);
  not (_03767_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_03768_, _03593_, _03767_);
  and (_03769_, _03768_, _03766_);
  nand (_03770_, _03769_, _03765_);
  nand (_03771_, _03770_, _03763_);
  nand (_03772_, _03771_, _03374_);
  not (_03773_, _03374_);
  not (_03774_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_03775_, _03760_, _03774_);
  not (_03776_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_03777_, _03593_, _03776_);
  and (_03778_, _03777_, _03766_);
  nand (_03779_, _03778_, _03775_);
  not (_03780_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_03781_, _03593_, _03780_);
  not (_03782_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_03783_, _03760_, _03782_);
  and (_03784_, _03783_, _03758_);
  nand (_03785_, _03784_, _03781_);
  nand (_03786_, _03785_, _03779_);
  nand (_03787_, _03786_, _03773_);
  nand (_03788_, _03787_, _03772_);
  nand (_03789_, _03788_, _03181_);
  not (_03790_, _03181_);
  not (_03791_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03792_, _03760_, _03791_);
  nand (_03793_, _03760_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03794_, _03793_, _03766_);
  nand (_03795_, _03794_, _03792_);
  not (_03796_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03797_, _03593_, _03796_);
  nand (_03798_, _03593_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03799_, _03798_, _03758_);
  nand (_03800_, _03799_, _03797_);
  nand (_03801_, _03800_, _03795_);
  nand (_03802_, _03801_, _03374_);
  not (_03803_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03804_, _03760_, _03803_);
  nand (_03805_, _03760_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03806_, _03805_, _03766_);
  nand (_03807_, _03806_, _03804_);
  not (_03808_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03809_, _03593_, _03808_);
  nand (_03810_, _03593_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_03811_, _03810_, _03758_);
  nand (_03812_, _03811_, _03809_);
  nand (_03813_, _03812_, _03807_);
  nand (_03814_, _03813_, _03773_);
  nand (_03815_, _03814_, _03802_);
  nand (_03816_, _03815_, _03790_);
  and (_03817_, _03816_, _03789_);
  and (_03818_, _02854_, _02890_);
  nor (_03819_, _03818_, _03384_);
  or (_03820_, _03819_, _03817_);
  not (_03821_, _02952_);
  nor (_03822_, _03821_, _02768_);
  not (_03823_, _03822_);
  not (_03824_, _02558_);
  and (_03825_, _02575_, _03383_);
  not (_03826_, _03825_);
  nor (_03827_, _03826_, _02768_);
  and (_03828_, _03827_, _02833_);
  or (_03829_, _03828_, _03824_);
  and (_03830_, _03393_, _03383_);
  nor (_03831_, _03830_, _03827_);
  or (_03832_, _03831_, _03829_);
  nor (_03833_, _02558_, _02877_);
  nor (_03834_, _03833_, _03394_);
  and (_03835_, _03834_, _03832_);
  and (_03836_, _03835_, _03823_);
  and (_03837_, _03836_, _03820_);
  and (_03838_, _03822_, _02833_);
  nor (_03839_, _03838_, _03837_);
  nor (_03840_, _03839_, _02894_);
  not (_03841_, _03840_);
  and (_03842_, _03841_, _02893_);
  nor (_03843_, _02556_, _02877_);
  nor (_03844_, _03843_, _03842_);
  nor (_03845_, _03327_, _02768_);
  and (_03846_, _03845_, _02832_);
  nor (_03847_, _03846_, _03412_);
  and (_03848_, _03847_, _03844_);
  not (_03849_, _03413_);
  nor (_03850_, _03817_, _03849_);
  not (_03851_, _03850_);
  and (_03852_, _03851_, _03848_);
  nor (_03853_, _02888_, _02768_);
  nor (_03854_, _02959_, _02768_);
  and (_03855_, _03854_, _02832_);
  nor (_03856_, _03855_, _03853_);
  and (_03857_, _03856_, _03852_);
  nor (_03858_, _03857_, _02889_);
  nor (_03859_, _03858_, _02886_);
  and (_03860_, _02886_, _02877_);
  or (_03861_, _03860_, _03859_);
  and (_03862_, _03861_, _02884_);
  nor (_03863_, _03862_, _02882_);
  and (_03864_, _03393_, _02980_);
  or (_03865_, _03864_, _03863_);
  nor (_03866_, _03865_, _02878_);
  and (_03867_, _02854_, _02980_);
  not (_03868_, _03817_);
  and (_03869_, _03868_, _03867_);
  nor (_03870_, _03869_, _03626_);
  and (_03871_, _03870_, _03866_);
  nor (_03872_, _03871_, _02876_);
  nor (_03873_, _03872_, _02578_);
  and (_03874_, _02578_, _02877_);
  nor (_03875_, _03874_, _03873_);
  and (_03876_, _03393_, _02516_);
  or (_03877_, _03876_, _03875_);
  nor (_03878_, _03877_, _02872_);
  and (_03879_, _02854_, _02516_);
  not (_03880_, _03879_);
  nor (_03881_, _03817_, _03880_);
  not (_03882_, _03881_);
  and (_03883_, _03882_, _03878_);
  not (_03884_, _03014_);
  nor (_03885_, _03884_, _02768_);
  and (_03886_, _03885_, _02832_);
  nor (_03887_, _03886_, _02517_);
  and (_03888_, _03887_, _03883_);
  and (_03889_, _02517_, _02877_);
  nor (_03890_, _03889_, _03888_);
  nor (_03891_, _03140_, _02768_);
  and (_03892_, _03131_, _03022_);
  nor (_03893_, _03892_, _02768_);
  nor (_03894_, _03893_, _03891_);
  nor (_03895_, _03894_, _02833_);
  nor (_03896_, _03895_, _02533_);
  not (_03897_, _03896_);
  nor (_03898_, _03897_, _03890_);
  and (_03899_, _02533_, _02877_);
  nor (_03900_, _03899_, _03898_);
  nor (_03901_, _03128_, _02768_);
  and (_03902_, _03901_, _02832_);
  nor (_03903_, _03902_, _03900_);
  and (_03904_, _03393_, _02370_);
  and (_03905_, _02531_, \oc8051_golden_model_1.SP [0]);
  nor (_03906_, _03905_, _03904_);
  and (_03907_, _03906_, _03903_);
  nor (_03908_, _03563_, _02768_);
  and (_03909_, _02854_, _02370_);
  not (_03910_, _03909_);
  nor (_03911_, _03817_, _03910_);
  nor (_03912_, _03911_, _03908_);
  and (_03913_, _03912_, _03907_);
  and (_03914_, _03908_, _02833_);
  nor (_03915_, _03914_, _03913_);
  nor (_03916_, _03004_, _02528_);
  nor (_03917_, _03916_, _02877_);
  nor (_03919_, _03917_, _03627_);
  not (_03920_, _03919_);
  nor (_03921_, _03920_, _03915_);
  nor (_03922_, _03921_, _02801_);
  and (_03923_, _03393_, _02525_);
  nor (_03924_, _03923_, _03922_);
  nor (_03925_, _03178_, _02768_);
  and (_03926_, _02854_, _02525_);
  not (_03927_, _03926_);
  nor (_03928_, _03817_, _03927_);
  nor (_03929_, _03928_, _03925_);
  and (_03930_, _03929_, _03924_);
  and (_03931_, _03925_, _02833_);
  nor (_03932_, _03931_, _03930_);
  not (_03933_, _03932_);
  and (_03934_, _03925_, _03672_);
  and (_03935_, _03631_, _02500_);
  not (_03936_, _03627_);
  not (_03937_, \oc8051_golden_model_1.SP [1]);
  and (_03938_, _03937_, \oc8051_golden_model_1.SP [0]);
  and (_03939_, \oc8051_golden_model_1.SP [1], _02877_);
  nor (_03940_, _03939_, _03938_);
  not (_03941_, _03940_);
  and (_03942_, _03941_, _02531_);
  and (_03943_, _03885_, _03672_);
  nor (_03944_, _02871_, _03672_);
  and (_03945_, _03631_, _02874_);
  and (_03946_, _03941_, _02886_);
  not (_03947_, _02886_);
  and (_03948_, _03822_, _03672_);
  not (_03949_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03950_, _03593_, _03949_);
  not (_03951_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_03952_, _03760_, _03951_);
  and (_03953_, _03952_, _03758_);
  nand (_03954_, _03953_, _03950_);
  not (_03955_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03956_, _03760_, _03955_);
  not (_03957_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03958_, _03593_, _03957_);
  and (_03959_, _03958_, _03766_);
  nand (_03960_, _03959_, _03956_);
  nand (_03961_, _03960_, _03954_);
  nand (_03962_, _03961_, _03374_);
  not (_03963_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03964_, _03760_, _03963_);
  not (_03965_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03966_, _03593_, _03965_);
  and (_03967_, _03966_, _03766_);
  nand (_03968_, _03967_, _03964_);
  not (_03969_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03970_, _03593_, _03969_);
  not (_03971_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03972_, _03760_, _03971_);
  and (_03973_, _03972_, _03758_);
  nand (_03974_, _03973_, _03970_);
  nand (_03975_, _03974_, _03968_);
  nand (_03976_, _03975_, _03773_);
  nand (_03977_, _03976_, _03962_);
  nand (_03978_, _03977_, _03181_);
  not (_03979_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03980_, _03760_, _03979_);
  nand (_03981_, _03760_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03982_, _03981_, _03766_);
  nand (_03983_, _03982_, _03980_);
  not (_03984_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_03985_, _03593_, _03984_);
  nand (_03986_, _03593_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03987_, _03986_, _03758_);
  nand (_03988_, _03987_, _03985_);
  nand (_03989_, _03988_, _03983_);
  nand (_03990_, _03989_, _03374_);
  not (_03991_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_03992_, _03760_, _03991_);
  nand (_03993_, _03760_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_03994_, _03993_, _03766_);
  nand (_03995_, _03994_, _03992_);
  not (_03996_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03997_, _03593_, _03996_);
  nand (_03998_, _03593_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_03999_, _03998_, _03758_);
  nand (_04000_, _03999_, _03997_);
  nand (_04001_, _04000_, _03995_);
  nand (_04002_, _04001_, _03773_);
  nand (_04003_, _04002_, _03990_);
  nand (_04004_, _04003_, _03790_);
  and (_04005_, _04004_, _03978_);
  or (_04006_, _04005_, _03819_);
  and (_04007_, _02497_, _02432_);
  and (_04008_, _04007_, _03383_);
  nor (_04009_, _04008_, _03827_);
  and (_04010_, _03827_, _03672_);
  or (_04011_, _04010_, _03824_);
  or (_04012_, _04011_, _04009_);
  and (_04013_, _03313_, _02890_);
  and (_04014_, _02862_, _02890_);
  and (_04015_, _02864_, _02890_);
  nor (_04016_, _04015_, _04014_);
  nor (_04017_, _03941_, _02558_);
  not (_04018_, _04017_);
  nand (_04019_, _04018_, _04016_);
  nor (_04020_, _04019_, _04013_);
  and (_04021_, _04020_, _04012_);
  and (_04022_, _04021_, _03823_);
  and (_04023_, _04022_, _04006_);
  nor (_04024_, _04023_, _03948_);
  nor (_04025_, _04024_, _02894_);
  nor (_04026_, _04025_, _03632_);
  nor (_04027_, _03941_, _02556_);
  nor (_04028_, _04027_, _04026_);
  and (_04029_, _03845_, _03671_);
  and (_04030_, _02864_, _02885_);
  not (_04031_, _04030_);
  and (_04032_, _02862_, _02885_);
  nor (_04033_, _04032_, _03362_);
  and (_04034_, _04033_, _04031_);
  not (_04035_, _04034_);
  nor (_04036_, _04035_, _04029_);
  and (_04037_, _04036_, _04028_);
  nand (_04038_, _04004_, _03978_);
  and (_04039_, _04038_, _03413_);
  nor (_04040_, _04039_, _03854_);
  and (_04041_, _04040_, _04037_);
  and (_04042_, _03854_, _03672_);
  nor (_04043_, _04042_, _04041_);
  and (_04044_, _03625_, _03853_);
  nor (_04045_, _04044_, _04043_);
  and (_04046_, _04045_, _03947_);
  nor (_04047_, _04046_, _03946_);
  and (_04048_, _03625_, _02883_);
  or (_04049_, _04048_, _04047_);
  nor (_04050_, _03941_, _02561_);
  and (_04051_, _04007_, _02980_);
  nor (_04052_, _04051_, _04050_);
  not (_04053_, _04052_);
  nor (_04054_, _04053_, _04049_);
  and (_04055_, _04038_, _03867_);
  nor (_04056_, _04055_, _03626_);
  and (_04057_, _04056_, _04054_);
  nor (_04058_, _04057_, _03945_);
  nor (_04059_, _04058_, _02578_);
  and (_04060_, _03941_, _02578_);
  nor (_04061_, _04060_, _04059_);
  and (_04062_, _04007_, _02516_);
  or (_04063_, _04062_, _04061_);
  nor (_04064_, _04063_, _03944_);
  and (_04065_, _04038_, _03879_);
  nor (_04066_, _04065_, _03885_);
  and (_04067_, _04066_, _04064_);
  nor (_04068_, _04067_, _03943_);
  nor (_04069_, _04068_, _02517_);
  and (_04070_, _03941_, _02517_);
  nor (_04071_, _04070_, _04069_);
  nor (_04072_, _03894_, _03672_);
  nor (_04073_, _04072_, _02533_);
  not (_04074_, _04073_);
  nor (_04075_, _04074_, _04071_);
  and (_04076_, _03941_, _02533_);
  nor (_04077_, _04076_, _04075_);
  and (_04078_, _03901_, _03671_);
  nor (_04079_, _04078_, _02531_);
  not (_04080_, _04079_);
  nor (_04081_, _04080_, _04077_);
  nor (_04082_, _04081_, _03942_);
  and (_04083_, _02864_, _02370_);
  nor (_04084_, _04083_, _03570_);
  not (_04085_, _04084_);
  nor (_04086_, _04085_, _03337_);
  not (_04087_, _04086_);
  nor (_04088_, _04087_, _04082_);
  and (_04089_, _04038_, _03909_);
  nor (_04090_, _04089_, _03908_);
  and (_04091_, _04090_, _04088_);
  and (_04092_, _03908_, _03672_);
  nor (_04093_, _04092_, _04091_);
  nor (_04094_, _03941_, _03916_);
  nor (_04095_, _04094_, _04093_);
  and (_04096_, _04095_, _03936_);
  nor (_04097_, _04096_, _03935_);
  and (_04098_, _04007_, _02525_);
  nor (_04099_, _04098_, _04097_);
  and (_04100_, _04038_, _03926_);
  nor (_04101_, _04100_, _03925_);
  and (_04102_, _04101_, _04099_);
  nor (_04103_, _04102_, _03934_);
  not (_04104_, _00000_);
  nor (_04105_, _03885_, _03853_);
  nor (_04106_, _03854_, _03845_);
  and (_04107_, _04106_, _04105_);
  nor (_04108_, _04030_, _03714_);
  and (_04109_, _03017_, _02980_);
  and (_04110_, _02842_, _02516_);
  and (_04111_, _04110_, _02502_);
  nor (_04112_, _04111_, _04109_);
  and (_04113_, _04112_, _04108_);
  not (_04114_, _04016_);
  and (_04115_, _04110_, _02572_);
  nor (_04116_, _04115_, _04114_);
  and (_04117_, _02981_, _02497_);
  not (_04118_, _04117_);
  and (_04120_, _04084_, _04118_);
  and (_04121_, _04120_, _04116_);
  and (_04122_, _04121_, _04113_);
  not (_04123_, _02517_);
  and (_04124_, _02534_, _04123_);
  not (_04125_, _02561_);
  nor (_04126_, _02578_, _04125_);
  and (_04127_, _04126_, _02559_);
  and (_04128_, _04127_, _04124_);
  and (_04129_, _04128_, _03309_);
  and (_04130_, _04129_, _04122_);
  and (_04131_, _02981_, _02496_);
  and (_04132_, _04131_, _02465_);
  not (_04133_, _04132_);
  nor (_04134_, _03030_, _02565_);
  not (_04135_, _04134_);
  and (_04136_, _02845_, _02525_);
  nor (_04137_, _04136_, _03584_);
  and (_04138_, _04137_, _04135_);
  and (_04139_, _04138_, _04133_);
  and (_04140_, _03010_, _02890_);
  not (_04141_, _02525_);
  nor (_04142_, _02975_, _04141_);
  nor (_04143_, _04142_, _04140_);
  and (_04144_, _02834_, _02516_);
  and (_04145_, _02834_, _03383_);
  nor (_04146_, _04145_, _04144_);
  and (_04147_, _04146_, _04143_);
  and (_04148_, _02842_, _02979_);
  and (_04149_, _04148_, _02525_);
  nor (_04150_, _04149_, _03867_);
  and (_04151_, _02842_, _03383_);
  nor (_04152_, _04151_, _04032_);
  and (_04153_, _04152_, _04150_);
  and (_04154_, _04153_, _04147_);
  nor (_04155_, _02976_, _02565_);
  not (_04156_, _04155_);
  and (_04157_, _04156_, _03338_);
  and (_04158_, _04157_, _04154_);
  not (_04159_, _03916_);
  nor (_04160_, _04159_, _03351_);
  and (_04161_, _04160_, _03927_);
  nor (_04162_, _03711_, _03413_);
  and (_04163_, _04162_, _03819_);
  nor (_04164_, _03909_, _03879_);
  nor (_04165_, _03362_, _02886_);
  and (_04166_, _04165_, _04164_);
  and (_04167_, _04166_, _04163_);
  and (_04168_, _04167_, _04161_);
  and (_04169_, _04168_, _04158_);
  and (_04170_, _04169_, _04139_);
  and (_04171_, _04170_, _04130_);
  not (_04172_, _04171_);
  nor (_04173_, _04172_, _03901_);
  and (_04174_, _04173_, _03628_);
  and (_04175_, _04174_, _04107_);
  not (_04176_, _03925_);
  nor (_04177_, _03908_, _02849_);
  and (_04178_, _04177_, _04176_);
  nor (_04179_, _03822_, _02894_);
  nor (_04180_, _03827_, _02883_);
  and (_04181_, _04180_, _04179_);
  and (_04182_, _04181_, _04178_);
  and (_04183_, _03894_, _02870_);
  and (_04184_, _04183_, _04182_);
  and (_04185_, _04184_, _04175_);
  nor (_04186_, _04185_, _04104_);
  not (_04187_, _04186_);
  nor (_04188_, _04187_, _04103_);
  and (_04189_, _04188_, _03933_);
  not (_04190_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04191_, _03593_, _04190_);
  not (_04192_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_04193_, _03760_, _04192_);
  and (_04194_, _04193_, _03758_);
  nand (_04195_, _04194_, _04191_);
  not (_04196_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_04197_, _03760_, _04196_);
  not (_04198_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04199_, _03593_, _04198_);
  and (_04200_, _04199_, _03766_);
  nand (_04201_, _04200_, _04197_);
  nand (_04202_, _04201_, _04195_);
  nand (_04203_, _04202_, _03374_);
  not (_04204_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04205_, _03760_, _04204_);
  not (_04206_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04207_, _03593_, _04206_);
  and (_04208_, _04207_, _03766_);
  nand (_04209_, _04208_, _04205_);
  not (_04210_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04211_, _03593_, _04210_);
  not (_04212_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04213_, _03760_, _04212_);
  and (_04214_, _04213_, _03758_);
  nand (_04215_, _04214_, _04211_);
  nand (_04216_, _04215_, _04209_);
  nand (_04217_, _04216_, _03773_);
  nand (_04218_, _04217_, _04203_);
  nand (_04219_, _04218_, _03181_);
  nand (_04220_, _03593_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04221_, _03760_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04222_, _04221_, _03766_);
  nand (_04223_, _04222_, _04220_);
  nand (_04224_, _03760_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04225_, _03593_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04226_, _04225_, _03758_);
  nand (_04227_, _04226_, _04224_);
  nand (_04228_, _04227_, _04223_);
  nand (_04229_, _04228_, _03374_);
  nand (_04230_, _03593_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04231_, _03760_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04232_, _04231_, _03766_);
  nand (_04233_, _04232_, _04230_);
  nand (_04234_, _03760_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_04235_, _03593_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04236_, _04235_, _03758_);
  nand (_04237_, _04236_, _04234_);
  nand (_04238_, _04237_, _04233_);
  nand (_04239_, _04238_, _03773_);
  nand (_04240_, _04239_, _04229_);
  nand (_04241_, _04240_, _03790_);
  nand (_04242_, _04241_, _04219_);
  and (_04243_, _04242_, _03926_);
  and (_04244_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04245_, _04244_, \oc8051_golden_model_1.SP [2]);
  or (_04246_, _04245_, \oc8051_golden_model_1.SP [3]);
  and (_04247_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04248_, _04247_, \oc8051_golden_model_1.SP [3]);
  nand (_04249_, _04248_, \oc8051_golden_model_1.SP [0]);
  and (_04250_, _04249_, _04246_);
  nor (_04251_, _04250_, _03916_);
  and (_04252_, _04242_, _03879_);
  not (_04253_, _04250_);
  nor (_04254_, _04253_, _02561_);
  and (_04255_, _04242_, _03413_);
  not (_04256_, _03845_);
  and (_04257_, _02932_, _02894_);
  nor (_04258_, _04253_, _02558_);
  nor (_04259_, _03384_, \oc8051_golden_model_1.PSW [3]);
  and (_04260_, _04242_, _03384_);
  or (_04261_, _04260_, _03827_);
  nor (_04262_, _04261_, _04259_);
  nor (_04263_, _03826_, _02800_);
  nor (_04264_, _04263_, _04262_);
  nor (_04265_, _04264_, _03824_);
  or (_04266_, _04265_, _03818_);
  nor (_04267_, _04266_, _04258_);
  and (_04268_, _04242_, _03818_);
  nor (_04269_, _04268_, _03822_);
  not (_04270_, _04269_);
  nor (_04271_, _04270_, _04267_);
  nor (_04272_, _03821_, _02800_);
  or (_04273_, _04272_, _02894_);
  nor (_04274_, _04273_, _04271_);
  nor (_04275_, _04274_, _04257_);
  and (_04276_, _04275_, _02556_);
  nor (_04277_, _04253_, _02556_);
  or (_04278_, _04277_, _04276_);
  and (_04279_, _04278_, _04256_);
  and (_04280_, _03845_, _02934_);
  or (_04281_, _04280_, _03413_);
  nor (_04282_, _04281_, _04279_);
  or (_04283_, _04282_, _03854_);
  nor (_04284_, _04283_, _04255_);
  and (_04285_, _03854_, _02934_);
  or (_04286_, _04285_, _03853_);
  nor (_04287_, _04286_, _04284_);
  and (_04288_, _02932_, _03853_);
  nor (_04289_, _04288_, _04287_);
  and (_04290_, _04289_, _03947_);
  and (_04291_, _04250_, _02886_);
  nor (_04292_, _04291_, _04290_);
  nor (_04293_, _04292_, _02883_);
  nor (_04294_, _02884_, _02936_);
  or (_04295_, _04294_, _04293_);
  and (_04296_, _04295_, _02561_);
  or (_04297_, _04296_, _03867_);
  nor (_04298_, _04297_, _04254_);
  and (_04299_, _04242_, _03867_);
  nor (_04300_, _04299_, _03626_);
  not (_04301_, _04300_);
  nor (_04302_, _04301_, _04298_);
  not (_04303_, _03626_);
  nor (_04304_, _04303_, _02936_);
  nor (_04305_, _04304_, _04302_);
  nor (_04306_, _04305_, _02578_);
  and (_04307_, _04250_, _02578_);
  not (_04308_, _04307_);
  and (_04309_, _04308_, _02871_);
  not (_04310_, _04309_);
  nor (_04311_, _04310_, _04306_);
  nor (_04312_, _02871_, _02934_);
  nor (_04313_, _04312_, _04311_);
  nor (_04314_, _04313_, _03879_);
  or (_04315_, _04314_, _03885_);
  nor (_04316_, _04315_, _04252_);
  and (_04317_, _03885_, _02934_);
  nor (_04318_, _04317_, _04316_);
  nor (_04319_, _04318_, _02517_);
  and (_04321_, _04250_, _02517_);
  not (_04322_, _04321_);
  and (_04323_, _04322_, _03894_);
  not (_04324_, _04323_);
  nor (_04325_, _04324_, _04319_);
  nor (_04326_, _03894_, _02934_);
  nor (_04327_, _04326_, _02533_);
  not (_04328_, _04327_);
  nor (_04329_, _04328_, _04325_);
  and (_04330_, _04250_, _02533_);
  nor (_04331_, _04330_, _03901_);
  not (_04332_, _04331_);
  nor (_04333_, _04332_, _04329_);
  and (_04334_, _03901_, _02799_);
  nor (_04335_, _04334_, _02531_);
  not (_04336_, _04335_);
  nor (_04337_, _04336_, _04333_);
  and (_04338_, _04250_, _02531_);
  nor (_04339_, _04338_, _03909_);
  not (_04340_, _04339_);
  nor (_04341_, _04340_, _04337_);
  and (_04342_, _04242_, _03909_);
  nor (_04343_, _04342_, _03908_);
  not (_04344_, _04343_);
  nor (_04345_, _04344_, _04341_);
  and (_04346_, _03908_, _02934_);
  nor (_04347_, _04346_, _04159_);
  not (_04348_, _04347_);
  nor (_04349_, _04348_, _04345_);
  or (_04350_, _04349_, _03627_);
  nor (_04351_, _04350_, _04251_);
  not (_04352_, _02932_);
  and (_04353_, _03627_, _04352_);
  or (_04354_, _04353_, _03926_);
  nor (_04355_, _04354_, _04351_);
  or (_04356_, _04355_, _03925_);
  nor (_04357_, _04356_, _04243_);
  and (_04358_, _03925_, _02934_);
  nor (_04359_, _04358_, _04357_);
  and (_04360_, _03925_, _03261_);
  and (_04361_, _03216_, _02500_);
  nor (_04362_, _04244_, \oc8051_golden_model_1.SP [2]);
  nor (_04363_, _04362_, _04245_);
  and (_04364_, _04363_, _02531_);
  and (_04365_, _03885_, _03261_);
  nor (_04366_, _02871_, _03261_);
  and (_04367_, _03216_, _02874_);
  and (_04369_, _04363_, _02886_);
  and (_04370_, _03822_, _03261_);
  not (_04372_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_04373_, _03593_, _04372_);
  not (_04375_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_04376_, _03760_, _04375_);
  and (_04378_, _04376_, _03758_);
  nand (_04379_, _04378_, _04373_);
  not (_04381_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_04382_, _03760_, _04381_);
  not (_04384_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04385_, _03593_, _04384_);
  and (_04387_, _04385_, _03766_);
  nand (_04388_, _04387_, _04382_);
  nand (_04390_, _04388_, _04379_);
  nand (_04391_, _04390_, _03374_);
  not (_04393_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_04394_, _03760_, _04393_);
  not (_04396_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04397_, _03593_, _04396_);
  and (_04399_, _04397_, _03766_);
  nand (_04400_, _04399_, _04394_);
  not (_04402_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04403_, _03593_, _04402_);
  not (_04405_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_04406_, _03760_, _04405_);
  and (_04407_, _04406_, _03758_);
  nand (_04408_, _04407_, _04403_);
  nand (_04409_, _04408_, _04400_);
  nand (_04410_, _04409_, _03773_);
  nand (_04411_, _04410_, _04391_);
  nand (_04412_, _04411_, _03181_);
  not (_04413_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_04414_, _03760_, _04413_);
  not (_04415_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04416_, _03593_, _04415_);
  and (_04417_, _04416_, _03766_);
  nand (_04418_, _04417_, _04414_);
  nand (_04419_, _03760_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_04420_, _03593_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04421_, _04420_, _03758_);
  nand (_04422_, _04421_, _04419_);
  nand (_04423_, _04422_, _04418_);
  nand (_04424_, _04423_, _03374_);
  not (_04425_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_04426_, _03760_, _04425_);
  not (_04427_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04428_, _03593_, _04427_);
  and (_04429_, _04428_, _03766_);
  nand (_04430_, _04429_, _04426_);
  nand (_04431_, _03760_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_04432_, _03593_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_04433_, _04432_, _03758_);
  nand (_04435_, _04433_, _04431_);
  nand (_04436_, _04435_, _04430_);
  nand (_04437_, _04436_, _03773_);
  nand (_04438_, _04437_, _04424_);
  nand (_04439_, _04438_, _03790_);
  nand (_04440_, _04439_, _04412_);
  not (_04441_, _04440_);
  or (_04442_, _04441_, _03819_);
  nor (_04443_, _04151_, _03827_);
  and (_04444_, _03827_, _03261_);
  or (_04445_, _04444_, _03824_);
  or (_04446_, _04445_, _04443_);
  nor (_04447_, _04363_, _02558_);
  not (_04448_, _04447_);
  nor (_04449_, _04114_, _04140_);
  and (_04450_, _04449_, _04448_);
  and (_04451_, _04450_, _04446_);
  and (_04452_, _04451_, _03823_);
  and (_04453_, _04452_, _04442_);
  nor (_04454_, _04453_, _04370_);
  nor (_04455_, _04454_, _02894_);
  nor (_04456_, _04455_, _03217_);
  nor (_04457_, _04363_, _02556_);
  nor (_04458_, _04457_, _04456_);
  and (_04459_, _03845_, _03260_);
  and (_04460_, _02842_, _02885_);
  nor (_04461_, _04460_, _04459_);
  and (_04462_, _04461_, _04458_);
  and (_04463_, _04440_, _03413_);
  nor (_04465_, _04463_, _03854_);
  and (_04467_, _04465_, _04462_);
  and (_04468_, _03854_, _03261_);
  nor (_04470_, _04468_, _04467_);
  and (_04471_, _03215_, _03853_);
  nor (_04473_, _04471_, _04470_);
  and (_04474_, _04473_, _03947_);
  nor (_04476_, _04474_, _04369_);
  and (_04477_, _02883_, _03215_);
  or (_04479_, _04477_, _04476_);
  nor (_04480_, _04363_, _02561_);
  nor (_04482_, _04480_, _02981_);
  not (_04483_, _04482_);
  nor (_04485_, _04483_, _04479_);
  and (_04486_, _04440_, _03867_);
  nor (_04488_, _04486_, _03626_);
  and (_04489_, _04488_, _04485_);
  nor (_04491_, _04489_, _04367_);
  nor (_04492_, _04491_, _02578_);
  and (_04494_, _04363_, _02578_);
  nor (_04495_, _04494_, _04492_);
  or (_04497_, _04495_, _04110_);
  nor (_04498_, _04497_, _04366_);
  and (_04499_, _04440_, _03879_);
  nor (_04500_, _04499_, _03885_);
  and (_04501_, _04500_, _04498_);
  nor (_04502_, _04501_, _04365_);
  nor (_04503_, _04502_, _02517_);
  and (_04504_, _04363_, _02517_);
  nor (_04505_, _04504_, _04503_);
  nor (_04506_, _03894_, _03261_);
  nor (_04507_, _04506_, _02533_);
  not (_04508_, _04507_);
  nor (_04509_, _04508_, _04505_);
  and (_04510_, _04363_, _02533_);
  nor (_04511_, _04510_, _04509_);
  and (_04512_, _03901_, _03260_);
  nor (_04513_, _04512_, _02531_);
  not (_04514_, _04513_);
  nor (_04515_, _04514_, _04511_);
  nor (_04516_, _04515_, _04364_);
  not (_04517_, _03711_);
  and (_04518_, _04084_, _04517_);
  not (_04519_, _04518_);
  nor (_04520_, _04519_, _04516_);
  and (_04521_, _04440_, _03909_);
  nor (_04522_, _04521_, _03908_);
  and (_04523_, _04522_, _04520_);
  and (_04524_, _03908_, _03261_);
  nor (_04525_, _04524_, _04523_);
  nor (_04526_, _04363_, _03916_);
  nor (_04527_, _04526_, _03627_);
  not (_04528_, _04527_);
  nor (_04529_, _04528_, _04525_);
  nor (_04530_, _04529_, _04361_);
  nor (_04531_, _04530_, _03580_);
  and (_04532_, _04440_, _03926_);
  nor (_04533_, _04532_, _03925_);
  and (_04534_, _04533_, _04531_);
  nor (_04535_, _04534_, _04360_);
  nor (_04536_, _04535_, _04187_);
  not (_04537_, _04536_);
  nor (_04538_, _04537_, _04359_);
  and (_04539_, _04538_, _04189_);
  or (_04540_, _04539_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04541_, _04247_, _02877_);
  nor (_04542_, _04363_, _03939_);
  nor (_04543_, _04542_, _04541_);
  and (_04544_, _04248_, _02877_);
  nor (_04545_, _04541_, _04250_);
  nor (_04546_, _04545_, _04544_);
  and (_04548_, _35422_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_04549_, _04548_);
  and (_04550_, _04128_, _03916_);
  nor (_04551_, _04550_, _04549_);
  and (_04552_, _04551_, _04546_);
  and (_04553_, _04552_, _04543_);
  and (_04554_, _04553_, _03938_);
  not (_04555_, _04554_);
  and (_04556_, _04555_, _04540_);
  nor (_04557_, _04549_, _04185_);
  not (_04558_, _04557_);
  nor (_04559_, _04558_, _03932_);
  not (_04560_, _04559_);
  nor (_04561_, _04560_, _04103_);
  not (_04562_, _04561_);
  not (_04563_, _04535_);
  nor (_04564_, _04558_, _04359_);
  nand (_04565_, _04564_, _04563_);
  or (_04566_, _04565_, _04562_);
  nand (_04567_, _03760_, \oc8051_golden_model_1.IRAM[0] [7]);
  nand (_04568_, _03593_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_04569_, _04568_, _03758_);
  nand (_04570_, _04569_, _04567_);
  not (_04571_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_04572_, _03760_, _04571_);
  not (_04573_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_04574_, _03593_, _04573_);
  and (_04575_, _04574_, _03766_);
  nand (_04576_, _04575_, _04572_);
  nand (_04577_, _04576_, _04570_);
  nand (_04578_, _04577_, _03374_);
  not (_04579_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_04580_, _03760_, _04579_);
  not (_04581_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04582_, _03593_, _04581_);
  and (_04583_, _04582_, _03766_);
  nand (_04584_, _04583_, _04580_);
  nand (_04585_, _03760_, \oc8051_golden_model_1.IRAM[4] [7]);
  nand (_04586_, _03593_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_04587_, _04586_, _03758_);
  nand (_04588_, _04587_, _04585_);
  nand (_04589_, _04588_, _04584_);
  nand (_04590_, _04589_, _03773_);
  nand (_04591_, _04590_, _04578_);
  nand (_04592_, _04591_, _03181_);
  not (_04593_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_04594_, _03760_, _04593_);
  not (_04595_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04596_, _03593_, _04595_);
  and (_04597_, _04596_, _03766_);
  nand (_04598_, _04597_, _04594_);
  not (_04599_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_04600_, _03593_, _04599_);
  not (_04601_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_04602_, _03760_, _04601_);
  and (_04603_, _04602_, _03758_);
  nand (_04604_, _04603_, _04600_);
  nand (_04605_, _04604_, _04598_);
  nand (_04606_, _04605_, _03374_);
  not (_04607_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_04608_, _03760_, _04607_);
  not (_04609_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04610_, _03593_, _04609_);
  and (_04611_, _04610_, _03766_);
  nand (_04612_, _04611_, _04608_);
  not (_04613_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_04614_, _03593_, _04613_);
  not (_04615_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_04616_, _03760_, _04615_);
  and (_04617_, _04616_, _03758_);
  nand (_04618_, _04617_, _04614_);
  nand (_04619_, _04618_, _04612_);
  nand (_04620_, _04619_, _03773_);
  nand (_04621_, _04620_, _04606_);
  nand (_04622_, _04621_, _03790_);
  nand (_04623_, _04622_, _04592_);
  nor (_04624_, _04623_, _02768_);
  not (_04625_, _04624_);
  and (_04626_, _02932_, _02768_);
  and (_04627_, _04626_, _03215_);
  and (_04628_, _04627_, _03625_);
  and (_04629_, _04628_, _02799_);
  nor (_04630_, _03671_, _02832_);
  and (_04631_, _04630_, _03260_);
  and (_04632_, _04631_, _04629_);
  and (_04633_, _04632_, \oc8051_golden_model_1.DPH [7]);
  not (_04634_, _04633_);
  and (_04635_, _03671_, _02832_);
  nor (_04636_, _03260_, _02799_);
  and (_04637_, _04636_, _04635_);
  and (_04638_, _04637_, _04628_);
  and (_04639_, _04638_, \oc8051_golden_model_1.TH0 [7]);
  not (_04640_, _04630_);
  nand (_04641_, _03260_, _02934_);
  nor (_04642_, _04641_, _04640_);
  and (_04643_, _04642_, _04628_);
  and (_04644_, _04643_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04645_, _04644_, _04639_);
  and (_04646_, _04645_, _04634_);
  and (_04647_, _03671_, _02833_);
  and (_04649_, _04647_, _03260_);
  and (_04650_, _04649_, _04629_);
  and (_04651_, _04650_, \oc8051_golden_model_1.SP [7]);
  nor (_04652_, _03671_, _02833_);
  and (_04653_, _04652_, _03260_);
  and (_04654_, _04653_, _04629_);
  and (_04655_, _04654_, \oc8051_golden_model_1.DPL [7]);
  nor (_04656_, _04655_, _04651_);
  and (_04657_, _04630_, _03261_);
  and (_04658_, _04657_, _04629_);
  and (_04659_, _04658_, \oc8051_golden_model_1.PCON [7]);
  not (_04660_, _04659_);
  and (_04661_, _04649_, _02934_);
  not (_04662_, _03625_);
  and (_04663_, _04662_, _03215_);
  and (_04664_, _04663_, _04626_);
  and (_04665_, _04664_, _04661_);
  and (_04666_, _04665_, \oc8051_golden_model_1.SBUF [7]);
  and (_04667_, _04635_, _03260_);
  and (_04668_, _04667_, _02934_);
  not (_04669_, _03215_);
  and (_04670_, _03625_, _04669_);
  and (_04671_, _04670_, _04626_);
  and (_04672_, _04671_, _04668_);
  and (_04673_, _04672_, \oc8051_golden_model_1.IE [7]);
  nor (_04674_, _04673_, _04666_);
  and (_04675_, _04674_, _04660_);
  and (_04676_, _04675_, _04656_);
  and (_04677_, _04676_, _04646_);
  not (_04678_, _04628_);
  not (_04679_, _04652_);
  or (_04680_, _04679_, _04641_);
  nor (_04681_, _04680_, _04678_);
  and (_04682_, _04681_, \oc8051_golden_model_1.TL0 [7]);
  and (_04683_, _04668_, _04664_);
  and (_04684_, _04683_, \oc8051_golden_model_1.SCON [7]);
  nor (_04685_, _04684_, _04682_);
  and (_04686_, _04647_, _04636_);
  and (_04687_, _04686_, _04628_);
  and (_04688_, _04687_, \oc8051_golden_model_1.TH1 [7]);
  not (_04689_, _04688_);
  and (_04690_, _04668_, _04628_);
  and (_04691_, _04690_, \oc8051_golden_model_1.TCON [7]);
  and (_04692_, _04661_, _04628_);
  and (_04693_, _04692_, \oc8051_golden_model_1.TMOD [7]);
  nor (_04694_, _04693_, _04691_);
  and (_04695_, _04694_, _04689_);
  and (_04696_, _04695_, _04685_);
  nor (_04697_, _03625_, _03215_);
  and (_04698_, _04697_, _04626_);
  and (_04699_, _04698_, _04668_);
  and (_04700_, _04699_, \oc8051_golden_model_1.IP [7]);
  and (_04701_, _03260_, _02799_);
  and (_04702_, _04701_, _04635_);
  nor (_04703_, _02932_, _02858_);
  and (_04704_, _04703_, _04697_);
  and (_04705_, _04704_, _04702_);
  and (_04706_, _04705_, \oc8051_golden_model_1.B [7]);
  nor (_04707_, _04706_, _04700_);
  and (_04708_, _04703_, _04663_);
  and (_04709_, _04708_, _04702_);
  and (_04710_, _04709_, \oc8051_golden_model_1.PSW [7]);
  and (_04711_, _04703_, _04670_);
  and (_04712_, _04711_, _04702_);
  and (_04713_, _04712_, \oc8051_golden_model_1.ACC [7]);
  nor (_04714_, _04713_, _04710_);
  and (_04715_, _04714_, _04707_);
  and (_04716_, _04702_, _04628_);
  and (_04717_, _04716_, \oc8051_golden_model_1.P0 [7]);
  not (_04718_, _04717_);
  and (_04719_, _04702_, _04664_);
  and (_04720_, _04719_, \oc8051_golden_model_1.P1 [7]);
  not (_04721_, _04720_);
  and (_04722_, _04702_, _04671_);
  and (_04723_, _04722_, \oc8051_golden_model_1.P2 [7]);
  and (_04724_, _04702_, _04698_);
  and (_04725_, _04724_, \oc8051_golden_model_1.P3 [7]);
  nor (_04726_, _04725_, _04723_);
  and (_04727_, _04726_, _04721_);
  and (_04728_, _04727_, _04718_);
  and (_04729_, _04728_, _04715_);
  and (_04730_, _04729_, _04696_);
  and (_04731_, _04730_, _04677_);
  and (_04732_, _04731_, _04625_);
  not (_04733_, _04732_);
  not (_04734_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_04735_, _03593_, _04734_);
  not (_04736_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_04737_, _03760_, _04736_);
  and (_04738_, _04737_, _03758_);
  nand (_04739_, _04738_, _04735_);
  not (_04740_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_04741_, _03760_, _04740_);
  not (_04742_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_04743_, _03593_, _04742_);
  and (_04744_, _04743_, _03766_);
  nand (_04745_, _04744_, _04741_);
  nand (_04746_, _04745_, _04739_);
  nand (_04747_, _04746_, _03374_);
  not (_04748_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_04750_, _03760_, _04748_);
  not (_04751_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_04752_, _03593_, _04751_);
  and (_04753_, _04752_, _03766_);
  nand (_04754_, _04753_, _04750_);
  not (_04755_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04756_, _03593_, _04755_);
  not (_04757_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_04758_, _03760_, _04757_);
  and (_04759_, _04758_, _03758_);
  nand (_04760_, _04759_, _04756_);
  nand (_04761_, _04760_, _04754_);
  nand (_04762_, _04761_, _03773_);
  nand (_04763_, _04762_, _04747_);
  nand (_04764_, _04763_, _03181_);
  nand (_04765_, _03593_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04766_, _03760_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04767_, _04766_, _03766_);
  nand (_04768_, _04767_, _04765_);
  nand (_04769_, _03760_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04770_, _03593_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04771_, _04770_, _03758_);
  nand (_04772_, _04771_, _04769_);
  nand (_04773_, _04772_, _04768_);
  nand (_04774_, _04773_, _03374_);
  nand (_04775_, _03593_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04776_, _03760_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04777_, _04776_, _03766_);
  nand (_04778_, _04777_, _04775_);
  nand (_04779_, _03760_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_04780_, _03593_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_04781_, _04780_, _03758_);
  nand (_04782_, _04781_, _04779_);
  nand (_04783_, _04782_, _04778_);
  nand (_04784_, _04783_, _03773_);
  nand (_04785_, _04784_, _04774_);
  nand (_04786_, _04785_, _03790_);
  nand (_04787_, _04786_, _04764_);
  or (_04788_, _04787_, _02768_);
  and (_04789_, _04650_, \oc8051_golden_model_1.SP [6]);
  not (_04790_, _04789_);
  and (_04791_, _04654_, \oc8051_golden_model_1.DPL [6]);
  and (_04792_, _04690_, \oc8051_golden_model_1.TCON [6]);
  nor (_04793_, _04792_, _04791_);
  and (_04794_, _04793_, _04790_);
  and (_04795_, _04716_, \oc8051_golden_model_1.P0 [6]);
  not (_04796_, _04795_);
  and (_04797_, _04719_, \oc8051_golden_model_1.P1 [6]);
  not (_04798_, _04797_);
  and (_04799_, _04722_, \oc8051_golden_model_1.P2 [6]);
  and (_04800_, _04724_, \oc8051_golden_model_1.P3 [6]);
  nor (_04801_, _04800_, _04799_);
  and (_04802_, _04801_, _04798_);
  and (_04803_, _04802_, _04796_);
  and (_04804_, _04803_, _04794_);
  and (_04805_, _04692_, \oc8051_golden_model_1.TMOD [6]);
  and (_04806_, _04687_, \oc8051_golden_model_1.TH1 [6]);
  nor (_04807_, _04806_, _04805_);
  and (_04808_, _04681_, \oc8051_golden_model_1.TL0 [6]);
  and (_04809_, _04643_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04810_, _04809_, _04808_);
  and (_04811_, _04810_, _04807_);
  and (_04812_, _04632_, \oc8051_golden_model_1.DPH [6]);
  not (_04813_, _04812_);
  and (_04814_, _04638_, \oc8051_golden_model_1.TH0 [6]);
  and (_04815_, _04683_, \oc8051_golden_model_1.SCON [6]);
  nor (_04816_, _04815_, _04814_);
  and (_04817_, _04816_, _04813_);
  and (_04818_, _04817_, _04811_);
  and (_04819_, _04658_, \oc8051_golden_model_1.PCON [6]);
  not (_04820_, _04819_);
  and (_04821_, _04709_, \oc8051_golden_model_1.PSW [6]);
  not (_04822_, _04821_);
  and (_04823_, _04699_, \oc8051_golden_model_1.IP [6]);
  and (_04824_, _04705_, \oc8051_golden_model_1.B [6]);
  nor (_04825_, _04824_, _04823_);
  and (_04826_, _04825_, _04822_);
  and (_04827_, _04665_, \oc8051_golden_model_1.SBUF [6]);
  not (_04828_, _04827_);
  and (_04829_, _04672_, \oc8051_golden_model_1.IE [6]);
  and (_04830_, _04712_, \oc8051_golden_model_1.ACC [6]);
  nor (_04831_, _04830_, _04829_);
  and (_04832_, _04831_, _04828_);
  and (_04833_, _04832_, _04826_);
  and (_04834_, _04833_, _04820_);
  and (_04835_, _04834_, _04818_);
  and (_04836_, _04835_, _04804_);
  and (_04837_, _04836_, _04788_);
  not (_04838_, _04837_);
  not (_04839_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_04840_, _03593_, _04839_);
  not (_04841_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_04842_, _03760_, _04841_);
  and (_04843_, _04842_, _03758_);
  nand (_04844_, _04843_, _04840_);
  not (_04845_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_04846_, _03760_, _04845_);
  not (_04847_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_04848_, _03593_, _04847_);
  and (_04849_, _04848_, _03766_);
  nand (_04851_, _04849_, _04846_);
  nand (_04852_, _04851_, _04844_);
  nand (_04853_, _04852_, _03374_);
  not (_04854_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_04855_, _03760_, _04854_);
  not (_04856_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_04857_, _03593_, _04856_);
  and (_04858_, _04857_, _03766_);
  nand (_04859_, _04858_, _04855_);
  not (_04860_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_04861_, _03593_, _04860_);
  not (_04862_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_04863_, _03760_, _04862_);
  and (_04864_, _04863_, _03758_);
  nand (_04865_, _04864_, _04861_);
  nand (_04866_, _04865_, _04859_);
  nand (_04867_, _04866_, _03773_);
  nand (_04868_, _04867_, _04853_);
  nand (_04869_, _04868_, _03181_);
  nand (_04870_, _03593_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_04871_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_04872_, _03593_, _04871_);
  and (_04873_, _04872_, _03766_);
  nand (_04874_, _04873_, _04870_);
  nand (_04875_, _03760_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_04876_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_04877_, _03760_, _04876_);
  and (_04878_, _04877_, _03758_);
  nand (_04879_, _04878_, _04875_);
  nand (_04880_, _04879_, _04874_);
  nand (_04881_, _04880_, _03374_);
  nand (_04882_, _03593_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_04883_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_04884_, _03593_, _04883_);
  and (_04885_, _04884_, _03766_);
  nand (_04886_, _04885_, _04882_);
  nand (_04887_, _03760_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_04888_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_04889_, _03760_, _04888_);
  and (_04890_, _04889_, _03758_);
  nand (_04891_, _04890_, _04887_);
  nand (_04892_, _04891_, _04886_);
  nand (_04893_, _04892_, _03773_);
  nand (_04894_, _04893_, _04881_);
  nand (_04895_, _04894_, _03790_);
  nand (_04896_, _04895_, _04869_);
  or (_04897_, _04896_, _02768_);
  and (_04898_, _04650_, \oc8051_golden_model_1.SP [5]);
  and (_04899_, _04654_, \oc8051_golden_model_1.DPL [5]);
  nor (_04900_, _04899_, _04898_);
  nand (_04901_, _04632_, \oc8051_golden_model_1.DPH [5]);
  and (_04902_, _04901_, _04900_);
  and (_04903_, _04690_, \oc8051_golden_model_1.TCON [5]);
  not (_04904_, _04903_);
  and (_04905_, _04681_, \oc8051_golden_model_1.TL0 [5]);
  and (_04906_, _04683_, \oc8051_golden_model_1.SCON [5]);
  nor (_04907_, _04906_, _04905_);
  and (_04908_, _04907_, _04904_);
  and (_04909_, _04638_, \oc8051_golden_model_1.TH0 [5]);
  and (_04910_, _04687_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04911_, _04910_, _04909_);
  and (_04912_, _04692_, \oc8051_golden_model_1.TMOD [5]);
  and (_04913_, _04643_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04914_, _04913_, _04912_);
  and (_04915_, _04914_, _04911_);
  and (_04916_, _04915_, _04908_);
  and (_04917_, _04916_, _04902_);
  and (_04918_, _04658_, \oc8051_golden_model_1.PCON [5]);
  not (_04919_, _04918_);
  and (_04920_, _04665_, \oc8051_golden_model_1.SBUF [5]);
  and (_04921_, _04672_, \oc8051_golden_model_1.IE [5]);
  nor (_04922_, _04921_, _04920_);
  and (_04923_, _04922_, _04919_);
  and (_04924_, _04716_, \oc8051_golden_model_1.P0 [5]);
  not (_04925_, _04924_);
  and (_04926_, _04709_, \oc8051_golden_model_1.PSW [5]);
  and (_04927_, _04712_, \oc8051_golden_model_1.ACC [5]);
  nor (_04928_, _04927_, _04926_);
  and (_04929_, _04699_, \oc8051_golden_model_1.IP [5]);
  and (_04930_, _04705_, \oc8051_golden_model_1.B [5]);
  nor (_04931_, _04930_, _04929_);
  and (_04932_, _04931_, _04928_);
  and (_04933_, _04719_, \oc8051_golden_model_1.P1 [5]);
  not (_04934_, _04933_);
  and (_04935_, _04722_, \oc8051_golden_model_1.P2 [5]);
  and (_04936_, _04724_, \oc8051_golden_model_1.P3 [5]);
  nor (_04937_, _04936_, _04935_);
  and (_04938_, _04937_, _04934_);
  and (_04939_, _04938_, _04932_);
  and (_04940_, _04939_, _04925_);
  and (_04941_, _04940_, _04923_);
  and (_04942_, _04941_, _04917_);
  and (_04943_, _04942_, _04897_);
  not (_04944_, _04943_);
  or (_04945_, _04242_, _02768_);
  and (_04946_, _04654_, \oc8051_golden_model_1.DPL [3]);
  not (_04947_, _04946_);
  and (_04948_, _04650_, \oc8051_golden_model_1.SP [3]);
  and (_04949_, _04690_, \oc8051_golden_model_1.TCON [3]);
  nor (_04950_, _04949_, _04948_);
  and (_04952_, _04950_, _04947_);
  and (_04953_, _04716_, \oc8051_golden_model_1.P0 [3]);
  not (_04954_, _04953_);
  and (_04955_, _04719_, \oc8051_golden_model_1.P1 [3]);
  not (_04956_, _04955_);
  and (_04957_, _04722_, \oc8051_golden_model_1.P2 [3]);
  and (_04958_, _04724_, \oc8051_golden_model_1.P3 [3]);
  nor (_04959_, _04958_, _04957_);
  and (_04960_, _04959_, _04956_);
  and (_04961_, _04960_, _04954_);
  and (_04962_, _04961_, _04952_);
  and (_04963_, _04643_, \oc8051_golden_model_1.TL1 [3]);
  and (_04964_, _04687_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04692_, \oc8051_golden_model_1.TMOD [3]);
  and (_04967_, _04683_, \oc8051_golden_model_1.SCON [3]);
  nor (_04968_, _04967_, _04966_);
  and (_04969_, _04968_, _04965_);
  and (_04970_, _04632_, \oc8051_golden_model_1.DPH [3]);
  not (_04971_, _04970_);
  and (_04972_, _04681_, \oc8051_golden_model_1.TL0 [3]);
  and (_04973_, _04638_, \oc8051_golden_model_1.TH0 [3]);
  nor (_04974_, _04973_, _04972_);
  and (_04975_, _04974_, _04971_);
  and (_04976_, _04975_, _04969_);
  and (_04977_, _04658_, \oc8051_golden_model_1.PCON [3]);
  not (_04978_, _04977_);
  and (_04979_, _04699_, \oc8051_golden_model_1.IP [3]);
  not (_04980_, _04979_);
  and (_04981_, _04709_, \oc8051_golden_model_1.PSW [3]);
  and (_04982_, _04705_, \oc8051_golden_model_1.B [3]);
  nor (_04983_, _04982_, _04981_);
  and (_04984_, _04983_, _04980_);
  and (_04985_, _04665_, \oc8051_golden_model_1.SBUF [3]);
  not (_04986_, _04985_);
  and (_04987_, _04672_, \oc8051_golden_model_1.IE [3]);
  and (_04988_, _04712_, \oc8051_golden_model_1.ACC [3]);
  nor (_04989_, _04988_, _04987_);
  and (_04990_, _04989_, _04986_);
  and (_04991_, _04990_, _04984_);
  and (_04992_, _04991_, _04978_);
  and (_04993_, _04992_, _04976_);
  and (_04994_, _04993_, _04962_);
  and (_04995_, _04994_, _04945_);
  not (_04996_, _04995_);
  nand (_04997_, _03817_, _02858_);
  and (_04998_, _04658_, \oc8051_golden_model_1.PCON [0]);
  not (_04999_, _04998_);
  and (_05000_, _04665_, \oc8051_golden_model_1.SBUF [0]);
  and (_05001_, _04672_, \oc8051_golden_model_1.IE [0]);
  nor (_05002_, _05001_, _05000_);
  and (_05003_, _05002_, _04999_);
  and (_05004_, _04722_, \oc8051_golden_model_1.P2 [0]);
  and (_05005_, _04724_, \oc8051_golden_model_1.P3 [0]);
  nor (_05006_, _05005_, _05004_);
  and (_05007_, _05006_, _05003_);
  and (_05008_, _04699_, \oc8051_golden_model_1.IP [0]);
  and (_05009_, _04705_, \oc8051_golden_model_1.B [0]);
  nor (_05010_, _05009_, _05008_);
  and (_05011_, _04709_, \oc8051_golden_model_1.PSW [0]);
  and (_05012_, _04712_, \oc8051_golden_model_1.ACC [0]);
  nor (_05013_, _05012_, _05011_);
  and (_05014_, _05013_, _05010_);
  and (_05015_, _04690_, \oc8051_golden_model_1.TCON [0]);
  and (_05016_, _04638_, \oc8051_golden_model_1.TH0 [0]);
  nor (_05017_, _05016_, _05015_);
  and (_05018_, _04719_, \oc8051_golden_model_1.P1 [0]);
  and (_05019_, _04643_, \oc8051_golden_model_1.TL1 [0]);
  nor (_05020_, _05019_, _05018_);
  and (_05021_, _05020_, _05017_);
  and (_05022_, _04683_, \oc8051_golden_model_1.SCON [0]);
  and (_05023_, _04687_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05024_, _05023_, _05022_);
  and (_05025_, _04681_, \oc8051_golden_model_1.TL0 [0]);
  and (_05026_, _04692_, \oc8051_golden_model_1.TMOD [0]);
  nor (_05027_, _05026_, _05025_);
  and (_05028_, _05027_, _05024_);
  and (_05029_, _05028_, _05021_);
  and (_05030_, _05029_, _05014_);
  and (_05031_, _05030_, _05007_);
  and (_05032_, _04716_, \oc8051_golden_model_1.P0 [0]);
  not (_05033_, _05032_);
  and (_05034_, _04650_, \oc8051_golden_model_1.SP [0]);
  and (_05035_, _04654_, \oc8051_golden_model_1.DPL [0]);
  nor (_05036_, _05035_, _05034_);
  and (_05037_, _04701_, _04630_);
  and (_05038_, _05037_, _04628_);
  and (_05039_, _05038_, \oc8051_golden_model_1.DPH [0]);
  not (_05040_, _05039_);
  and (_05041_, _05040_, _05036_);
  and (_05042_, _05041_, _05033_);
  and (_05043_, _05042_, _05031_);
  and (_05044_, _05043_, _04997_);
  or (_05045_, _04038_, _02768_);
  and (_05046_, _04654_, \oc8051_golden_model_1.DPL [1]);
  not (_05047_, _05046_);
  and (_05048_, _04650_, \oc8051_golden_model_1.SP [1]);
  and (_05049_, _04690_, \oc8051_golden_model_1.TCON [1]);
  nor (_05050_, _05049_, _05048_);
  and (_05051_, _05050_, _05047_);
  and (_05053_, _04716_, \oc8051_golden_model_1.P0 [1]);
  not (_05054_, _05053_);
  and (_05055_, _04719_, \oc8051_golden_model_1.P1 [1]);
  not (_05056_, _05055_);
  and (_05057_, _04722_, \oc8051_golden_model_1.P2 [1]);
  and (_05058_, _04724_, \oc8051_golden_model_1.P3 [1]);
  nor (_05059_, _05058_, _05057_);
  and (_05060_, _05059_, _05056_);
  and (_05061_, _05060_, _05054_);
  and (_05062_, _05061_, _05051_);
  and (_05063_, _04692_, \oc8051_golden_model_1.TMOD [1]);
  and (_05064_, _04687_, \oc8051_golden_model_1.TH1 [1]);
  nor (_05065_, _05064_, _05063_);
  and (_05066_, _04681_, \oc8051_golden_model_1.TL0 [1]);
  and (_05067_, _04643_, \oc8051_golden_model_1.TL1 [1]);
  nor (_05068_, _05067_, _05066_);
  and (_05069_, _05068_, _05065_);
  and (_05070_, _04632_, \oc8051_golden_model_1.DPH [1]);
  not (_05071_, _05070_);
  and (_05072_, _04638_, \oc8051_golden_model_1.TH0 [1]);
  and (_05073_, _04683_, \oc8051_golden_model_1.SCON [1]);
  nor (_05074_, _05073_, _05072_);
  and (_05075_, _05074_, _05071_);
  and (_05076_, _05075_, _05069_);
  and (_05077_, _04658_, \oc8051_golden_model_1.PCON [1]);
  not (_05078_, _05077_);
  and (_05079_, _04709_, \oc8051_golden_model_1.PSW [1]);
  not (_05080_, _05079_);
  and (_05081_, _04699_, \oc8051_golden_model_1.IP [1]);
  and (_05082_, _04705_, \oc8051_golden_model_1.B [1]);
  nor (_05083_, _05082_, _05081_);
  and (_05084_, _05083_, _05080_);
  and (_05085_, _04665_, \oc8051_golden_model_1.SBUF [1]);
  not (_05086_, _05085_);
  and (_05087_, _04672_, \oc8051_golden_model_1.IE [1]);
  and (_05088_, _04712_, \oc8051_golden_model_1.ACC [1]);
  nor (_05089_, _05088_, _05087_);
  and (_05090_, _05089_, _05086_);
  and (_05091_, _05090_, _05084_);
  and (_05092_, _05091_, _05078_);
  and (_05093_, _05092_, _05076_);
  and (_05094_, _05093_, _05062_);
  and (_05095_, _05094_, _05045_);
  nor (_05096_, _05095_, _05044_);
  or (_05097_, _04440_, _02768_);
  and (_05098_, _04658_, \oc8051_golden_model_1.PCON [2]);
  not (_05099_, _05098_);
  and (_05100_, _04665_, \oc8051_golden_model_1.SBUF [2]);
  and (_05101_, _04672_, \oc8051_golden_model_1.IE [2]);
  nor (_05102_, _05101_, _05100_);
  and (_05103_, _05102_, _05099_);
  and (_05104_, _04722_, \oc8051_golden_model_1.P2 [2]);
  and (_05105_, _04724_, \oc8051_golden_model_1.P3 [2]);
  nor (_05106_, _05105_, _05104_);
  and (_05107_, _05106_, _05103_);
  and (_05108_, _04699_, \oc8051_golden_model_1.IP [2]);
  and (_05109_, _04712_, \oc8051_golden_model_1.ACC [2]);
  nor (_05110_, _05109_, _05108_);
  and (_05111_, _04709_, \oc8051_golden_model_1.PSW [2]);
  and (_05112_, _04705_, \oc8051_golden_model_1.B [2]);
  nor (_05113_, _05112_, _05111_);
  and (_05114_, _05113_, _05110_);
  and (_05115_, _04690_, \oc8051_golden_model_1.TCON [2]);
  and (_05116_, _04638_, \oc8051_golden_model_1.TH0 [2]);
  nor (_05117_, _05116_, _05115_);
  and (_05118_, _04719_, \oc8051_golden_model_1.P1 [2]);
  and (_05119_, _04643_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05120_, _05119_, _05118_);
  and (_05121_, _05120_, _05117_);
  and (_05122_, _04683_, \oc8051_golden_model_1.SCON [2]);
  and (_05123_, _04687_, \oc8051_golden_model_1.TH1 [2]);
  nor (_05124_, _05123_, _05122_);
  and (_05125_, _04692_, \oc8051_golden_model_1.TMOD [2]);
  and (_05126_, _04681_, \oc8051_golden_model_1.TL0 [2]);
  nor (_05127_, _05126_, _05125_);
  and (_05128_, _05127_, _05124_);
  and (_05129_, _05128_, _05121_);
  and (_05130_, _05129_, _05114_);
  and (_05131_, _05130_, _05107_);
  and (_05132_, _04716_, \oc8051_golden_model_1.P0 [2]);
  not (_05133_, _05132_);
  and (_05134_, _04650_, \oc8051_golden_model_1.SP [2]);
  and (_05135_, _04654_, \oc8051_golden_model_1.DPL [2]);
  nor (_05136_, _05135_, _05134_);
  and (_05137_, _05038_, \oc8051_golden_model_1.DPH [2]);
  not (_05138_, _05137_);
  and (_05139_, _05138_, _05136_);
  and (_05140_, _05139_, _05133_);
  and (_05141_, _05140_, _05131_);
  and (_05142_, _05141_, _05097_);
  not (_05143_, _05142_);
  and (_05144_, _05143_, _05096_);
  and (_05145_, _05144_, _04996_);
  not (_05146_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_05147_, _03593_, _05146_);
  not (_05148_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05149_, _03760_, _05148_);
  and (_05150_, _05149_, _03758_);
  nand (_05151_, _05150_, _05147_);
  not (_05152_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_05153_, _03760_, _05152_);
  not (_05154_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05155_, _03593_, _05154_);
  and (_05156_, _05155_, _03766_);
  nand (_05157_, _05156_, _05153_);
  nand (_05158_, _05157_, _05151_);
  nand (_05159_, _05158_, _03374_);
  not (_05160_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05161_, _03760_, _05160_);
  not (_05162_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05163_, _03593_, _05162_);
  and (_05164_, _05163_, _03766_);
  nand (_05165_, _05164_, _05161_);
  not (_05166_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05167_, _03593_, _05166_);
  not (_05168_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05169_, _03760_, _05168_);
  and (_05170_, _05169_, _03758_);
  nand (_05171_, _05170_, _05167_);
  nand (_05172_, _05171_, _05165_);
  nand (_05173_, _05172_, _03773_);
  nand (_05174_, _05173_, _05159_);
  nand (_05175_, _05174_, _03181_);
  nand (_05176_, _03593_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_05177_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05178_, _03593_, _05177_);
  and (_05179_, _05178_, _03766_);
  nand (_05180_, _05179_, _05176_);
  nand (_05181_, _03760_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_05182_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05183_, _03760_, _05182_);
  and (_05184_, _05183_, _03758_);
  nand (_05185_, _05184_, _05181_);
  nand (_05186_, _05185_, _05180_);
  nand (_05187_, _05186_, _03374_);
  nand (_05188_, _03593_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_05189_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05190_, _03593_, _05189_);
  and (_05191_, _05190_, _03766_);
  nand (_05192_, _05191_, _05188_);
  nand (_05193_, _03760_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_05194_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05195_, _03760_, _05194_);
  and (_05196_, _05195_, _03758_);
  nand (_05197_, _05196_, _05193_);
  nand (_05198_, _05197_, _05192_);
  nand (_05199_, _05198_, _03773_);
  nand (_05200_, _05199_, _05187_);
  nand (_05201_, _05200_, _03790_);
  nand (_05202_, _05201_, _05175_);
  or (_05203_, _05202_, _02768_);
  and (_05204_, _04638_, \oc8051_golden_model_1.TH0 [4]);
  and (_05205_, _04665_, \oc8051_golden_model_1.SBUF [4]);
  nor (_05206_, _05205_, _05204_);
  and (_05207_, _04692_, \oc8051_golden_model_1.TMOD [4]);
  and (_05208_, _04683_, \oc8051_golden_model_1.SCON [4]);
  nor (_05209_, _05208_, _05207_);
  and (_05210_, _05209_, _05206_);
  and (_05211_, _04632_, \oc8051_golden_model_1.DPH [4]);
  not (_05212_, _05211_);
  and (_05213_, _04681_, \oc8051_golden_model_1.TL0 [4]);
  and (_05214_, _04672_, \oc8051_golden_model_1.IE [4]);
  nor (_05215_, _05214_, _05213_);
  and (_05216_, _04643_, \oc8051_golden_model_1.TL1 [4]);
  and (_05217_, _04687_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05218_, _05217_, _05216_);
  and (_05219_, _05218_, _05215_);
  and (_05220_, _05219_, _05212_);
  and (_05221_, _05220_, _05210_);
  and (_05222_, _04716_, \oc8051_golden_model_1.P0 [4]);
  not (_05223_, _05222_);
  and (_05224_, _04658_, \oc8051_golden_model_1.PCON [4]);
  not (_05225_, _05224_);
  and (_05226_, _04709_, \oc8051_golden_model_1.PSW [4]);
  and (_05227_, _04705_, \oc8051_golden_model_1.B [4]);
  nor (_05228_, _05227_, _05226_);
  and (_05229_, _04699_, \oc8051_golden_model_1.IP [4]);
  and (_05230_, _04712_, \oc8051_golden_model_1.ACC [4]);
  nor (_05231_, _05230_, _05229_);
  and (_05232_, _05231_, _05228_);
  and (_05233_, _05232_, _05225_);
  and (_05234_, _05233_, _05223_);
  and (_05235_, _04650_, \oc8051_golden_model_1.SP [4]);
  and (_05236_, _04654_, \oc8051_golden_model_1.DPL [4]);
  nor (_05237_, _05236_, _05235_);
  and (_05238_, _04719_, \oc8051_golden_model_1.P1 [4]);
  not (_05239_, _05238_);
  and (_05240_, _04690_, \oc8051_golden_model_1.TCON [4]);
  not (_05241_, _05240_);
  and (_05242_, _04722_, \oc8051_golden_model_1.P2 [4]);
  and (_05243_, _04724_, \oc8051_golden_model_1.P3 [4]);
  nor (_05244_, _05243_, _05242_);
  and (_05245_, _05244_, _05241_);
  and (_05246_, _05245_, _05239_);
  and (_05247_, _05246_, _05237_);
  and (_05248_, _05247_, _05234_);
  and (_05249_, _05248_, _05221_);
  and (_05250_, _05249_, _05203_);
  not (_05251_, _05250_);
  and (_05252_, _05251_, _05145_);
  and (_05253_, _05252_, _04944_);
  and (_05254_, _05253_, _04838_);
  nor (_05255_, _05254_, _04733_);
  and (_05256_, _05254_, _04733_);
  nor (_05257_, _05256_, _05255_);
  and (_05258_, _05257_, _03925_);
  not (_05259_, _04623_);
  and (_05260_, _05202_, _04896_);
  nor (_05261_, _04005_, _03817_);
  and (_05262_, _04440_, _04242_);
  and (_05263_, _05262_, _05261_);
  and (_05264_, _05263_, _05260_);
  and (_05265_, _05264_, _04787_);
  or (_05266_, _05265_, _05259_);
  nand (_05267_, _05265_, _05259_);
  and (_05268_, _05267_, _05266_);
  and (_05269_, _02834_, _02370_);
  nor (_05270_, _03711_, _05269_);
  and (_05271_, _05270_, _04084_);
  or (_05272_, _05271_, _05268_);
  not (_05273_, _03891_);
  not (_05274_, _03020_);
  nor (_05275_, _05274_, _02768_);
  not (_05276_, _05275_);
  nor (_05277_, _03131_, _02768_);
  not (_05278_, _05277_);
  not (_05279_, _03021_);
  nor (_05280_, _05279_, _02768_);
  and (_05281_, _03096_, _01085_);
  and (_05282_, _03094_, _01157_);
  nor (_05283_, _05282_, _05281_);
  and (_05284_, _03083_, _01170_);
  and (_05285_, _03063_, _01140_);
  nor (_05286_, _05285_, _05284_);
  and (_05287_, _05286_, _05283_);
  and (_05288_, _03112_, _01137_);
  and (_05289_, _03102_, _01119_);
  nor (_05290_, _05289_, _05288_);
  and (_05291_, _03086_, _01125_);
  and (_05292_, _03068_, _01154_);
  nor (_05293_, _05292_, _05291_);
  and (_05294_, _05293_, _05290_);
  and (_05295_, _05294_, _05287_);
  and (_05296_, _03107_, _33937_);
  and (_05297_, _03074_, _01164_);
  nor (_05298_, _05297_, _05296_);
  and (_05299_, _03081_, _01167_);
  and (_05300_, _03114_, _01115_);
  nor (_05301_, _05300_, _05299_);
  and (_05302_, _05301_, _05298_);
  and (_05303_, _03100_, _01161_);
  and (_05304_, _03076_, _01147_);
  nor (_05305_, _05304_, _05303_);
  and (_05306_, _03109_, _01129_);
  and (_05307_, _03088_, _01134_);
  nor (_05308_, _05307_, _05306_);
  and (_05309_, _05308_, _05305_);
  and (_05310_, _05309_, _05302_);
  and (_05311_, _05310_, _05295_);
  and (_05312_, _05311_, _04732_);
  nor (_05313_, _05311_, _04732_);
  nor (_05314_, _05313_, _05312_);
  and (_05315_, _05314_, _05280_);
  and (_05316_, _03029_, _02516_);
  not (_05317_, _05316_);
  or (_05318_, _03017_, _03313_);
  and (_05319_, _05318_, _02516_);
  nor (_05320_, _05319_, _04110_);
  and (_05321_, _05320_, _03880_);
  and (_05322_, _05321_, _05317_);
  and (_05323_, _05322_, _03884_);
  or (_05324_, _05323_, _02768_);
  not (_05325_, _02578_);
  nor (_05326_, _03631_, _03501_);
  and (_05327_, _03219_, _02936_);
  and (_05328_, _05327_, _05326_);
  and (_05329_, _04708_, _05328_);
  and (_05330_, _05329_, \oc8051_golden_model_1.PSW [7]);
  and (_05331_, _04711_, _05328_);
  and (_05332_, _05331_, \oc8051_golden_model_1.ACC [7]);
  nor (_05333_, _05332_, _05330_);
  nor (_05334_, _03216_, _02936_);
  and (_05335_, _05334_, _05326_);
  and (_05336_, _05335_, _04698_);
  and (_05337_, _05336_, \oc8051_golden_model_1.IP [7]);
  and (_05338_, _04704_, _05328_);
  and (_05339_, _05338_, \oc8051_golden_model_1.B [7]);
  nor (_05340_, _05339_, _05337_);
  and (_05341_, _05340_, _05333_);
  and (_05342_, _04629_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05343_, _05342_);
  and (_05344_, _04664_, _05328_);
  and (_05345_, _05344_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05346_, _04671_, _05328_);
  and (_05347_, _05346_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05348_, _05347_, _05345_);
  and (_05349_, _05348_, _05343_);
  and (_05350_, _05335_, _04664_);
  and (_05351_, _05350_, \oc8051_golden_model_1.SCON [7]);
  and (_05352_, _05335_, _04671_);
  and (_05353_, _05352_, \oc8051_golden_model_1.IE [7]);
  nor (_05354_, _05353_, _05351_);
  and (_05355_, _05335_, _04628_);
  and (_05356_, _05355_, \oc8051_golden_model_1.TCON [7]);
  and (_05357_, _04698_, _05328_);
  and (_05358_, _05357_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05359_, _05358_, _05356_);
  and (_05360_, _05359_, _05354_);
  and (_05361_, _05360_, _05349_);
  and (_05362_, _05361_, _05341_);
  and (_05363_, _05362_, _04625_);
  nor (_05364_, _05363_, _04657_);
  and (_05365_, _04657_, \oc8051_golden_model_1.PSW [7]);
  nor (_05366_, _05365_, _05364_);
  nor (_05367_, _05366_, _04303_);
  not (_05368_, _03853_);
  and (_05369_, _05357_, \oc8051_golden_model_1.P3 [7]);
  and (_05370_, _05346_, \oc8051_golden_model_1.P2 [7]);
  or (_05371_, _05370_, _05369_);
  nor (_05372_, _05371_, _05356_);
  and (_05373_, _05344_, \oc8051_golden_model_1.P1 [7]);
  and (_05374_, _04629_, \oc8051_golden_model_1.P0 [7]);
  nor (_05375_, _05374_, _05373_);
  and (_05376_, _05375_, _05354_);
  and (_05377_, _05376_, _05341_);
  and (_05378_, _05377_, _05372_);
  and (_05379_, _05378_, _04625_);
  nor (_05380_, _05379_, _04657_);
  or (_05381_, _05380_, _05368_);
  not (_05382_, _02556_);
  not (_05383_, _02894_);
  not (_05384_, _04657_);
  nand (_05385_, _05379_, _05384_);
  or (_05386_, _05385_, _05383_);
  and (_05387_, _04449_, _03309_);
  or (_05388_, _05387_, _05268_);
  and (_05389_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05390_, _05389_, \oc8051_golden_model_1.PC [6]);
  and (_05391_, _05390_, _02674_);
  and (_05392_, _05391_, \oc8051_golden_model_1.PC [7]);
  nor (_05393_, _05391_, \oc8051_golden_model_1.PC [7]);
  nor (_05394_, _05393_, _05392_);
  not (_05395_, _05394_);
  nor (_05396_, _05395_, _02558_);
  and (_05397_, _02558_, \oc8051_golden_model_1.ACC [7]);
  nor (_05398_, _05397_, _05396_);
  nand (_05399_, _05398_, _05387_);
  and (_05400_, _05399_, _05388_);
  or (_05401_, _05400_, _03818_);
  not (_05402_, _03818_);
  nor (_05403_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05404_, _05403_, _03326_);
  nor (_05405_, _05404_, _02946_);
  nor (_05406_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05407_, _05406_, _02946_);
  and (_05408_, _05407_, _02877_);
  nor (_05409_, _05408_, _05405_);
  nor (_05410_, _05409_, _03328_);
  not (_05411_, _05410_);
  not (_05412_, _04242_);
  or (_05413_, _05412_, _03867_);
  not (_05414_, _03328_);
  and (_05415_, _03867_, _02799_);
  nor (_05416_, _05415_, _05414_);
  nand (_05417_, _05416_, _05413_);
  and (_05418_, _05417_, _05411_);
  nor (_05419_, _05403_, _03326_);
  nor (_05420_, _05419_, _05404_);
  nor (_05421_, _05420_, _03328_);
  not (_05422_, _05421_);
  or (_05423_, _04441_, _03867_);
  and (_05424_, _03867_, _03260_);
  nor (_05425_, _05424_, _05414_);
  nand (_05426_, _05425_, _05423_);
  and (_05427_, _05426_, _05422_);
  not (_05428_, _05427_);
  nor (_05429_, _03940_, _03328_);
  not (_05430_, _05429_);
  nor (_05431_, _04038_, _03867_);
  and (_05432_, _03672_, _03867_);
  or (_05433_, _05432_, _05414_);
  or (_05434_, _05433_, _05431_);
  nand (_05435_, _05434_, _05430_);
  or (_05436_, _03817_, _03867_);
  and (_05437_, _03867_, _02832_);
  nor (_05438_, _05437_, _05414_);
  nand (_05439_, _05438_, _05436_);
  nor (_05440_, _03328_, \oc8051_golden_model_1.SP [0]);
  not (_05441_, _05440_);
  and (_05442_, _05441_, _05439_);
  and (_05443_, _05442_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_05444_, _05441_, _05439_);
  and (_05445_, _05444_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_05446_, _05445_, _05443_);
  and (_05447_, _05446_, _05435_);
  and (_05448_, _05434_, _05430_);
  and (_05449_, _05442_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_05450_, _05444_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_05451_, _05450_, _05449_);
  and (_05452_, _05451_, _05448_);
  or (_05453_, _05452_, _05447_);
  nor (_05454_, _05453_, _05428_);
  and (_05455_, _05442_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_05456_, _05444_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _05435_);
  and (_05459_, _05442_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_05460_, _05444_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_05461_, _05460_, _05459_);
  and (_05462_, _05461_, _05448_);
  or (_05463_, _05462_, _05458_);
  nor (_05464_, _05463_, _05427_);
  nor (_05465_, _05464_, _05454_);
  nor (_05466_, _05465_, _05418_);
  not (_05467_, _05418_);
  and (_05468_, _05444_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_05469_, _05442_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_05470_, _05469_, _05468_);
  and (_05471_, _05470_, _05435_);
  and (_05472_, _05442_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_05473_, _05444_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_05474_, _05473_, _05472_);
  and (_05475_, _05474_, _05448_);
  or (_05476_, _05475_, _05471_);
  nor (_05477_, _05476_, _05428_);
  and (_05478_, _05442_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_05479_, _05444_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_05480_, _05479_, _05478_);
  and (_05481_, _05480_, _05435_);
  and (_05482_, _05442_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_05483_, _05444_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_05484_, _05483_, _05482_);
  and (_05485_, _05484_, _05448_);
  or (_05486_, _05485_, _05481_);
  nor (_05487_, _05486_, _05427_);
  nor (_05488_, _05487_, _05477_);
  nor (_05489_, _05488_, _05467_);
  nor (_05490_, _05489_, _05466_);
  or (_05491_, _05490_, _05402_);
  and (_05492_, _05491_, _05401_);
  or (_05493_, _05492_, _03822_);
  and (_05494_, _05250_, _04943_);
  and (_05495_, _05095_, _05044_);
  and (_05496_, _05142_, _04995_);
  and (_05497_, _05496_, _05495_);
  and (_05498_, _05497_, _05494_);
  and (_05499_, _05498_, _04837_);
  nor (_05500_, _05499_, _04733_);
  and (_05501_, _05499_, _04733_);
  nor (_05502_, _05501_, _05500_);
  or (_05503_, _05502_, _03823_);
  and (_05504_, _05503_, _05493_);
  or (_05505_, _05504_, _02894_);
  and (_05506_, _05505_, _05386_);
  or (_05507_, _05506_, _05382_);
  nor (_05508_, _05394_, _02556_);
  nor (_05509_, _05508_, _03845_);
  and (_05510_, _05509_, _05507_);
  nor (_05511_, _04623_, _04256_);
  or (_05512_, _05511_, _03853_);
  or (_05513_, _05512_, _05510_);
  and (_05514_, _05513_, _05381_);
  or (_05515_, _05514_, _02886_);
  and (_05516_, _04716_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05517_, _05516_);
  and (_05518_, _04719_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05519_, _05518_);
  and (_05520_, _04722_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05521_, _04724_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05522_, _05521_, _05520_);
  and (_05523_, _05522_, _05519_);
  and (_05524_, _05523_, _04715_);
  and (_05525_, _05524_, _05517_);
  and (_05526_, _05525_, _04696_);
  and (_05527_, _05526_, _04677_);
  and (_05528_, _05527_, _04625_);
  nand (_05529_, _05528_, _02886_);
  and (_05530_, _05529_, _02884_);
  and (_05531_, _05530_, _05515_);
  nor (_05532_, _05379_, _05384_);
  not (_05533_, _05532_);
  and (_05534_, _05533_, _05385_);
  and (_05535_, _05534_, _02883_);
  or (_05536_, _05535_, _05531_);
  and (_05537_, _05536_, _02561_);
  or (_05538_, _05395_, _02561_);
  nand (_05539_, _05538_, _02983_);
  or (_05540_, _05539_, _05537_);
  nand (_05541_, _05528_, _02984_);
  and (_05542_, _05541_, _05540_);
  or (_05543_, _05542_, _03867_);
  and (_05544_, _05490_, _02858_);
  nand (_05545_, _05527_, _03867_);
  or (_05546_, _05545_, _05544_);
  and (_05547_, _05546_, _04303_);
  and (_05548_, _05547_, _05543_);
  or (_05549_, _05548_, _05367_);
  and (_05550_, _05549_, _05325_);
  nor (_05551_, _02868_, _02849_);
  nand (_05552_, _05394_, _02578_);
  nand (_05553_, _05552_, _05551_);
  or (_05554_, _05553_, _05550_);
  or (_05555_, _05259_, _05551_);
  and (_05556_, _05555_, _05554_);
  or (_05557_, _05556_, _02857_);
  not (_05558_, _02857_);
  or (_05559_, _05490_, _05558_);
  and (_05560_, _05559_, _02853_);
  and (_05561_, _05560_, _05557_);
  not (_05562_, _05322_);
  not (_05563_, _05311_);
  nor (_05564_, _05563_, _04623_);
  not (_05565_, _05564_);
  not (_05566_, _03492_);
  and (_05567_, _03705_, _05566_);
  and (_05568_, _03063_, _01550_);
  and (_05569_, _03076_, _01548_);
  nor (_05570_, _05569_, _05568_);
  and (_05571_, _03100_, _01542_);
  and (_05572_, _03102_, _01538_);
  nor (_05573_, _05572_, _05571_);
  and (_05574_, _05573_, _05570_);
  and (_05575_, _03109_, _01546_);
  and (_05576_, _03086_, _01559_);
  nor (_05577_, _05576_, _05575_);
  and (_05578_, _03094_, _01540_);
  and (_05579_, _03096_, _01578_);
  nor (_05580_, _05579_, _05578_);
  and (_05581_, _05580_, _05577_);
  and (_05582_, _05581_, _05574_);
  and (_05583_, _03083_, _01571_);
  and (_05584_, _03112_, _01554_);
  nor (_05585_, _05584_, _05583_);
  and (_05586_, _03074_, _01567_);
  and (_05587_, _03114_, _01565_);
  nor (_05588_, _05587_, _05586_);
  and (_05589_, _05588_, _05585_);
  and (_05590_, _03088_, _01561_);
  and (_05591_, _03068_, _01576_);
  nor (_05592_, _05591_, _05590_);
  and (_05593_, _03107_, _33986_);
  and (_05594_, _03081_, _01569_);
  nor (_05595_, _05594_, _05593_);
  and (_05596_, _05595_, _05592_);
  and (_05597_, _05596_, _05589_);
  and (_05598_, _05597_, _05582_);
  and (_05599_, _05598_, _05563_);
  and (_05600_, _03083_, _01456_);
  and (_05601_, _03112_, _01466_);
  nor (_05602_, _05601_, _05600_);
  and (_05603_, _03107_, _33972_);
  and (_05604_, _03074_, _01460_);
  nor (_05605_, _05604_, _05603_);
  and (_05606_, _05605_, _05602_);
  and (_05607_, _03088_, _01480_);
  and (_05608_, _03094_, _01486_);
  nor (_05609_, _05608_, _05607_);
  and (_05610_, _03063_, _01464_);
  and (_05611_, _03086_, _01475_);
  nor (_05612_, _05611_, _05610_);
  and (_05613_, _05612_, _05609_);
  and (_05614_, _05613_, _05606_);
  and (_05615_, _03114_, _01450_);
  and (_05616_, _03096_, _01471_);
  nor (_05617_, _05616_, _05615_);
  and (_05618_, _03102_, _01448_);
  and (_05619_, _03076_, _01478_);
  nor (_05620_, _05619_, _05618_);
  and (_05621_, _05620_, _05617_);
  and (_05622_, _03081_, _01458_);
  and (_05623_, _03068_, _01488_);
  nor (_05624_, _05623_, _05622_);
  and (_05625_, _03100_, _01452_);
  and (_05626_, _03109_, _01473_);
  nor (_05627_, _05626_, _05625_);
  and (_05628_, _05627_, _05624_);
  and (_05629_, _05628_, _05621_);
  and (_05630_, _05629_, _05614_);
  and (_05631_, _03063_, _01509_);
  and (_05632_, _03076_, _01523_);
  nor (_05633_, _05632_, _05631_);
  and (_05634_, _03074_, _01503_);
  and (_05635_, _03114_, _01495_);
  nor (_05636_, _05635_, _05634_);
  and (_05637_, _05636_, _05633_);
  and (_05638_, _03109_, _01518_);
  and (_05639_, _03086_, _01520_);
  nor (_05640_, _05639_, _05638_);
  and (_05641_, _03094_, _01531_);
  and (_05642_, _03096_, _01516_);
  nor (_05643_, _05642_, _05641_);
  and (_05644_, _05643_, _05640_);
  and (_05645_, _05644_, _05637_);
  and (_05646_, _03081_, _01505_);
  and (_05647_, _03112_, _01501_);
  nor (_05648_, _05647_, _05646_);
  and (_05649_, _03107_, _33979_);
  and (_05650_, _03083_, _01511_);
  nor (_05651_, _05650_, _05649_);
  and (_05652_, _05651_, _05648_);
  and (_05653_, _03088_, _01525_);
  and (_05654_, _03068_, _01533_);
  nor (_05655_, _05654_, _05653_);
  and (_05656_, _03100_, _01497_);
  and (_05657_, _03102_, _01493_);
  nor (_05658_, _05657_, _05656_);
  and (_05659_, _05658_, _05655_);
  and (_05660_, _05659_, _05652_);
  and (_05661_, _05660_, _05645_);
  and (_05662_, _05661_, _05630_);
  and (_05663_, _05662_, _05599_);
  not (_05664_, _03120_);
  and (_05665_, _03302_, _05664_);
  and (_05666_, _05665_, _05663_);
  and (_05667_, _05666_, _05567_);
  and (_05668_, _05667_, \oc8051_golden_model_1.TMOD [7]);
  and (_05669_, _03302_, _03120_);
  nor (_05670_, _03705_, _03492_);
  and (_05671_, _05670_, _05663_);
  and (_05672_, _05671_, _05669_);
  and (_05673_, _05672_, \oc8051_golden_model_1.DPH [7]);
  nor (_05674_, _05673_, _05668_);
  not (_05675_, _03705_);
  and (_05676_, _05675_, _03492_);
  and (_05677_, _05676_, _05666_);
  and (_05678_, _05677_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05679_, _03302_, _03120_);
  and (_05680_, _05679_, _05663_);
  and (_05681_, _05680_, _05567_);
  and (_05682_, _05681_, \oc8051_golden_model_1.TH1 [7]);
  nor (_05683_, _05682_, _05678_);
  and (_05684_, _05683_, _05674_);
  and (_05685_, _03705_, _03492_);
  and (_05686_, _05685_, _05665_);
  nor (_05687_, _05661_, _05630_);
  and (_05688_, _05687_, _05599_);
  and (_05689_, _05688_, _05686_);
  and (_05690_, _05689_, \oc8051_golden_model_1.IP [7]);
  and (_05691_, _05685_, _05669_);
  nor (_05692_, _05598_, _05311_);
  and (_05693_, _05692_, _05691_);
  and (_05694_, _05693_, _05687_);
  and (_05695_, _05694_, \oc8051_golden_model_1.B [7]);
  nor (_05696_, _05695_, _05690_);
  not (_05697_, _05630_);
  and (_05698_, _05661_, _05697_);
  and (_05699_, _05698_, _05693_);
  and (_05700_, _05699_, \oc8051_golden_model_1.PSW [7]);
  not (_05701_, _05661_);
  and (_05702_, _05701_, _05630_);
  and (_05703_, _05702_, _05693_);
  and (_05704_, _05703_, \oc8051_golden_model_1.ACC [7]);
  nor (_05705_, _05704_, _05700_);
  and (_05706_, _05705_, _05696_);
  and (_05707_, _05702_, _05599_);
  and (_05708_, _05707_, _05686_);
  and (_05709_, _05708_, \oc8051_golden_model_1.IE [7]);
  and (_05710_, _05698_, _05599_);
  and (_05711_, _05665_, _05567_);
  and (_05712_, _05711_, _05710_);
  and (_05713_, _05712_, \oc8051_golden_model_1.SBUF [7]);
  and (_05714_, _05710_, _05686_);
  and (_05715_, _05714_, \oc8051_golden_model_1.SCON [7]);
  or (_05716_, _05715_, _05713_);
  nor (_05717_, _05716_, _05709_);
  and (_05718_, _05717_, _05706_);
  and (_05719_, _05718_, _05684_);
  and (_05720_, _05685_, _05680_);
  and (_05721_, _05720_, \oc8051_golden_model_1.TH0 [7]);
  and (_05722_, _05671_, _05665_);
  and (_05723_, _05722_, \oc8051_golden_model_1.TL1 [7]);
  nor (_05724_, _05723_, _05721_);
  and (_05725_, _05686_, _05663_);
  and (_05726_, _05725_, \oc8051_golden_model_1.TCON [7]);
  not (_05727_, _03302_);
  and (_05728_, _05727_, _03120_);
  and (_05729_, _05728_, _05671_);
  and (_05730_, _05729_, \oc8051_golden_model_1.PCON [7]);
  nor (_05731_, _05730_, _05726_);
  and (_05732_, _05731_, _05724_);
  and (_05733_, _05710_, _05691_);
  and (_05734_, _05733_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05735_, _05734_);
  and (_05736_, _05691_, _05663_);
  and (_05737_, _05736_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05738_, _05737_);
  and (_05739_, _05707_, _05691_);
  and (_05740_, _05739_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05741_, _05691_, _05688_);
  and (_05742_, _05741_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05743_, _05742_, _05740_);
  and (_05744_, _05743_, _05738_);
  and (_05745_, _05744_, _05735_);
  and (_05746_, _05669_, _05663_);
  and (_05747_, _05746_, _05567_);
  and (_05748_, _05747_, \oc8051_golden_model_1.SP [7]);
  and (_05749_, _05746_, _05676_);
  and (_05750_, _05749_, \oc8051_golden_model_1.DPL [7]);
  nor (_05751_, _05750_, _05748_);
  and (_05752_, _05751_, _05745_);
  and (_05753_, _05752_, _05732_);
  and (_05754_, _05753_, _05719_);
  and (_05755_, _05754_, _05565_);
  nor (_05756_, _05755_, _02853_);
  or (_05757_, _05756_, _05562_);
  or (_05758_, _05757_, _05561_);
  and (_05759_, _05758_, _05324_);
  and (_05760_, _05563_, _03885_);
  or (_05761_, _05760_, _02517_);
  or (_05762_, _05761_, _05759_);
  and (_05763_, _05395_, _02517_);
  nor (_05764_, _05763_, _05280_);
  and (_05765_, _05764_, _05762_);
  or (_05766_, _05765_, _05315_);
  and (_05767_, _05766_, _05278_);
  not (_05768_, \oc8051_golden_model_1.ACC [7]);
  nor (_05769_, _04732_, _05768_);
  and (_05770_, _04732_, _05768_);
  nor (_05771_, _05770_, _05769_);
  and (_05772_, _05771_, _05277_);
  or (_05773_, _05772_, _05767_);
  and (_05774_, _05773_, _05276_);
  and (_05775_, _05313_, _05275_);
  or (_05776_, _05775_, _05774_);
  and (_05777_, _05776_, _05273_);
  and (_05778_, _05769_, _03891_);
  or (_05779_, _05778_, _02533_);
  or (_05780_, _05779_, _05777_);
  not (_05781_, _03036_);
  nor (_05782_, _05781_, _02768_);
  and (_05783_, _05395_, _02533_);
  nor (_05784_, _05783_, _05782_);
  and (_05785_, _05784_, _05780_);
  not (_05786_, _03127_);
  nor (_05787_, _05786_, _02768_);
  not (_05788_, _05782_);
  nor (_05789_, _05312_, _05788_);
  or (_05790_, _05789_, _05787_);
  or (_05791_, _05790_, _05785_);
  not (_05792_, _02531_);
  nand (_05793_, _05770_, _05787_);
  and (_05794_, _05793_, _05792_);
  and (_05795_, _05794_, _05791_);
  nand (_05796_, _05394_, _02531_);
  nand (_05797_, _05796_, _05271_);
  or (_05798_, _05797_, _05795_);
  and (_05799_, _05798_, _05272_);
  or (_05800_, _05799_, _03909_);
  not (_05801_, _03908_);
  not (_05802_, _05490_);
  or (_05803_, _05442_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_05804_, _05444_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_05805_, _05804_, _05435_);
  and (_05806_, _05805_, _05803_);
  or (_05807_, _05444_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05808_, _05442_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_05809_, _05808_, _05448_);
  and (_05810_, _05809_, _05807_);
  nor (_05811_, _05810_, _05806_);
  nand (_05812_, _05811_, _05427_);
  or (_05813_, _05442_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_05814_, _05444_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_05815_, _05814_, _05435_);
  and (_05816_, _05815_, _05813_);
  or (_05817_, _05444_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05818_, _05442_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_05819_, _05818_, _05448_);
  and (_05820_, _05819_, _05817_);
  nor (_05821_, _05820_, _05816_);
  nand (_05822_, _05821_, _05428_);
  nand (_05823_, _05822_, _05812_);
  nand (_05824_, _05823_, _05467_);
  or (_05825_, _05442_, _04736_);
  or (_05826_, _05444_, _04734_);
  and (_05827_, _05826_, _05435_);
  nand (_05828_, _05827_, _05825_);
  or (_05829_, _05444_, _04742_);
  or (_05830_, _05442_, _04740_);
  and (_05831_, _05830_, _05448_);
  nand (_05832_, _05831_, _05829_);
  nand (_05833_, _05832_, _05828_);
  nand (_05834_, _05833_, _05427_);
  or (_05835_, _05444_, _04755_);
  or (_05836_, _05442_, _04757_);
  and (_05837_, _05836_, _05435_);
  nand (_05838_, _05837_, _05835_);
  or (_05839_, _05444_, _04751_);
  or (_05840_, _05442_, _04748_);
  and (_05841_, _05840_, _05448_);
  nand (_05842_, _05841_, _05839_);
  nand (_05843_, _05842_, _05838_);
  nand (_05844_, _05843_, _05428_);
  nand (_05845_, _05844_, _05834_);
  nand (_05846_, _05845_, _05418_);
  and (_05847_, _05846_, _05824_);
  not (_05848_, _05847_);
  or (_05849_, _05442_, \oc8051_golden_model_1.IRAM[9] [1]);
  or (_05850_, _05444_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_05851_, _05850_, _05435_);
  and (_05852_, _05851_, _05849_);
  or (_05853_, _05444_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_05854_, _05442_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_05855_, _05854_, _05448_);
  and (_05856_, _05855_, _05853_);
  nor (_05857_, _05856_, _05852_);
  nand (_05858_, _05857_, _05427_);
  or (_05859_, _05442_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_05860_, _05444_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_05861_, _05860_, _05435_);
  and (_05862_, _05861_, _05859_);
  or (_05863_, _05444_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_05864_, _05442_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_05865_, _05864_, _05448_);
  and (_05866_, _05865_, _05863_);
  nor (_05867_, _05866_, _05862_);
  nand (_05868_, _05867_, _05428_);
  nand (_05869_, _05868_, _05858_);
  nand (_05870_, _05869_, _05467_);
  or (_05871_, _05442_, _03951_);
  or (_05872_, _05444_, _03949_);
  and (_05873_, _05872_, _05435_);
  nand (_05874_, _05873_, _05871_);
  or (_05875_, _05444_, _03957_);
  or (_05876_, _05442_, _03955_);
  and (_05877_, _05876_, _05448_);
  nand (_05878_, _05877_, _05875_);
  nand (_05879_, _05878_, _05874_);
  nand (_05880_, _05879_, _05427_);
  or (_05881_, _05444_, _03969_);
  or (_05882_, _05442_, _03971_);
  and (_05883_, _05882_, _05435_);
  nand (_05884_, _05883_, _05881_);
  or (_05885_, _05444_, _03965_);
  or (_05886_, _05442_, _03963_);
  and (_05887_, _05886_, _05448_);
  nand (_05888_, _05887_, _05885_);
  nand (_05889_, _05888_, _05884_);
  nand (_05890_, _05889_, _05428_);
  nand (_05891_, _05890_, _05880_);
  nand (_05892_, _05891_, _05418_);
  nand (_05893_, _05892_, _05870_);
  or (_05894_, _05442_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_05895_, _05444_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_05896_, _05895_, _05435_);
  and (_05897_, _05896_, _05894_);
  or (_05898_, _05444_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_05899_, _05442_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_05900_, _05899_, _05448_);
  and (_05901_, _05900_, _05898_);
  nor (_05902_, _05901_, _05897_);
  nand (_05903_, _05902_, _05427_);
  or (_05904_, _05442_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_05905_, _05444_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_05906_, _05905_, _05435_);
  and (_05907_, _05906_, _05904_);
  or (_05908_, _05444_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_05909_, _05442_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_05910_, _05909_, _05448_);
  and (_05911_, _05910_, _05908_);
  nor (_05912_, _05911_, _05907_);
  nand (_05913_, _05912_, _05428_);
  nand (_05914_, _05913_, _05903_);
  nand (_05915_, _05914_, _05467_);
  or (_05916_, _05442_, _03759_);
  or (_05917_, _05444_, _03375_);
  and (_05918_, _05917_, _05435_);
  nand (_05919_, _05918_, _05916_);
  or (_05920_, _05444_, _03767_);
  or (_05921_, _05442_, _03764_);
  and (_05922_, _05921_, _05448_);
  nand (_05923_, _05922_, _05920_);
  nand (_05924_, _05923_, _05919_);
  nand (_05925_, _05924_, _05427_);
  or (_05926_, _05444_, _03780_);
  or (_05927_, _05442_, _03782_);
  and (_05928_, _05927_, _05435_);
  nand (_05929_, _05928_, _05926_);
  or (_05930_, _05444_, _03776_);
  or (_05931_, _05442_, _03774_);
  and (_05932_, _05931_, _05448_);
  nand (_05933_, _05932_, _05930_);
  nand (_05934_, _05933_, _05929_);
  nand (_05935_, _05934_, _05428_);
  nand (_05936_, _05935_, _05925_);
  nand (_05937_, _05936_, _05418_);
  nand (_05938_, _05937_, _05915_);
  and (_05939_, _05938_, _05893_);
  or (_05940_, _05442_, \oc8051_golden_model_1.IRAM[9] [3]);
  or (_05941_, _05444_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_05942_, _05941_, _05435_);
  and (_05943_, _05942_, _05940_);
  or (_05944_, _05444_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05945_, _05442_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_05946_, _05945_, _05448_);
  and (_05947_, _05946_, _05944_);
  nor (_05948_, _05947_, _05943_);
  nand (_05949_, _05948_, _05427_);
  or (_05950_, _05442_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_05951_, _05444_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_05952_, _05951_, _05435_);
  and (_05953_, _05952_, _05950_);
  or (_05954_, _05444_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05955_, _05442_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_05956_, _05955_, _05448_);
  and (_05957_, _05956_, _05954_);
  nor (_05958_, _05957_, _05953_);
  nand (_05959_, _05958_, _05428_);
  nand (_05960_, _05959_, _05949_);
  nand (_05961_, _05960_, _05467_);
  or (_05962_, _05442_, _04192_);
  or (_05963_, _05444_, _04190_);
  and (_05964_, _05963_, _05435_);
  nand (_05965_, _05964_, _05962_);
  or (_05966_, _05444_, _04198_);
  or (_05967_, _05442_, _04196_);
  and (_05968_, _05967_, _05448_);
  nand (_05969_, _05968_, _05966_);
  nand (_05970_, _05969_, _05965_);
  nand (_05971_, _05970_, _05427_);
  or (_05972_, _05444_, _04210_);
  or (_05973_, _05442_, _04212_);
  and (_05974_, _05973_, _05435_);
  nand (_05975_, _05974_, _05972_);
  or (_05976_, _05444_, _04206_);
  or (_05977_, _05442_, _04204_);
  and (_05978_, _05977_, _05448_);
  nand (_05979_, _05978_, _05976_);
  nand (_05980_, _05979_, _05975_);
  nand (_05981_, _05980_, _05428_);
  nand (_05982_, _05981_, _05971_);
  nand (_05983_, _05982_, _05418_);
  nand (_05984_, _05983_, _05961_);
  or (_05985_, _05442_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_05986_, _05444_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_05987_, _05986_, _05435_);
  and (_05988_, _05987_, _05985_);
  or (_05989_, _05444_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_05990_, _05442_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_05991_, _05990_, _05448_);
  and (_05992_, _05991_, _05989_);
  nor (_05993_, _05992_, _05988_);
  nand (_05994_, _05993_, _05427_);
  or (_05995_, _05442_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_05996_, _05444_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_05997_, _05996_, _05435_);
  and (_05998_, _05997_, _05995_);
  or (_05999_, _05444_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_06000_, _05442_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_06001_, _06000_, _05448_);
  and (_06002_, _06001_, _05999_);
  nor (_06003_, _06002_, _05998_);
  nand (_06004_, _06003_, _05428_);
  nand (_06005_, _06004_, _05994_);
  nand (_06006_, _06005_, _05467_);
  or (_06007_, _05442_, _04375_);
  or (_06008_, _05444_, _04372_);
  and (_06009_, _06008_, _05435_);
  nand (_06010_, _06009_, _06007_);
  or (_06011_, _05444_, _04384_);
  or (_06012_, _05442_, _04381_);
  and (_06013_, _06012_, _05448_);
  nand (_06014_, _06013_, _06011_);
  nand (_06015_, _06014_, _06010_);
  nand (_06016_, _06015_, _05427_);
  or (_06017_, _05444_, _04402_);
  or (_06018_, _05442_, _04405_);
  and (_06019_, _06018_, _05435_);
  nand (_06020_, _06019_, _06017_);
  or (_06021_, _05444_, _04396_);
  or (_06022_, _05442_, _04393_);
  and (_06023_, _06022_, _05448_);
  nand (_06024_, _06023_, _06021_);
  nand (_06025_, _06024_, _06020_);
  nand (_06026_, _06025_, _05428_);
  nand (_06027_, _06026_, _06016_);
  nand (_06028_, _06027_, _05418_);
  nand (_06029_, _06028_, _06006_);
  and (_06030_, _06029_, _05984_);
  and (_06031_, _06030_, _05939_);
  or (_06032_, _05442_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_06033_, _05444_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_06034_, _06033_, _05435_);
  and (_06035_, _06034_, _06032_);
  or (_06036_, _05444_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06037_, _05442_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_06038_, _06037_, _05448_);
  and (_06039_, _06038_, _06036_);
  nor (_06040_, _06039_, _06035_);
  nand (_06041_, _06040_, _05427_);
  or (_06042_, _05442_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_06043_, _05444_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_06044_, _06043_, _05435_);
  and (_06045_, _06044_, _06042_);
  or (_06046_, _05444_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06047_, _05442_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_06048_, _06047_, _05448_);
  and (_06049_, _06048_, _06046_);
  nor (_06050_, _06049_, _06045_);
  nand (_06051_, _06050_, _05428_);
  nand (_06052_, _06051_, _06041_);
  nand (_06053_, _06052_, _05467_);
  or (_06054_, _05442_, _04841_);
  or (_06055_, _05444_, _04839_);
  and (_06056_, _06055_, _05435_);
  nand (_06057_, _06056_, _06054_);
  or (_06058_, _05444_, _04847_);
  or (_06059_, _05442_, _04845_);
  and (_06060_, _06059_, _05448_);
  nand (_06061_, _06060_, _06058_);
  nand (_06062_, _06061_, _06057_);
  nand (_06063_, _06062_, _05427_);
  or (_06064_, _05444_, _04860_);
  or (_06065_, _05442_, _04862_);
  and (_06066_, _06065_, _05435_);
  nand (_06067_, _06066_, _06064_);
  or (_06068_, _05444_, _04856_);
  or (_06069_, _05442_, _04854_);
  and (_06070_, _06069_, _05448_);
  nand (_06071_, _06070_, _06068_);
  nand (_06072_, _06071_, _06067_);
  nand (_06073_, _06072_, _05428_);
  nand (_06074_, _06073_, _06063_);
  nand (_06075_, _06074_, _05418_);
  nand (_06076_, _06075_, _06053_);
  or (_06077_, _05442_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_06078_, _05444_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_06079_, _06078_, _05435_);
  and (_06080_, _06079_, _06077_);
  or (_06081_, _05444_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06082_, _05442_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_06083_, _06082_, _05448_);
  and (_06084_, _06083_, _06081_);
  nor (_06085_, _06084_, _06080_);
  nand (_06086_, _06085_, _05427_);
  or (_06087_, _05442_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_06088_, _05444_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_06089_, _06088_, _05435_);
  and (_06090_, _06089_, _06087_);
  or (_06091_, _05444_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06092_, _05442_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_06093_, _06092_, _05448_);
  and (_06094_, _06093_, _06091_);
  nor (_06095_, _06094_, _06090_);
  nand (_06096_, _06095_, _05428_);
  nand (_06097_, _06096_, _06086_);
  nand (_06098_, _06097_, _05467_);
  or (_06099_, _05442_, _05148_);
  or (_06100_, _05444_, _05146_);
  and (_06101_, _06100_, _05435_);
  nand (_06102_, _06101_, _06099_);
  or (_06103_, _05444_, _05154_);
  or (_06104_, _05442_, _05152_);
  and (_06105_, _06104_, _05448_);
  nand (_06106_, _06105_, _06103_);
  nand (_06107_, _06106_, _06102_);
  nand (_06108_, _06107_, _05427_);
  or (_06109_, _05444_, _05166_);
  or (_06110_, _05442_, _05168_);
  and (_06111_, _06110_, _05435_);
  nand (_06112_, _06111_, _06109_);
  or (_06113_, _05444_, _05162_);
  or (_06114_, _05442_, _05160_);
  and (_06115_, _06114_, _05448_);
  nand (_06116_, _06115_, _06113_);
  nand (_06117_, _06116_, _06112_);
  nand (_06118_, _06117_, _05428_);
  nand (_06119_, _06118_, _06108_);
  nand (_06120_, _06119_, _05418_);
  nand (_06121_, _06120_, _06098_);
  and (_06122_, _06121_, _06076_);
  and (_06123_, _06122_, _06031_);
  and (_06124_, _06123_, _05848_);
  nor (_06125_, _06124_, _05802_);
  and (_06126_, _06124_, _05802_);
  or (_06127_, _06126_, _06125_);
  or (_06128_, _06127_, _03910_);
  and (_06129_, _06128_, _05801_);
  and (_06130_, _06129_, _05800_);
  and (_06131_, _05502_, _03908_);
  or (_06132_, _06131_, _03004_);
  or (_06133_, _06132_, _06130_);
  and (_06134_, _02251_, _02232_);
  and (_06135_, _06134_, _05390_);
  and (_06136_, _06135_, \oc8051_golden_model_1.PC [7]);
  nor (_06137_, _06135_, \oc8051_golden_model_1.PC [7]);
  nor (_06138_, _06137_, _06136_);
  not (_06139_, _06138_);
  nand (_06140_, _06139_, _03004_);
  and (_06141_, _06140_, _06133_);
  or (_06142_, _06141_, _02528_);
  and (_06143_, _05395_, _02528_);
  nor (_06144_, _06143_, _03627_);
  and (_06145_, _06144_, _06142_);
  and (_06146_, _05364_, _03627_);
  and (_06147_, _02862_, _02525_);
  and (_06148_, _02864_, _02525_);
  nor (_06149_, _06148_, _06147_);
  not (_06150_, _04142_);
  nand (_06151_, _03010_, _02525_);
  and (_06152_, _06151_, _03585_);
  and (_06153_, _06152_, _06150_);
  and (_06154_, _06153_, _06149_);
  not (_06155_, _06154_);
  or (_06156_, _06155_, _06146_);
  or (_06157_, _06156_, _06145_);
  not (_06158_, _04787_);
  not (_06159_, _04896_);
  not (_06160_, _05202_);
  and (_06161_, _04005_, _03817_);
  nor (_06162_, _04440_, _04242_);
  and (_06163_, _06162_, _06161_);
  and (_06164_, _06163_, _06160_);
  and (_06165_, _06164_, _06159_);
  and (_06166_, _06165_, _06158_);
  and (_06167_, _06166_, _04623_);
  nor (_06168_, _06166_, _04623_);
  or (_06169_, _06168_, _06167_);
  or (_06170_, _06169_, _06154_);
  and (_06171_, _06170_, _06157_);
  or (_06172_, _06171_, _03926_);
  and (_06173_, _05892_, _05870_);
  and (_06174_, _05937_, _05915_);
  and (_06175_, _06174_, _06173_);
  and (_06176_, _05983_, _05961_);
  and (_06177_, _06028_, _06006_);
  and (_06178_, _06177_, _06176_);
  and (_06179_, _06178_, _06175_);
  and (_06180_, _06075_, _06053_);
  and (_06181_, _06120_, _06098_);
  and (_06182_, _06181_, _06180_);
  and (_06183_, _06182_, _06179_);
  and (_06184_, _06183_, _05847_);
  and (_06185_, _06184_, _05490_);
  nor (_06186_, _06184_, _05490_);
  nor (_06187_, _06186_, _06185_);
  or (_06188_, _06187_, _03927_);
  and (_06189_, _06188_, _04176_);
  and (_06190_, _06189_, _06172_);
  or (_06191_, _06190_, _05258_);
  and (_06192_, _06191_, _04557_);
  or (_06193_, _06192_, _04566_);
  and (_06194_, _06193_, _04556_);
  not (_06195_, _03004_);
  and (_06196_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06197_, _06196_, \oc8051_golden_model_1.PC [10]);
  and (_06198_, _06197_, _06136_);
  and (_06199_, _06198_, \oc8051_golden_model_1.PC [11]);
  and (_06200_, _06199_, \oc8051_golden_model_1.PC [12]);
  and (_06201_, _06200_, \oc8051_golden_model_1.PC [13]);
  and (_06202_, _06201_, \oc8051_golden_model_1.PC [14]);
  nor (_06203_, _06202_, \oc8051_golden_model_1.PC [15]);
  and (_06204_, _06196_, _06136_);
  and (_06205_, _06204_, \oc8051_golden_model_1.PC [10]);
  and (_06206_, _06205_, \oc8051_golden_model_1.PC [11]);
  and (_06207_, _06206_, \oc8051_golden_model_1.PC [12]);
  and (_06208_, _06207_, \oc8051_golden_model_1.PC [13]);
  and (_06209_, _06208_, \oc8051_golden_model_1.PC [14]);
  and (_06210_, _06209_, \oc8051_golden_model_1.PC [15]);
  nor (_06211_, _06210_, _06203_);
  or (_06212_, _06211_, _06195_);
  and (_06213_, _06197_, _05392_);
  and (_06214_, _06213_, \oc8051_golden_model_1.PC [11]);
  and (_06215_, _06214_, \oc8051_golden_model_1.PC [12]);
  and (_06216_, _06215_, \oc8051_golden_model_1.PC [13]);
  and (_06217_, _06216_, \oc8051_golden_model_1.PC [14]);
  nor (_06218_, _06217_, \oc8051_golden_model_1.PC [15]);
  and (_06219_, _05392_, \oc8051_golden_model_1.PC [8]);
  and (_06220_, _06219_, \oc8051_golden_model_1.PC [9]);
  and (_06221_, _06220_, \oc8051_golden_model_1.PC [10]);
  and (_06222_, _06221_, \oc8051_golden_model_1.PC [11]);
  and (_06223_, _06222_, \oc8051_golden_model_1.PC [12]);
  and (_06224_, _06223_, \oc8051_golden_model_1.PC [13]);
  and (_06225_, _06224_, \oc8051_golden_model_1.PC [14]);
  and (_06226_, _06225_, \oc8051_golden_model_1.PC [15]);
  nor (_06227_, _06226_, _06218_);
  or (_06228_, _06227_, _03004_);
  and (_06229_, _06228_, _06212_);
  and (_06230_, _06229_, _04551_);
  and (_06231_, _06230_, _04554_);
  or (_32484_, _06231_, _06194_);
  not (_06232_, \oc8051_golden_model_1.B [7]);
  nor (_06233_, _34698_, _06232_);
  nor (_06234_, _04705_, _06232_);
  not (_06235_, _04705_);
  nor (_06236_, _06235_, _04623_);
  or (_06237_, _06236_, _06234_);
  and (_06238_, _04148_, _02520_);
  not (_06239_, _02520_);
  nor (_06240_, _02977_, _06239_);
  nor (_06241_, _06240_, _06238_);
  or (_06242_, _06241_, _06237_);
  nor (_06243_, _05338_, _06232_);
  and (_06244_, _05380_, _05338_);
  or (_06245_, _06244_, _06243_);
  and (_06246_, _06245_, _02887_);
  and (_06247_, _05502_, _04705_);
  or (_06248_, _06247_, _06234_);
  or (_06249_, _06248_, _03821_);
  and (_06250_, _04705_, \oc8051_golden_model_1.ACC [7]);
  or (_06251_, _06250_, _06234_);
  and (_06252_, _06251_, _03825_);
  nor (_06253_, _03825_, _06232_);
  or (_06254_, _06253_, _02952_);
  or (_06255_, _06254_, _06252_);
  and (_06256_, _06255_, _02892_);
  and (_06257_, _06256_, _06249_);
  and (_06258_, _05385_, _05338_);
  or (_06259_, _06258_, _06243_);
  and (_06260_, _06259_, _02891_);
  or (_06261_, _06260_, _02947_);
  or (_06262_, _06261_, _06257_);
  or (_06263_, _06237_, _03327_);
  and (_06264_, _06263_, _06262_);
  or (_06265_, _06264_, _02950_);
  or (_06266_, _06251_, _02959_);
  and (_06267_, _06266_, _02888_);
  and (_06268_, _06267_, _06265_);
  or (_06269_, _06268_, _06246_);
  and (_06270_, _06269_, _02881_);
  and (_06271_, _03024_, _02980_);
  or (_06272_, _06243_, _05533_);
  and (_06273_, _06272_, _02880_);
  and (_06274_, _06273_, _06259_);
  or (_06275_, _06274_, _06271_);
  or (_06276_, _06275_, _06270_);
  not (_06277_, _06271_);
  and (_06278_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06279_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06280_, _06279_, _06278_);
  and (_06281_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06282_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_06283_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_06284_, _06283_, _06282_);
  nor (_06285_, _06284_, _06280_);
  and (_06286_, _06285_, _06281_);
  nor (_06287_, _06286_, _06280_);
  and (_06288_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06289_, _06288_, _06283_);
  and (_06290_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06291_, _06290_, _06278_);
  nor (_06292_, _06291_, _06289_);
  not (_06293_, _06292_);
  nor (_06294_, _06293_, _06287_);
  and (_06295_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06296_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06297_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06298_, _06297_, _06296_);
  nor (_06299_, _06297_, _06296_);
  nor (_06300_, _06299_, _06298_);
  and (_06301_, _06300_, _06295_);
  nor (_06302_, _06300_, _06295_);
  nor (_06303_, _06302_, _06301_);
  and (_06304_, _06293_, _06287_);
  nor (_06305_, _06304_, _06294_);
  and (_06306_, _06305_, _06303_);
  nor (_06307_, _06306_, _06294_);
  not (_06308_, _06283_);
  and (_06309_, _06288_, _06308_);
  and (_06310_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06311_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06312_, _06311_, _06296_);
  and (_06313_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06314_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06315_, _06314_, _06313_);
  nor (_06316_, _06315_, _06312_);
  and (_06317_, _06316_, _06310_);
  nor (_06318_, _06316_, _06310_);
  nor (_06319_, _06318_, _06317_);
  and (_06320_, _06319_, _06309_);
  nor (_06321_, _06319_, _06309_);
  nor (_06322_, _06321_, _06320_);
  not (_06323_, _06322_);
  nor (_06324_, _06323_, _06307_);
  and (_06325_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06326_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06327_, _06326_, _06325_);
  nor (_06328_, _06301_, _06298_);
  and (_06329_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06330_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06331_, _06330_, _06329_);
  nor (_06332_, _06330_, _06329_);
  nor (_06333_, _06332_, _06331_);
  not (_06334_, _06333_);
  nor (_06335_, _06334_, _06328_);
  and (_06336_, _06334_, _06328_);
  nor (_06337_, _06336_, _06335_);
  and (_06338_, _06337_, _06327_);
  nor (_06339_, _06337_, _06327_);
  nor (_06340_, _06339_, _06338_);
  and (_06341_, _06323_, _06307_);
  nor (_06342_, _06341_, _06324_);
  and (_06343_, _06342_, _06340_);
  nor (_06344_, _06343_, _06324_);
  nor (_06345_, _06317_, _06312_);
  and (_06346_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06347_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06348_, _06347_, _06346_);
  nor (_06349_, _06347_, _06346_);
  nor (_06350_, _06349_, _06348_);
  not (_06351_, _06350_);
  nor (_06352_, _06351_, _06345_);
  and (_06353_, _06351_, _06345_);
  nor (_06354_, _06353_, _06352_);
  and (_06355_, _06354_, _06331_);
  nor (_06356_, _06354_, _06331_);
  nor (_06357_, _06356_, _06355_);
  nor (_06358_, _06320_, _06289_);
  and (_06359_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_06360_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_06361_, _06360_, _06311_);
  nor (_06362_, _06360_, _06311_);
  nor (_06363_, _06362_, _06361_);
  and (_06364_, _06363_, _06359_);
  nor (_06365_, _06363_, _06359_);
  nor (_06366_, _06365_, _06364_);
  not (_06367_, _06366_);
  nor (_06368_, _06367_, _06358_);
  and (_06369_, _06367_, _06358_);
  nor (_06370_, _06369_, _06368_);
  and (_06371_, _06370_, _06357_);
  nor (_06372_, _06370_, _06357_);
  nor (_06373_, _06372_, _06371_);
  not (_06374_, _06373_);
  nor (_06375_, _06374_, _06344_);
  nor (_06376_, _06338_, _06335_);
  not (_06377_, _06376_);
  and (_06378_, _06374_, _06344_);
  nor (_06379_, _06378_, _06375_);
  and (_06380_, _06379_, _06377_);
  nor (_06381_, _06380_, _06375_);
  nor (_06382_, _06355_, _06352_);
  not (_06383_, _06382_);
  nor (_06384_, _06371_, _06368_);
  not (_06385_, _06384_);
  and (_06386_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_06387_, _06386_, _06311_);
  and (_06388_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_06389_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_06390_, _06389_, _06388_);
  nor (_06391_, _06390_, _06387_);
  nor (_06392_, _06364_, _06361_);
  and (_06393_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_06394_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_06395_, _06394_, _06393_);
  nor (_06396_, _06394_, _06393_);
  nor (_06397_, _06396_, _06395_);
  not (_06398_, _06397_);
  nor (_06399_, _06398_, _06392_);
  and (_06400_, _06398_, _06392_);
  nor (_06401_, _06400_, _06399_);
  and (_06402_, _06401_, _06348_);
  nor (_06403_, _06401_, _06348_);
  nor (_06404_, _06403_, _06402_);
  and (_06405_, _06404_, _06391_);
  nor (_06406_, _06404_, _06391_);
  nor (_06407_, _06406_, _06405_);
  and (_06408_, _06407_, _06385_);
  nor (_06409_, _06407_, _06385_);
  nor (_06410_, _06409_, _06408_);
  and (_06411_, _06410_, _06383_);
  nor (_06412_, _06410_, _06383_);
  nor (_06413_, _06412_, _06411_);
  not (_06414_, _06413_);
  nor (_06415_, _06414_, _06381_);
  nor (_06416_, _06411_, _06408_);
  nor (_06417_, _06402_, _06399_);
  not (_06418_, _06417_);
  and (_06419_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_06420_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_06421_, _06420_, _06419_);
  nor (_06422_, _06420_, _06419_);
  nor (_06423_, _06422_, _06421_);
  and (_06424_, _06423_, _06387_);
  nor (_06425_, _06423_, _06387_);
  nor (_06426_, _06425_, _06424_);
  and (_06427_, _06426_, _06395_);
  nor (_06428_, _06426_, _06395_);
  nor (_06429_, _06428_, _06427_);
  and (_06430_, _06429_, _06386_);
  nor (_06431_, _06429_, _06386_);
  nor (_06432_, _06431_, _06430_);
  and (_06433_, _06432_, _06405_);
  nor (_06434_, _06432_, _06405_);
  nor (_06435_, _06434_, _06433_);
  and (_06436_, _06435_, _06418_);
  nor (_06437_, _06435_, _06418_);
  nor (_06438_, _06437_, _06436_);
  not (_06439_, _06438_);
  nor (_06440_, _06439_, _06416_);
  and (_06441_, _06439_, _06416_);
  nor (_06442_, _06441_, _06440_);
  and (_06443_, _06442_, _06415_);
  nor (_06444_, _06436_, _06433_);
  nor (_06445_, _06427_, _06424_);
  not (_06446_, _06445_);
  and (_06447_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_06448_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_06449_, _06448_, _06447_);
  nor (_06450_, _06448_, _06447_);
  nor (_06451_, _06450_, _06449_);
  and (_06452_, _06451_, _06421_);
  nor (_06453_, _06451_, _06421_);
  nor (_06454_, _06453_, _06452_);
  and (_06455_, _06454_, _06430_);
  nor (_06456_, _06454_, _06430_);
  nor (_06457_, _06456_, _06455_);
  and (_06458_, _06457_, _06446_);
  nor (_06459_, _06457_, _06446_);
  nor (_06460_, _06459_, _06458_);
  not (_06461_, _06460_);
  nor (_06462_, _06461_, _06444_);
  and (_06463_, _06461_, _06444_);
  nor (_06464_, _06463_, _06462_);
  and (_06465_, _06464_, _06440_);
  nor (_06466_, _06464_, _06440_);
  nor (_06467_, _06466_, _06465_);
  and (_06468_, _06467_, _06443_);
  nor (_06469_, _06467_, _06443_);
  nor (_06470_, _06469_, _06468_);
  and (_06471_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_06472_, _06471_, _06283_);
  and (_06473_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_06474_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_06475_, _06474_, _06279_);
  nor (_06476_, _06475_, _06472_);
  and (_06477_, _06476_, _06473_);
  nor (_06478_, _06477_, _06472_);
  not (_06479_, _06478_);
  nor (_06480_, _06285_, _06281_);
  nor (_06481_, _06480_, _06286_);
  and (_06482_, _06481_, _06479_);
  and (_06483_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_06484_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_06485_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_06486_, _06485_, _06484_);
  nor (_06487_, _06485_, _06484_);
  nor (_06488_, _06487_, _06486_);
  and (_06489_, _06488_, _06483_);
  nor (_06490_, _06488_, _06483_);
  nor (_06491_, _06490_, _06489_);
  nor (_06492_, _06481_, _06479_);
  nor (_06493_, _06492_, _06482_);
  and (_06494_, _06493_, _06491_);
  nor (_06495_, _06494_, _06482_);
  nor (_06496_, _06305_, _06303_);
  nor (_06497_, _06496_, _06306_);
  not (_06498_, _06497_);
  nor (_06499_, _06498_, _06495_);
  and (_06500_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_06501_, _06500_, _06326_);
  nor (_06502_, _06489_, _06486_);
  nor (_06503_, _06326_, _06325_);
  nor (_06504_, _06503_, _06327_);
  not (_06505_, _06504_);
  nor (_06506_, _06505_, _06502_);
  and (_06507_, _06505_, _06502_);
  nor (_06508_, _06507_, _06506_);
  and (_06509_, _06508_, _06501_);
  nor (_06510_, _06508_, _06501_);
  nor (_06511_, _06510_, _06509_);
  and (_06512_, _06498_, _06495_);
  nor (_06513_, _06512_, _06499_);
  and (_06514_, _06513_, _06511_);
  nor (_06515_, _06514_, _06499_);
  nor (_06516_, _06342_, _06340_);
  nor (_06517_, _06516_, _06343_);
  not (_06518_, _06517_);
  nor (_06519_, _06518_, _06515_);
  nor (_06520_, _06509_, _06506_);
  not (_06521_, _06520_);
  and (_06522_, _06518_, _06515_);
  nor (_06523_, _06522_, _06519_);
  and (_06524_, _06523_, _06521_);
  nor (_06525_, _06524_, _06519_);
  nor (_06526_, _06379_, _06377_);
  nor (_06527_, _06526_, _06380_);
  not (_06528_, _06527_);
  nor (_06529_, _06528_, _06525_);
  and (_06530_, _06414_, _06381_);
  nor (_06531_, _06530_, _06415_);
  and (_06532_, _06531_, _06529_);
  nor (_06533_, _06442_, _06415_);
  nor (_06534_, _06533_, _06443_);
  and (_06535_, _06534_, _06532_);
  and (_06536_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_06537_, _06536_, _06471_);
  and (_06538_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_06539_, _06536_, _06471_);
  nor (_06540_, _06539_, _06537_);
  and (_06541_, _06540_, _06538_);
  nor (_06542_, _06541_, _06537_);
  not (_06543_, _06542_);
  nor (_06544_, _06476_, _06473_);
  nor (_06545_, _06544_, _06477_);
  and (_06546_, _06545_, _06543_);
  and (_06547_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_06548_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_06549_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_06550_, _06549_, _06548_);
  nor (_06551_, _06549_, _06548_);
  nor (_06552_, _06551_, _06550_);
  and (_06553_, _06552_, _06547_);
  nor (_06554_, _06552_, _06547_);
  nor (_06555_, _06554_, _06553_);
  nor (_06556_, _06545_, _06543_);
  nor (_06557_, _06556_, _06546_);
  and (_06558_, _06557_, _06555_);
  nor (_06559_, _06558_, _06546_);
  not (_06560_, _06559_);
  nor (_06561_, _06493_, _06491_);
  nor (_06562_, _06561_, _06494_);
  and (_06563_, _06562_, _06560_);
  nor (_06564_, _06553_, _06550_);
  and (_06565_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_06566_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_06567_, _06566_, _06565_);
  nor (_06568_, _06567_, _06501_);
  not (_06569_, _06568_);
  nor (_06570_, _06569_, _06564_);
  and (_06571_, _06569_, _06564_);
  nor (_06572_, _06571_, _06570_);
  nor (_06573_, _06562_, _06560_);
  nor (_06574_, _06573_, _06563_);
  and (_06575_, _06574_, _06572_);
  nor (_06576_, _06575_, _06563_);
  nor (_06577_, _06513_, _06511_);
  nor (_06578_, _06577_, _06514_);
  not (_06579_, _06578_);
  nor (_06580_, _06579_, _06576_);
  and (_06581_, _06579_, _06576_);
  nor (_06582_, _06581_, _06580_);
  and (_06583_, _06582_, _06570_);
  nor (_06584_, _06583_, _06580_);
  nor (_06585_, _06523_, _06521_);
  nor (_06586_, _06585_, _06524_);
  not (_06587_, _06586_);
  nor (_06588_, _06587_, _06584_);
  and (_06589_, _06528_, _06525_);
  nor (_06590_, _06589_, _06529_);
  and (_06591_, _06590_, _06588_);
  nor (_06592_, _06531_, _06529_);
  nor (_06593_, _06592_, _06532_);
  and (_06594_, _06593_, _06591_);
  nor (_06595_, _06593_, _06591_);
  nor (_06596_, _06595_, _06594_);
  and (_06597_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_06598_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_06599_, _06598_, _06597_);
  and (_06600_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06601_, _06598_, _06597_);
  nor (_06602_, _06601_, _06599_);
  and (_06603_, _06602_, _06600_);
  nor (_06604_, _06603_, _06599_);
  not (_06605_, _06604_);
  nor (_06606_, _06540_, _06538_);
  nor (_06607_, _06606_, _06541_);
  and (_06608_, _06607_, _06605_);
  and (_06609_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_06610_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_06611_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_06612_, _06611_, _06610_);
  nor (_06613_, _06611_, _06610_);
  nor (_06614_, _06613_, _06612_);
  and (_06615_, _06614_, _06609_);
  nor (_06616_, _06614_, _06609_);
  nor (_06617_, _06616_, _06615_);
  nor (_06618_, _06607_, _06605_);
  nor (_06619_, _06618_, _06608_);
  and (_06620_, _06619_, _06617_);
  nor (_06621_, _06620_, _06608_);
  not (_06622_, _06621_);
  nor (_06623_, _06557_, _06555_);
  nor (_06624_, _06623_, _06558_);
  and (_06625_, _06624_, _06622_);
  not (_06626_, _06500_);
  nor (_06627_, _06615_, _06612_);
  nor (_06628_, _06627_, _06626_);
  and (_06629_, _06627_, _06626_);
  nor (_06630_, _06629_, _06628_);
  nor (_06631_, _06624_, _06622_);
  nor (_06632_, _06631_, _06625_);
  and (_06633_, _06632_, _06630_);
  nor (_06634_, _06633_, _06625_);
  not (_06635_, _06634_);
  nor (_06636_, _06574_, _06572_);
  nor (_06637_, _06636_, _06575_);
  and (_06638_, _06637_, _06635_);
  nor (_06639_, _06637_, _06635_);
  nor (_06640_, _06639_, _06638_);
  and (_06641_, _06640_, _06628_);
  nor (_06642_, _06641_, _06638_);
  nor (_06643_, _06582_, _06570_);
  nor (_06644_, _06643_, _06583_);
  not (_06645_, _06644_);
  nor (_06646_, _06645_, _06642_);
  and (_06647_, _06587_, _06584_);
  nor (_06648_, _06647_, _06588_);
  and (_06649_, _06648_, _06646_);
  nor (_06650_, _06590_, _06588_);
  nor (_06651_, _06650_, _06591_);
  and (_06652_, _06651_, _06649_);
  nor (_06653_, _06651_, _06649_);
  nor (_06654_, _06653_, _06652_);
  and (_06655_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_06656_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_06657_, _06656_, _06655_);
  and (_06658_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06659_, _06656_, _06655_);
  nor (_06660_, _06659_, _06657_);
  and (_06661_, _06660_, _06658_);
  nor (_06662_, _06661_, _06657_);
  not (_06663_, _06662_);
  nor (_06664_, _06602_, _06600_);
  nor (_06665_, _06664_, _06603_);
  and (_06666_, _06665_, _06663_);
  and (_06667_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_06668_, _06667_, _06611_);
  and (_06669_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_06670_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_06671_, _06670_, _06669_);
  nor (_06672_, _06671_, _06668_);
  nor (_06673_, _06665_, _06663_);
  nor (_06674_, _06673_, _06666_);
  and (_06675_, _06674_, _06672_);
  nor (_06676_, _06675_, _06666_);
  not (_06677_, _06676_);
  nor (_06678_, _06619_, _06617_);
  nor (_06679_, _06678_, _06620_);
  and (_06680_, _06679_, _06677_);
  nor (_06681_, _06679_, _06677_);
  nor (_06682_, _06681_, _06680_);
  and (_06683_, _06682_, _06668_);
  nor (_06684_, _06683_, _06680_);
  not (_06685_, _06684_);
  nor (_06686_, _06632_, _06630_);
  nor (_06687_, _06686_, _06633_);
  and (_06688_, _06687_, _06685_);
  nor (_06689_, _06640_, _06628_);
  nor (_06690_, _06689_, _06641_);
  and (_06691_, _06690_, _06688_);
  and (_06692_, _06645_, _06642_);
  nor (_06693_, _06692_, _06646_);
  and (_06694_, _06693_, _06691_);
  nor (_06695_, _06648_, _06646_);
  nor (_06696_, _06695_, _06649_);
  nor (_06697_, _06696_, _06694_);
  and (_06698_, _06696_, _06694_);
  not (_06699_, _06698_);
  and (_06700_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_06701_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_06702_, _06701_, _06700_);
  and (_06703_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_06704_, _06701_, _06700_);
  nor (_06705_, _06704_, _06702_);
  and (_06706_, _06705_, _06703_);
  nor (_06707_, _06706_, _06702_);
  not (_06708_, _06707_);
  nor (_06709_, _06660_, _06658_);
  nor (_06710_, _06709_, _06661_);
  and (_06711_, _06710_, _06708_);
  nor (_06712_, _06710_, _06708_);
  nor (_06713_, _06712_, _06711_);
  and (_06714_, _06713_, _06667_);
  nor (_06715_, _06714_, _06711_);
  not (_06716_, _06715_);
  nor (_06717_, _06674_, _06672_);
  nor (_06718_, _06717_, _06675_);
  and (_06719_, _06718_, _06716_);
  nor (_06720_, _06682_, _06668_);
  nor (_06721_, _06720_, _06683_);
  and (_06722_, _06721_, _06719_);
  nor (_06723_, _06687_, _06685_);
  nor (_06724_, _06723_, _06688_);
  and (_06725_, _06724_, _06722_);
  nor (_06726_, _06690_, _06688_);
  nor (_06727_, _06726_, _06691_);
  and (_06728_, _06727_, _06725_);
  nor (_06729_, _06693_, _06691_);
  nor (_06730_, _06729_, _06694_);
  and (_06731_, _06730_, _06728_);
  and (_06732_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_06733_, _06732_, _06701_);
  nor (_06734_, _06705_, _06703_);
  nor (_06735_, _06734_, _06706_);
  and (_06736_, _06735_, _06733_);
  nor (_06737_, _06713_, _06667_);
  nor (_06738_, _06737_, _06714_);
  and (_06739_, _06738_, _06736_);
  nor (_06740_, _06718_, _06716_);
  nor (_06741_, _06740_, _06719_);
  and (_06743_, _06741_, _06739_);
  nor (_06744_, _06721_, _06719_);
  nor (_06745_, _06744_, _06722_);
  and (_06746_, _06745_, _06743_);
  nor (_06747_, _06724_, _06722_);
  nor (_06748_, _06747_, _06725_);
  and (_06749_, _06748_, _06746_);
  nor (_06750_, _06727_, _06725_);
  nor (_06751_, _06750_, _06728_);
  and (_06752_, _06751_, _06749_);
  nor (_06753_, _06730_, _06728_);
  nor (_06754_, _06753_, _06731_);
  and (_06755_, _06754_, _06752_);
  nor (_06756_, _06755_, _06731_);
  and (_06757_, _06756_, _06699_);
  nor (_06758_, _06757_, _06697_);
  and (_06759_, _06758_, _06654_);
  nor (_06760_, _06759_, _06652_);
  not (_06761_, _06760_);
  and (_06762_, _06761_, _06596_);
  nor (_06763_, _06762_, _06594_);
  not (_06764_, _06763_);
  nor (_06765_, _06534_, _06532_);
  nor (_06766_, _06765_, _06535_);
  and (_06767_, _06766_, _06764_);
  nor (_06768_, _06767_, _06535_);
  not (_06769_, _06768_);
  and (_06770_, _06769_, _06470_);
  nor (_06771_, _06770_, _06468_);
  not (_06772_, _06771_);
  and (_06773_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_06774_, _06773_);
  nor (_06775_, _06774_, _06420_);
  nor (_06776_, _06775_, _06452_);
  nor (_06777_, _06458_, _06455_);
  nor (_06778_, _06777_, _06776_);
  and (_06779_, _06777_, _06776_);
  nor (_06780_, _06779_, _06778_);
  not (_06781_, _06780_);
  nor (_06782_, _06465_, _06462_);
  nor (_06783_, _06782_, _06781_);
  and (_06784_, _06782_, _06781_);
  nor (_06785_, _06784_, _06783_);
  and (_06786_, _06785_, _06772_);
  or (_06787_, _06778_, _06449_);
  or (_06788_, _06787_, _06783_);
  or (_06789_, _06788_, _06786_);
  or (_06790_, _06789_, _06277_);
  and (_06791_, _06790_, _02875_);
  and (_06792_, _06791_, _06276_);
  not (_06793_, _06241_);
  not (_06794_, _05338_);
  nor (_06795_, _05366_, _06794_);
  or (_06796_, _06795_, _06243_);
  and (_06797_, _06796_, _02874_);
  or (_06798_, _06797_, _06793_);
  or (_06799_, _06798_, _06792_);
  and (_06800_, _06799_, _06242_);
  or (_06801_, _06800_, _02855_);
  and (_06802_, _05490_, _04705_);
  or (_06803_, _06234_, _02856_);
  or (_06804_, _06803_, _06802_);
  and (_06805_, _06804_, _02851_);
  and (_06806_, _06805_, _06801_);
  and (_06807_, _03024_, _02520_);
  nor (_06808_, _05755_, _06235_);
  or (_06809_, _06808_, _06234_);
  and (_06810_, _06809_, _02576_);
  or (_06811_, _06810_, _06807_);
  or (_06812_, _06811_, _06806_);
  not (_06813_, _06807_);
  not (_06814_, \oc8051_golden_model_1.B [1]);
  nor (_06815_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor (_06816_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and (_06817_, _06816_, _06815_);
  and (_06818_, _06817_, _06814_);
  nor (_06819_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_06820_, \oc8051_golden_model_1.B [0]);
  and (_06821_, _06820_, \oc8051_golden_model_1.ACC [7]);
  and (_06822_, _06821_, _06819_);
  and (_06823_, _06822_, _06818_);
  and (_06824_, _06819_, _06818_);
  nor (_06825_, _06824_, _05768_);
  not (_06826_, \oc8051_golden_model_1.B [2]);
  not (_06827_, \oc8051_golden_model_1.B [3]);
  nor (_06828_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06829_, _06828_, _06815_);
  and (_06830_, _06829_, _06827_);
  and (_06831_, _06830_, _06826_);
  not (_06832_, _06831_);
  not (_06833_, \oc8051_golden_model_1.ACC [6]);
  and (_06834_, \oc8051_golden_model_1.B [0], _06833_);
  nor (_06835_, _06834_, _05768_);
  nor (_06836_, _06835_, _06814_);
  nor (_06837_, _06836_, _06832_);
  not (_06838_, _06837_);
  and (_06839_, _06838_, _06825_);
  nor (_06840_, _06839_, _06823_);
  and (_06841_, _06837_, \oc8051_golden_model_1.B [0]);
  nor (_06842_, _06841_, _06833_);
  and (_06843_, _06842_, _06814_);
  nor (_06844_, _06842_, _06814_);
  nor (_06845_, _06844_, _06843_);
  nor (_06846_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06847_, _06846_, _06471_);
  nor (_06848_, _06847_, \oc8051_golden_model_1.ACC [4]);
  nor (_06849_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_06850_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06851_, _06850_, _06820_);
  nor (_06852_, _06851_, _06849_);
  nor (_06853_, _06852_, _06848_);
  not (_06854_, _06853_);
  and (_06855_, _06854_, _06845_);
  not (_06856_, _06855_);
  nor (_06857_, _06840_, \oc8051_golden_model_1.B [2]);
  nor (_06858_, _06857_, _06843_);
  and (_06859_, _06858_, _06856_);
  and (_06860_, \oc8051_golden_model_1.B [2], _05768_);
  nor (_06861_, _06860_, \oc8051_golden_model_1.B [7]);
  and (_06862_, _06861_, _06817_);
  not (_06863_, _06862_);
  nor (_06864_, _06863_, _06859_);
  nor (_06865_, _06864_, _06840_);
  nor (_06866_, _06865_, _06823_);
  and (_06867_, _06829_, \oc8051_golden_model_1.ACC [7]);
  nor (_06868_, _06867_, _06830_);
  nor (_06869_, _06854_, _06845_);
  nor (_06870_, _06869_, _06855_);
  not (_06871_, _06870_);
  and (_06872_, _06871_, _06864_);
  nor (_06873_, _06864_, _06842_);
  nor (_06874_, _06873_, _06872_);
  and (_06875_, _06874_, _06826_);
  nor (_06876_, _06874_, _06826_);
  nor (_06877_, _06876_, _06875_);
  not (_06878_, _06877_);
  not (_06879_, \oc8051_golden_model_1.ACC [5]);
  nor (_06880_, _06864_, _06879_);
  and (_06881_, _06864_, _06847_);
  or (_06882_, _06881_, _06880_);
  and (_06883_, _06882_, _06814_);
  nor (_06884_, _06882_, _06814_);
  not (_06885_, \oc8051_golden_model_1.ACC [4]);
  and (_06886_, \oc8051_golden_model_1.B [0], _06885_);
  nor (_06887_, _06886_, _06884_);
  nor (_06888_, _06887_, _06883_);
  nor (_06889_, _06888_, _06878_);
  nor (_06890_, _06866_, \oc8051_golden_model_1.B [3]);
  nor (_06891_, _06890_, _06875_);
  not (_06892_, _06891_);
  nor (_06893_, _06892_, _06889_);
  nor (_06894_, _06893_, _06868_);
  nor (_06895_, _06894_, _06866_);
  nor (_06896_, _06895_, _06823_);
  not (_06897_, _06894_);
  and (_06898_, _06888_, _06878_);
  nor (_06899_, _06898_, _06889_);
  nor (_06900_, _06899_, _06897_);
  nor (_06901_, _06894_, _06874_);
  nor (_06902_, _06901_, _06900_);
  and (_06903_, _06902_, _06827_);
  nor (_06904_, _06902_, _06827_);
  nor (_06905_, _06904_, _06903_);
  not (_06906_, _06905_);
  nor (_06907_, _06894_, _06882_);
  nor (_06908_, _06884_, _06883_);
  and (_06909_, _06908_, _06886_);
  nor (_06910_, _06908_, _06886_);
  nor (_06911_, _06910_, _06909_);
  and (_06912_, _06911_, _06894_);
  or (_06913_, _06912_, _06907_);
  nor (_06914_, _06913_, \oc8051_golden_model_1.B [2]);
  and (_06915_, _06913_, \oc8051_golden_model_1.B [2]);
  nor (_06916_, _06894_, _06885_);
  nor (_06917_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06918_, _06917_, _06597_);
  and (_06919_, _06894_, _06918_);
  or (_06920_, _06919_, _06916_);
  and (_06921_, _06920_, _06814_);
  nor (_06922_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06923_, _06922_, _06655_);
  nor (_06924_, _06923_, \oc8051_golden_model_1.ACC [2]);
  nor (_06925_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06926_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06927_, _06926_, _06820_);
  nor (_06928_, _06927_, _06925_);
  nor (_06929_, _06928_, _06924_);
  not (_06930_, _06929_);
  nor (_06931_, _06920_, _06814_);
  nor (_06932_, _06931_, _06921_);
  and (_06933_, _06932_, _06930_);
  nor (_06934_, _06933_, _06921_);
  nor (_06935_, _06934_, _06915_);
  nor (_06936_, _06935_, _06914_);
  nor (_06937_, _06936_, _06906_);
  nor (_06938_, _06896_, \oc8051_golden_model_1.B [4]);
  nor (_06939_, _06938_, _06903_);
  not (_06940_, _06939_);
  nor (_06941_, _06940_, _06937_);
  not (_06942_, \oc8051_golden_model_1.B [5]);
  and (_06943_, _06828_, _06942_);
  and (_06944_, \oc8051_golden_model_1.B [4], _05768_);
  not (_06945_, _06944_);
  and (_06946_, _06945_, _06943_);
  not (_06947_, _06946_);
  nor (_06948_, _06947_, _06941_);
  nor (_06949_, _06948_, _06896_);
  nor (_06950_, _06949_, _06823_);
  not (_06951_, \oc8051_golden_model_1.B [4]);
  and (_06952_, _06936_, _06906_);
  nor (_06953_, _06952_, _06937_);
  not (_06954_, _06953_);
  and (_06955_, _06954_, _06948_);
  nor (_06956_, _06948_, _06902_);
  nor (_06957_, _06956_, _06955_);
  and (_06958_, _06957_, _06951_);
  nor (_06959_, _06957_, _06951_);
  nor (_06960_, _06959_, _06958_);
  not (_06961_, _06960_);
  nor (_06962_, _06948_, _06913_);
  nor (_06963_, _06915_, _06914_);
  and (_06964_, _06963_, _06934_);
  nor (_06965_, _06963_, _06934_);
  nor (_06966_, _06965_, _06964_);
  not (_06967_, _06966_);
  and (_06968_, _06967_, _06948_);
  nor (_06969_, _06968_, _06962_);
  nor (_06970_, _06969_, \oc8051_golden_model_1.B [3]);
  and (_06971_, _06969_, \oc8051_golden_model_1.B [3]);
  nor (_06972_, _06932_, _06930_);
  nor (_06973_, _06972_, _06933_);
  not (_06974_, _06973_);
  and (_06975_, _06974_, _06948_);
  nor (_06976_, _06948_, _06920_);
  nor (_06977_, _06976_, _06975_);
  and (_06978_, _06977_, _06826_);
  nor (_06979_, _06948_, _02701_);
  and (_06980_, _06948_, _06923_);
  or (_06981_, _06980_, _06979_);
  and (_06982_, _06981_, _06814_);
  nor (_06983_, _06981_, _06814_);
  not (_06984_, \oc8051_golden_model_1.ACC [2]);
  and (_06985_, \oc8051_golden_model_1.B [0], _06984_);
  nor (_06986_, _06985_, _06983_);
  nor (_06987_, _06986_, _06982_);
  nor (_06988_, _06977_, _06826_);
  nor (_06989_, _06988_, _06978_);
  not (_06990_, _06989_);
  nor (_06991_, _06990_, _06987_);
  nor (_06992_, _06991_, _06978_);
  nor (_06993_, _06992_, _06971_);
  nor (_06994_, _06993_, _06970_);
  nor (_06995_, _06994_, _06961_);
  nor (_06996_, _06950_, \oc8051_golden_model_1.B [5]);
  nor (_06997_, _06996_, _06958_);
  not (_06998_, _06997_);
  nor (_06999_, _06998_, _06995_);
  not (_07000_, _06999_);
  not (_07001_, _06828_);
  and (_07002_, \oc8051_golden_model_1.B [5], _05768_);
  nor (_07003_, _07002_, _07001_);
  and (_07004_, _07003_, _07000_);
  nor (_07005_, _07004_, _06950_);
  nor (_07006_, _07005_, _06823_);
  not (_07007_, _07004_);
  and (_07008_, _06994_, _06961_);
  nor (_07009_, _07008_, _06995_);
  nor (_07010_, _07009_, _07007_);
  nor (_07011_, _07004_, _06957_);
  nor (_07012_, _07011_, _07010_);
  and (_07013_, _07012_, _06942_);
  nor (_07014_, _07012_, _06942_);
  nor (_07015_, _07014_, _07013_);
  nor (_07016_, _06971_, _06970_);
  nor (_07017_, _07016_, _06992_);
  and (_07018_, _07016_, _06992_);
  or (_07019_, _07018_, _07017_);
  nor (_07020_, _07019_, _07007_);
  and (_07021_, _07007_, _06969_);
  nor (_07022_, _07021_, _07020_);
  and (_07023_, _07022_, _06951_);
  nor (_07024_, _07022_, _06951_);
  and (_07025_, _06990_, _06987_);
  nor (_07026_, _07025_, _06991_);
  nor (_07027_, _07026_, _07007_);
  nor (_07028_, _07004_, _06977_);
  nor (_07029_, _07028_, _07027_);
  and (_07030_, _07029_, _06827_);
  nor (_07031_, _06983_, _06982_);
  nor (_07032_, _07031_, _06985_);
  and (_07033_, _07031_, _06985_);
  or (_07034_, _07033_, _07032_);
  nor (_07035_, _07034_, _07007_);
  nor (_07036_, _07004_, _06981_);
  nor (_07037_, _07036_, _07035_);
  and (_07038_, _07037_, _06826_);
  nor (_07039_, _07037_, _06826_);
  nor (_07040_, _07004_, \oc8051_golden_model_1.ACC [2]);
  nor (_07041_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_07042_, _07041_, _06700_);
  nor (_07043_, _07007_, _07042_);
  nor (_07044_, _07043_, _07040_);
  and (_07045_, _07044_, _06814_);
  and (_07046_, \oc8051_golden_model_1.B [0], _02618_);
  not (_07047_, _07046_);
  nor (_07048_, _07044_, _06814_);
  nor (_07049_, _07048_, _07045_);
  and (_07050_, _07049_, _07047_);
  nor (_07051_, _07050_, _07045_);
  nor (_07052_, _07051_, _07039_);
  nor (_07053_, _07052_, _07038_);
  not (_07054_, _07053_);
  nor (_07055_, _07029_, _06827_);
  nor (_07056_, _07055_, _07030_);
  and (_07057_, _07056_, _07054_);
  nor (_07058_, _07057_, _07030_);
  nor (_07059_, _07058_, _07024_);
  nor (_07060_, _07059_, _07023_);
  not (_07061_, _07060_);
  and (_07062_, _07061_, _07015_);
  nor (_07063_, _07006_, \oc8051_golden_model_1.B [6]);
  or (_07064_, _07063_, _07013_);
  or (_07065_, _07064_, _07062_);
  not (_07066_, \oc8051_golden_model_1.B [6]);
  or (_07067_, _07066_, \oc8051_golden_model_1.ACC [7]);
  and (_07068_, _07067_, _06232_);
  and (_07069_, _07068_, _07065_);
  nor (_07070_, _07069_, _07006_);
  or (_07071_, _07070_, _06823_);
  nor (_07072_, _07071_, \oc8051_golden_model_1.B [7]);
  nor (_07073_, _07072_, _06773_);
  nor (_07074_, _07061_, _07015_);
  nor (_07075_, _07074_, _07062_);
  and (_07076_, _07075_, _07069_);
  not (_07077_, _07012_);
  nor (_07078_, _07069_, _07077_);
  nor (_07079_, _07078_, _07076_);
  and (_07080_, _07079_, \oc8051_golden_model_1.B [6]);
  not (_07081_, _07080_);
  nor (_07082_, _07081_, _07073_);
  nor (_07083_, _07039_, _07038_);
  and (_07084_, _07083_, _07051_);
  nor (_07085_, _07083_, _07051_);
  or (_07086_, _07085_, _07084_);
  and (_07087_, _07086_, _07069_);
  not (_07088_, _07037_);
  nor (_07089_, _07069_, _07088_);
  nor (_07090_, _07089_, _07087_);
  and (_07091_, _07090_, \oc8051_golden_model_1.B [3]);
  nor (_07092_, _07090_, \oc8051_golden_model_1.B [3]);
  nor (_07093_, _07092_, _07091_);
  nor (_07094_, _07049_, _07047_);
  nor (_07095_, _07094_, _07050_);
  and (_07096_, _07095_, _07069_);
  not (_07097_, _07044_);
  nor (_07098_, _07069_, _07097_);
  nor (_07099_, _07098_, _07096_);
  and (_07100_, _07099_, \oc8051_golden_model_1.B [2]);
  nor (_07101_, _07099_, \oc8051_golden_model_1.B [2]);
  nor (_07102_, _07101_, _07100_);
  and (_07103_, _07102_, _07093_);
  or (_07104_, _07069_, \oc8051_golden_model_1.ACC [1]);
  and (_07105_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07106_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07107_, _07106_, _07105_);
  nand (_07108_, _07069_, _07107_);
  and (_07109_, _07108_, _07104_);
  and (_07110_, _07109_, _06814_);
  nor (_07111_, _07109_, _06814_);
  and (_07112_, _06820_, \oc8051_golden_model_1.ACC [0]);
  not (_07113_, _07112_);
  nor (_07114_, _07113_, _07111_);
  nor (_07115_, _07114_, _07110_);
  and (_07116_, _07115_, _07103_);
  not (_07117_, _07116_);
  and (_07118_, _07100_, _07093_);
  nor (_07119_, _07118_, _07091_);
  and (_07120_, _07119_, _07117_);
  nor (_07121_, _07079_, \oc8051_golden_model_1.B [6]);
  nor (_07122_, _07121_, _07080_);
  not (_07123_, _07122_);
  nor (_07124_, _07123_, _07073_);
  nor (_07125_, _07056_, _07054_);
  nor (_07126_, _07125_, _07057_);
  and (_07127_, _07126_, _07069_);
  not (_07128_, _07029_);
  nor (_07129_, _07069_, _07128_);
  nor (_07130_, _07129_, _07127_);
  and (_07131_, _07130_, \oc8051_golden_model_1.B [4]);
  nor (_07132_, _07130_, \oc8051_golden_model_1.B [4]);
  nor (_07133_, _07132_, _07131_);
  nor (_07134_, _07024_, _07023_);
  nor (_07135_, _07134_, _07058_);
  and (_07136_, _07134_, _07058_);
  or (_07137_, _07136_, _07135_);
  and (_07138_, _07137_, _07069_);
  not (_07139_, _07022_);
  nor (_07140_, _07069_, _07139_);
  nor (_07141_, _07140_, _07138_);
  and (_07142_, _07141_, \oc8051_golden_model_1.B [5]);
  nor (_07143_, _07141_, \oc8051_golden_model_1.B [5]);
  nor (_07144_, _07143_, _07142_);
  and (_07145_, _07144_, _07133_);
  and (_07146_, _07145_, _07124_);
  not (_07147_, _07146_);
  nor (_07148_, _07147_, _07120_);
  and (_07149_, _07006_, \oc8051_golden_model_1.B [7]);
  and (_07150_, _07144_, _07131_);
  nor (_07151_, _07150_, _07142_);
  not (_07152_, _07151_);
  and (_07153_, _07152_, _07124_);
  or (_07154_, _07153_, _07149_);
  or (_07155_, _07154_, _07148_);
  nor (_07156_, _07155_, _07082_);
  and (_07157_, \oc8051_golden_model_1.B [0], _02549_);
  not (_07158_, _07157_);
  nor (_07159_, _07111_, _07110_);
  and (_07160_, _07159_, _07158_);
  and (_07161_, _07160_, _07113_);
  and (_07162_, _07161_, _07103_);
  and (_07163_, _07162_, _07146_);
  nor (_07164_, _07163_, _07156_);
  or (_07165_, _07164_, _06823_);
  and (_07166_, _07165_, _07071_);
  or (_07167_, _07166_, _06813_);
  and (_07168_, _07167_, _06812_);
  or (_07169_, _07168_, _03014_);
  and (_07170_, _05563_, _04705_);
  or (_07171_, _07170_, _06234_);
  or (_07172_, _07171_, _03884_);
  and (_07173_, _07172_, _05279_);
  and (_07174_, _07173_, _07169_);
  and (_07175_, _05314_, _04705_);
  or (_07176_, _07175_, _06234_);
  and (_07177_, _07176_, _03021_);
  or (_07178_, _07177_, _03130_);
  or (_07179_, _07178_, _07174_);
  and (_07180_, _05771_, _04705_);
  or (_07181_, _06234_, _03131_);
  or (_07182_, _07181_, _07180_);
  and (_07183_, _07182_, _05274_);
  and (_07184_, _07183_, _07179_);
  or (_07185_, _06234_, _04733_);
  and (_07186_, _07171_, _03020_);
  and (_07187_, _07186_, _07185_);
  or (_07188_, _07187_, _07184_);
  and (_07189_, _07188_, _03140_);
  and (_07190_, _06251_, _03139_);
  and (_07191_, _07190_, _07185_);
  or (_07192_, _07191_, _03036_);
  or (_07193_, _07192_, _07189_);
  nor (_07194_, _05312_, _06235_);
  or (_07195_, _06234_, _05781_);
  or (_07196_, _07195_, _07194_);
  and (_07197_, _07196_, _05786_);
  and (_07198_, _07197_, _07193_);
  nor (_07199_, _05770_, _06235_);
  or (_07200_, _07199_, _06234_);
  and (_07201_, _07200_, _03127_);
  or (_07202_, _07201_, _03166_);
  or (_07203_, _07202_, _07198_);
  or (_07204_, _06248_, _03563_);
  and (_07205_, _07204_, _02501_);
  and (_07206_, _07205_, _07203_);
  and (_07207_, _06245_, _02500_);
  or (_07208_, _07207_, _03174_);
  or (_07209_, _07208_, _07206_);
  and (_07210_, _05257_, _04705_);
  or (_07211_, _06234_, _03178_);
  or (_07212_, _07211_, _07210_);
  and (_07213_, _07212_, _34698_);
  and (_07214_, _07213_, _07209_);
  or (_07215_, _07214_, _06233_);
  and (_32485_, _07215_, _36029_);
  nor (_07216_, _34698_, _05768_);
  and (_07217_, _02854_, _02535_);
  and (_07218_, _04623_, _05768_);
  nor (_07219_, _04623_, _05768_);
  nor (_07220_, _07219_, _07218_);
  nor (_07221_, _04787_, _06833_);
  and (_07222_, _04787_, _06833_);
  nor (_07223_, _07222_, _07221_);
  nor (_07224_, _04896_, _06879_);
  and (_07225_, _04896_, _06879_);
  nor (_07226_, _07225_, _07224_);
  not (_07227_, _07226_);
  nor (_07228_, _05202_, _06885_);
  and (_07229_, _05202_, _06885_);
  nor (_07230_, _07229_, _07228_);
  and (_07231_, _04242_, _02701_);
  not (_07232_, _07231_);
  nor (_07233_, _04242_, _02701_);
  not (_07234_, _07233_);
  nor (_07235_, _04440_, _06984_);
  and (_07236_, _04440_, _06984_);
  nor (_07237_, _07236_, _07235_);
  not (_07238_, _07237_);
  and (_07239_, _04005_, \oc8051_golden_model_1.ACC [1]);
  and (_07240_, _04038_, _02618_);
  nor (_07241_, _07240_, _07239_);
  and (_07242_, _03817_, \oc8051_golden_model_1.ACC [0]);
  and (_07243_, _07242_, _07241_);
  nor (_07244_, _07243_, _07239_);
  nor (_07245_, _07244_, _07238_);
  nor (_07246_, _07245_, _07235_);
  nand (_07247_, _07246_, _07234_);
  and (_07248_, _07247_, _07232_);
  and (_07249_, _07248_, _07230_);
  nor (_07250_, _07249_, _07228_);
  nor (_07251_, _07250_, _07227_);
  or (_07252_, _07251_, _07224_);
  and (_07253_, _07252_, _07223_);
  nor (_07254_, _07253_, _07221_);
  nor (_07255_, _07254_, _07220_);
  and (_07256_, _07254_, _07220_);
  or (_07257_, _07256_, _07255_);
  and (_07258_, _02535_, _02432_);
  not (_07259_, _07258_);
  or (_07260_, _07259_, _07257_);
  and (_07261_, _02845_, _02537_);
  nor (_07262_, _07261_, _03360_);
  not (_07263_, _07262_);
  nand (_07264_, _07263_, _07218_);
  not (_07265_, _03513_);
  and (_07266_, _05490_, \oc8051_golden_model_1.ACC [7]);
  or (_07267_, _07266_, _07265_);
  nor (_07268_, _04712_, _05768_);
  and (_07269_, _05314_, _04712_);
  nor (_07270_, _07269_, _07268_);
  nand (_07271_, _07270_, _03021_);
  not (_07272_, _04712_);
  nor (_07273_, _07272_, _04623_);
  nor (_07274_, _07273_, _07268_);
  nand (_07275_, _07274_, _06793_);
  and (_07276_, _03024_, _02577_);
  not (_07277_, _07276_);
  and (_07278_, _04630_, \oc8051_golden_model_1.PSW [7]);
  and (_07279_, _07278_, _04636_);
  and (_07280_, _07279_, _04697_);
  and (_07281_, _07280_, _04352_);
  nor (_07282_, _07281_, _02858_);
  and (_07283_, _07280_, _02933_);
  nor (_07284_, _07283_, _07282_);
  and (_07285_, _07284_, \oc8051_golden_model_1.ACC [7]);
  nor (_07286_, _07284_, \oc8051_golden_model_1.ACC [7]);
  nor (_07287_, _07286_, _07285_);
  not (_07288_, _07287_);
  nor (_07289_, _07280_, _04352_);
  nor (_07290_, _07289_, _07281_);
  nor (_07291_, _07290_, _06833_);
  and (_07292_, _07290_, _06833_);
  nor (_07293_, _07291_, _07292_);
  and (_07294_, _07279_, _04662_);
  nor (_07295_, _07294_, _04669_);
  nor (_07296_, _07295_, _07280_);
  nor (_07297_, _07296_, _06879_);
  and (_07298_, _07296_, _06879_);
  nor (_07299_, _07298_, _07297_);
  nor (_07300_, _07279_, _04662_);
  nor (_07301_, _07300_, _07294_);
  nor (_07302_, _07301_, _06885_);
  and (_07303_, _07301_, _06885_);
  nor (_07304_, _07303_, _07302_);
  and (_07305_, _07304_, _07299_);
  nor (_07306_, _05365_, _02934_);
  nor (_07307_, _07306_, _07279_);
  and (_07308_, _07307_, _02701_);
  nor (_07309_, _07307_, _02701_);
  nor (_07310_, _07278_, _03261_);
  nor (_07311_, _07310_, _05365_);
  nor (_07312_, _07311_, _06984_);
  nor (_07313_, _07312_, _07309_);
  or (_07314_, _07313_, _07308_);
  nor (_07315_, _07308_, _07309_);
  and (_07316_, _07311_, _06984_);
  nor (_07317_, _07316_, _07312_);
  and (_07318_, _07317_, _07315_);
  not (_07319_, \oc8051_golden_model_1.PSW [7]);
  nor (_07320_, _02832_, _07319_);
  nor (_07321_, _07320_, _03672_);
  nor (_07322_, _07321_, _07278_);
  and (_07323_, _07322_, _02618_);
  nor (_07324_, _07322_, _02618_);
  nor (_07325_, _02832_, \oc8051_golden_model_1.PSW [7]);
  and (_07326_, _02832_, \oc8051_golden_model_1.PSW [7]);
  nor (_07327_, _07326_, _07325_);
  or (_07328_, _07327_, \oc8051_golden_model_1.ACC [0]);
  nor (_07329_, _07328_, _07324_);
  nor (_07330_, _07329_, _07323_);
  nand (_07331_, _07330_, _07318_);
  and (_07332_, _07331_, _07314_);
  not (_07333_, _07332_);
  and (_07334_, _07333_, _07305_);
  nor (_07335_, _07302_, _07297_);
  nor (_07336_, _07335_, _07298_);
  or (_07337_, _07336_, _07334_);
  and (_07338_, _07337_, _07293_);
  or (_07339_, _07338_, _07291_);
  and (_07340_, _07339_, _07288_);
  nor (_07341_, _07339_, _07288_);
  or (_07342_, _07341_, _07340_);
  or (_07343_, _07342_, _07277_);
  not (_07344_, _03441_);
  and (_07345_, _06184_, \oc8051_golden_model_1.PSW [7]);
  nor (_07346_, _07345_, _05490_);
  and (_07347_, _06185_, \oc8051_golden_model_1.PSW [7]);
  nor (_07348_, _07347_, _07346_);
  nor (_07349_, _07348_, _05768_);
  and (_07350_, _07348_, _05768_);
  nor (_07351_, _07350_, _07349_);
  not (_07352_, _07351_);
  and (_07353_, _06179_, _06181_);
  and (_07354_, _07353_, \oc8051_golden_model_1.PSW [7]);
  and (_07355_, _07354_, _06180_);
  nor (_07356_, _07355_, _05847_);
  nor (_07357_, _07356_, _07345_);
  nor (_07358_, _07357_, _06833_);
  and (_07359_, _07357_, _06833_);
  nor (_07360_, _07354_, _06180_);
  nor (_07361_, _07360_, _07355_);
  and (_07362_, _07361_, _06879_);
  nor (_07363_, _07361_, _06879_);
  and (_07364_, _06175_, \oc8051_golden_model_1.PSW [7]);
  and (_07365_, _07364_, _06178_);
  nor (_07366_, _07365_, _06181_);
  nor (_07367_, _07366_, _07354_);
  nor (_07368_, _07367_, _06885_);
  nor (_07369_, _07368_, _07363_);
  nor (_07370_, _07369_, _07362_);
  nor (_07371_, _07363_, _07362_);
  and (_07372_, _07367_, _06885_);
  nor (_07373_, _07372_, _07368_);
  and (_07374_, _07373_, _07371_);
  not (_07375_, _07374_);
  and (_07376_, _06175_, _06177_);
  and (_07377_, _07376_, \oc8051_golden_model_1.PSW [7]);
  nor (_07378_, _07377_, _06176_);
  nor (_07379_, _07378_, _07365_);
  nor (_07380_, _07379_, _02701_);
  and (_07381_, _07379_, _02701_);
  nor (_07382_, _07381_, _07380_);
  nor (_07383_, _07364_, _06177_);
  nor (_07384_, _07383_, _07377_);
  nor (_07385_, _07384_, _06984_);
  and (_07386_, _07384_, _06984_);
  nor (_07387_, _07386_, _07385_);
  and (_07388_, _07387_, _07382_);
  and (_07389_, _06174_, \oc8051_golden_model_1.PSW [7]);
  nor (_07390_, _07389_, _06173_);
  nor (_07391_, _07390_, _07364_);
  and (_07392_, _07391_, _02618_);
  nor (_07393_, _07391_, _02618_);
  and (_07394_, _05938_, _07319_);
  nor (_07395_, _07394_, _07389_);
  nor (_07396_, _07395_, _02549_);
  nor (_07397_, _07396_, _07393_);
  nor (_07398_, _07397_, _07392_);
  not (_07399_, _07398_);
  and (_07400_, _07399_, _07388_);
  not (_07401_, _07400_);
  and (_07402_, _07386_, _07382_);
  nor (_07403_, _07402_, _07381_);
  and (_07404_, _07403_, _07401_);
  nor (_07405_, _07392_, _07393_);
  and (_07406_, _07395_, _02549_);
  nor (_07407_, _07396_, _07406_);
  and (_07408_, _07407_, _07405_);
  and (_07409_, _07408_, _07388_);
  nor (_07410_, _07409_, _07404_);
  nor (_07411_, _07410_, _07375_);
  nor (_07412_, _07411_, _07370_);
  nor (_07413_, _07412_, _07359_);
  or (_07414_, _07413_, _07358_);
  and (_07415_, _07414_, _07352_);
  nor (_07416_, _07414_, _07352_);
  or (_07417_, _07416_, _07415_);
  or (_07418_, _07417_, _07344_);
  nor (_07419_, _02975_, _03316_);
  not (_07420_, _07419_);
  nor (_07421_, _03011_, _03316_);
  not (_07422_, _07421_);
  and (_07423_, _02864_, _02577_);
  nor (_07424_, _07423_, _03444_);
  and (_07425_, _07424_, _07422_);
  and (_07426_, _07425_, _07420_);
  not (_07427_, _07426_);
  not (_07428_, _03336_);
  and (_07429_, _04108_, _07428_);
  and (_07430_, _07429_, _04033_);
  not (_07431_, _07430_);
  nand (_07432_, _07431_, _04623_);
  not (_07433_, _02954_);
  nor (_07434_, _05528_, _07433_);
  and (_07435_, _02854_, _02953_);
  not (_07436_, _07435_);
  or (_07437_, _05490_, _07436_);
  and (_07438_, _02842_, _02953_);
  not (_07439_, _07438_);
  and (_07440_, _07439_, _03324_);
  nor (_07441_, _07440_, _04623_);
  and (_07442_, _03024_, _03383_);
  nor (_07443_, _07442_, \oc8051_golden_model_1.ACC [7]);
  and (_07444_, _07442_, \oc8051_golden_model_1.ACC [7]);
  nor (_07445_, _07444_, _07443_);
  nand (_07446_, _07445_, _07440_);
  nand (_07447_, _07446_, _07436_);
  or (_07448_, _07447_, _07441_);
  and (_07449_, _07448_, _07433_);
  and (_07450_, _07449_, _07437_);
  or (_07451_, _07450_, _07434_);
  and (_07452_, _03024_, _02953_);
  nor (_07453_, _07452_, _02952_);
  and (_07454_, _07453_, _07451_);
  and (_07455_, _03024_, _02890_);
  and (_07456_, _05502_, _04712_);
  nor (_07457_, _07456_, _07268_);
  nor (_07458_, _07457_, _03821_);
  or (_07459_, _07458_, _07455_);
  or (_07460_, _07459_, _07454_);
  nor (_07461_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07462_, _07461_, _02701_);
  and (_07463_, _07462_, _06850_);
  and (_07464_, _07463_, \oc8051_golden_model_1.ACC [6]);
  and (_07465_, _07464_, \oc8051_golden_model_1.ACC [7]);
  nor (_07466_, _07464_, \oc8051_golden_model_1.ACC [7]);
  nor (_07467_, _07466_, _07465_);
  and (_07468_, _07462_, \oc8051_golden_model_1.ACC [4]);
  nor (_07469_, _07468_, \oc8051_golden_model_1.ACC [5]);
  nor (_07470_, _07469_, _07463_);
  nor (_07471_, _07463_, \oc8051_golden_model_1.ACC [6]);
  nor (_07472_, _07471_, _07464_);
  nor (_07473_, _07472_, _07470_);
  not (_07474_, _07473_);
  and (_07475_, _07474_, _07467_);
  nor (_07476_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_07477_, _07476_, _07473_);
  nor (_07478_, _07477_, _07467_);
  nor (_07479_, _07478_, _07475_);
  not (_07480_, _07479_);
  nand (_07481_, _07480_, _07455_);
  and (_07482_, _07481_, _02951_);
  and (_07483_, _07482_, _07460_);
  nor (_07484_, _05331_, _05768_);
  and (_07485_, _05385_, _05331_);
  nor (_07486_, _07485_, _07484_);
  nor (_07487_, _07486_, _02892_);
  nor (_07488_, _07274_, _03327_);
  or (_07489_, _07488_, _07431_);
  or (_07490_, _07489_, _07487_);
  or (_07491_, _07490_, _07483_);
  and (_07492_, _07491_, _07432_);
  or (_07493_, _07492_, _03413_);
  or (_07494_, _05490_, _03849_);
  and (_07495_, _07494_, _02959_);
  and (_07496_, _07495_, _07493_);
  and (_07497_, _03024_, _02885_);
  nor (_07498_, _05528_, _02959_);
  or (_07499_, _07498_, _07497_);
  or (_07500_, _07499_, _07496_);
  nand (_07501_, _07497_, _02701_);
  and (_07502_, _07501_, _07500_);
  or (_07503_, _07502_, _02887_);
  and (_07504_, _05380_, _05331_);
  nor (_07505_, _07504_, _07484_);
  nand (_07506_, _07505_, _02887_);
  and (_07507_, _07506_, _02881_);
  and (_07508_, _07507_, _07503_);
  and (_07509_, _07485_, _05533_);
  nor (_07510_, _07509_, _07484_);
  nor (_07511_, _07510_, _02881_);
  or (_07512_, _07511_, _06271_);
  or (_07513_, _07512_, _07508_);
  nor (_07514_, _06751_, _06749_);
  nor (_07515_, _07514_, _06752_);
  or (_07516_, _07515_, _06277_);
  and (_07517_, _07516_, _07513_);
  or (_07518_, _07517_, _07427_);
  and (_07519_, _06166_, \oc8051_golden_model_1.PSW [7]);
  nor (_07520_, _07519_, _04623_);
  and (_07521_, _07519_, _04623_);
  nor (_07522_, _07521_, _07520_);
  and (_07523_, _07522_, \oc8051_golden_model_1.ACC [7]);
  nor (_07524_, _07522_, \oc8051_golden_model_1.ACC [7]);
  nor (_07525_, _07524_, _07523_);
  and (_07526_, _06165_, \oc8051_golden_model_1.PSW [7]);
  nor (_07527_, _07526_, _06158_);
  nor (_07528_, _07527_, _07519_);
  nor (_07529_, _07528_, _06833_);
  and (_07530_, _07528_, _06833_);
  and (_07531_, _06164_, \oc8051_golden_model_1.PSW [7]);
  nor (_07532_, _07531_, _06159_);
  nor (_07533_, _07532_, _07526_);
  and (_07534_, _07533_, _06879_);
  nor (_07535_, _07533_, _06879_);
  nor (_07536_, _07535_, _07534_);
  and (_07537_, _06161_, \oc8051_golden_model_1.PSW [7]);
  and (_07538_, _07537_, _06162_);
  nor (_07539_, _07538_, _06160_);
  nor (_07540_, _07539_, _07531_);
  nor (_07541_, _07540_, _06885_);
  and (_07542_, _07540_, _06885_);
  nor (_07543_, _07542_, _07541_);
  and (_07544_, _07543_, _07536_);
  not (_07545_, _07544_);
  and (_07546_, _06161_, _04441_);
  and (_07547_, _07546_, \oc8051_golden_model_1.PSW [7]);
  nor (_07548_, _07547_, _05412_);
  nor (_07549_, _07548_, _07538_);
  nor (_07550_, _07549_, _02701_);
  and (_07551_, _07549_, _02701_);
  nor (_07552_, _07551_, _07550_);
  nor (_07553_, _07537_, _04441_);
  nor (_07554_, _07553_, _07547_);
  nor (_07555_, _07554_, _06984_);
  and (_07556_, _07554_, _06984_);
  nor (_07557_, _07556_, _07555_);
  and (_07558_, _07557_, _07552_);
  and (_07559_, _03817_, \oc8051_golden_model_1.PSW [7]);
  nor (_07560_, _07559_, _04005_);
  nor (_07561_, _07560_, _07537_);
  and (_07562_, _07561_, _02618_);
  nor (_07563_, _07561_, _02618_);
  nor (_07564_, _03817_, \oc8051_golden_model_1.PSW [7]);
  nor (_07565_, _07564_, _07559_);
  nor (_07566_, _07565_, _02549_);
  nor (_07567_, _07566_, _07563_);
  nor (_07568_, _07567_, _07562_);
  not (_07569_, _07568_);
  and (_07570_, _07569_, _07558_);
  not (_07571_, _07570_);
  and (_07572_, _07556_, _07552_);
  nor (_07573_, _07572_, _07551_);
  and (_07574_, _07573_, _07571_);
  nor (_07575_, _07562_, _07563_);
  and (_07576_, _07565_, _02549_);
  nor (_07577_, _07566_, _07576_);
  and (_07578_, _07577_, _07575_);
  and (_07579_, _07578_, _07558_);
  nor (_07580_, _07579_, _07574_);
  nor (_07581_, _07580_, _07545_);
  not (_07582_, _07581_);
  and (_07583_, _07541_, _07536_);
  nor (_07584_, _07583_, _07535_);
  and (_07585_, _07584_, _07582_);
  nor (_07586_, _07585_, _07530_);
  or (_07587_, _07586_, _07529_);
  nor (_07588_, _07587_, _07525_);
  and (_07589_, _07587_, _07525_);
  nor (_07590_, _07589_, _07588_);
  or (_07591_, _07590_, _07426_);
  and (_07592_, _07591_, _07518_);
  or (_07593_, _07592_, _03441_);
  and (_07594_, _07593_, _02997_);
  and (_07595_, _07594_, _07418_);
  nor (_07596_, _07276_, _02992_);
  not (_07597_, _07596_);
  and (_07598_, _05528_, _05768_);
  nor (_07599_, _05528_, _05768_);
  nor (_07600_, _07599_, _07598_);
  and (_07601_, _04722_, \oc8051_golden_model_1.P2INREG [6]);
  and (_07602_, _04724_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_07603_, _07602_, _07601_);
  and (_07604_, _04716_, \oc8051_golden_model_1.P0INREG [6]);
  and (_07605_, _04719_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_07606_, _07605_, _07604_);
  and (_07607_, _07606_, _07603_);
  and (_07608_, _07607_, _04794_);
  and (_07609_, _07608_, _04835_);
  and (_07610_, _07609_, _04788_);
  and (_07611_, _07610_, \oc8051_golden_model_1.ACC [6]);
  nor (_07612_, _07610_, \oc8051_golden_model_1.ACC [6]);
  nor (_07613_, _07612_, _07611_);
  and (_07614_, _04722_, \oc8051_golden_model_1.P2INREG [5]);
  and (_07615_, _04724_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_07616_, _07615_, _07614_);
  and (_07617_, _04716_, \oc8051_golden_model_1.P0INREG [5]);
  and (_07618_, _04719_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_07619_, _07618_, _07617_);
  and (_07620_, _07619_, _07616_);
  and (_07621_, _07620_, _04932_);
  and (_07622_, _07621_, _04923_);
  and (_07623_, _07622_, _04917_);
  and (_07624_, _07623_, _04897_);
  and (_07625_, _07624_, \oc8051_golden_model_1.ACC [5]);
  nor (_07626_, _07624_, \oc8051_golden_model_1.ACC [5]);
  and (_07627_, _04716_, \oc8051_golden_model_1.P0INREG [4]);
  not (_07628_, _07627_);
  and (_07629_, _07628_, _05233_);
  and (_07630_, _04719_, \oc8051_golden_model_1.P1INREG [4]);
  not (_07631_, _07630_);
  and (_07632_, _04722_, \oc8051_golden_model_1.P2INREG [4]);
  and (_07633_, _04724_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_07634_, _07633_, _07632_);
  and (_07635_, _07634_, _05241_);
  and (_07636_, _07635_, _07631_);
  and (_07637_, _07636_, _05237_);
  and (_07638_, _07637_, _07629_);
  and (_07639_, _07638_, _05221_);
  and (_07640_, _07639_, _05203_);
  and (_07641_, _07640_, \oc8051_golden_model_1.ACC [4]);
  and (_07642_, _04722_, \oc8051_golden_model_1.P2INREG [3]);
  and (_07643_, _04724_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_07644_, _07643_, _07642_);
  and (_07645_, _04716_, \oc8051_golden_model_1.P0INREG [3]);
  and (_07646_, _04719_, \oc8051_golden_model_1.P1INREG [3]);
  nor (_07647_, _07646_, _07645_);
  and (_07648_, _07647_, _07644_);
  and (_07649_, _07648_, _04952_);
  and (_07650_, _07649_, _04993_);
  and (_07651_, _07650_, _04945_);
  and (_07652_, _07651_, \oc8051_golden_model_1.ACC [3]);
  nor (_07653_, _07651_, \oc8051_golden_model_1.ACC [3]);
  not (_07654_, _05115_);
  nor (_07655_, _05119_, _05116_);
  and (_07656_, _07655_, _05127_);
  and (_07657_, _07656_, _07654_);
  and (_07658_, _07657_, _05139_);
  and (_07659_, _05124_, _05103_);
  and (_07660_, _04722_, \oc8051_golden_model_1.P2INREG [2]);
  and (_07661_, _04724_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_07662_, _07661_, _07660_);
  and (_07663_, _04719_, \oc8051_golden_model_1.P1INREG [2]);
  and (_07664_, _04716_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_07665_, _07664_, _07663_);
  and (_07666_, _07665_, _07662_);
  and (_07667_, _07666_, _05114_);
  and (_07668_, _07667_, _07659_);
  and (_07669_, _07668_, _07658_);
  and (_07670_, _07669_, _05097_);
  and (_07671_, _07670_, \oc8051_golden_model_1.ACC [2]);
  and (_07672_, _04722_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07673_, _04724_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_07674_, _07673_, _07672_);
  and (_07675_, _04716_, \oc8051_golden_model_1.P0INREG [1]);
  and (_07676_, _04719_, \oc8051_golden_model_1.P1INREG [1]);
  nor (_07677_, _07676_, _07675_);
  and (_07678_, _07677_, _07674_);
  and (_07679_, _07678_, _05051_);
  and (_07680_, _07679_, _05093_);
  and (_07681_, _07680_, _05045_);
  and (_07682_, _07681_, \oc8051_golden_model_1.ACC [1]);
  nor (_07683_, _07681_, \oc8051_golden_model_1.ACC [1]);
  not (_07684_, _05015_);
  nor (_07685_, _05019_, _05016_);
  and (_07686_, _07685_, _05027_);
  and (_07687_, _07686_, _07684_);
  and (_07688_, _07687_, _05041_);
  and (_07689_, _05024_, _05003_);
  and (_07690_, _04722_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07691_, _04724_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07692_, _07691_, _07690_);
  and (_07693_, _04719_, \oc8051_golden_model_1.P1INREG [0]);
  and (_07694_, _04716_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_07695_, _07694_, _07693_);
  and (_07696_, _07695_, _07692_);
  and (_07697_, _07696_, _05014_);
  and (_07698_, _07697_, _07689_);
  and (_07699_, _07698_, _07688_);
  and (_07700_, _07699_, _04997_);
  nor (_07701_, _07700_, \oc8051_golden_model_1.ACC [0]);
  nor (_07702_, _07701_, _07683_);
  or (_07703_, _07702_, _07682_);
  nor (_07704_, _07670_, \oc8051_golden_model_1.ACC [2]);
  nor (_07705_, _07704_, _07671_);
  and (_07706_, _07705_, _07703_);
  nor (_07707_, _07706_, _07671_);
  nor (_07708_, _07707_, _07653_);
  or (_07709_, _07708_, _07652_);
  nor (_07710_, _07640_, \oc8051_golden_model_1.ACC [4]);
  nor (_07711_, _07710_, _07641_);
  and (_07712_, _07711_, _07709_);
  nor (_07713_, _07712_, _07641_);
  nor (_07714_, _07713_, _07626_);
  or (_07715_, _07714_, _07625_);
  and (_07716_, _07715_, _07613_);
  nor (_07717_, _07716_, _07611_);
  and (_07718_, _07717_, _07600_);
  nor (_07719_, _07717_, _07600_);
  nor (_07720_, _07719_, _07718_);
  not (_07721_, _07720_);
  nor (_07722_, _07715_, _07613_);
  nor (_07723_, _07722_, _07716_);
  nor (_07724_, _07625_, _07626_);
  nor (_07725_, _07724_, _07713_);
  and (_07726_, _07724_, _07713_);
  or (_07727_, _07726_, _07725_);
  nor (_07728_, _07711_, _07709_);
  nor (_07729_, _07728_, _07712_);
  nor (_07730_, _07652_, _07653_);
  and (_07731_, _07730_, _07705_);
  nor (_07732_, _07682_, _07683_);
  and (_07733_, _07700_, \oc8051_golden_model_1.ACC [0]);
  nor (_07734_, _07733_, _07701_);
  and (_07735_, _07734_, _07732_);
  and (_07736_, _07735_, _07731_);
  and (_07737_, _07736_, \oc8051_golden_model_1.PSW [7]);
  not (_07738_, _07737_);
  nor (_07739_, _07738_, _07729_);
  not (_07740_, _07739_);
  nor (_07741_, _07740_, _07727_);
  not (_07742_, _07741_);
  nor (_07743_, _07742_, _07723_);
  nor (_07744_, _07743_, _07721_);
  and (_07745_, _07743_, _07721_);
  or (_07746_, _07745_, _07276_);
  or (_07747_, _07746_, _07744_);
  and (_07748_, _07747_, _07597_);
  or (_07749_, _07748_, _07595_);
  and (_07750_, _07749_, _07343_);
  or (_07751_, _07750_, _02585_);
  or (_07752_, _02768_, _02586_);
  and (_07753_, _07752_, _02875_);
  and (_07754_, _07753_, _07751_);
  not (_07755_, _05331_);
  nor (_07756_, _05366_, _07755_);
  nor (_07757_, _07756_, _07484_);
  nor (_07758_, _07757_, _02875_);
  or (_07759_, _07758_, _06793_);
  or (_07760_, _07759_, _07754_);
  and (_07761_, _07760_, _07275_);
  or (_07762_, _07761_, _02855_);
  and (_07763_, _05490_, _04712_);
  or (_07764_, _07763_, _07268_);
  or (_07765_, _07764_, _02856_);
  and (_07766_, _07765_, _02851_);
  and (_07767_, _07766_, _07762_);
  nor (_07768_, _05755_, _07272_);
  nor (_07769_, _07768_, _07268_);
  nor (_07770_, _07769_, _02851_);
  or (_07771_, _07770_, _06807_);
  or (_07772_, _07771_, _07767_);
  and (_07773_, \oc8051_golden_model_1.B [0], _05768_);
  not (_07774_, _07773_);
  and (_07775_, _07774_, _06824_);
  or (_07776_, _07775_, _06813_);
  and (_07777_, _07776_, _07772_);
  and (_07778_, _07777_, _02584_);
  and (_07779_, _02768_, _02548_);
  or (_07780_, _07779_, _03014_);
  or (_07781_, _07780_, _07778_);
  and (_07782_, _03024_, _02516_);
  not (_07783_, _07782_);
  and (_07784_, _05563_, _04712_);
  nor (_07785_, _07784_, _07268_);
  nand (_07786_, _07785_, _03014_);
  and (_07787_, _07786_, _07783_);
  and (_07788_, _07787_, _07781_);
  and (_07789_, _07782_, _02768_);
  not (_07790_, _02511_);
  nor (_07791_, _02975_, _07790_);
  not (_07792_, _07791_);
  nor (_07793_, _03011_, _07790_);
  and (_07794_, _02862_, _02511_);
  and (_07795_, _02864_, _02511_);
  or (_07796_, _07795_, _07794_);
  nor (_07797_, _07796_, _07793_);
  and (_07798_, _07797_, _07792_);
  not (_07799_, _07798_);
  or (_07800_, _07799_, _07789_);
  or (_07801_, _07800_, _07788_);
  and (_07802_, _02854_, _02511_);
  not (_07803_, _07802_);
  or (_07804_, _07798_, _07220_);
  and (_07805_, _07804_, _07803_);
  and (_07806_, _07805_, _07801_);
  nor (_07807_, _05490_, \oc8051_golden_model_1.ACC [7]);
  nor (_07808_, _07807_, _07266_);
  and (_07809_, _07808_, _07802_);
  or (_07810_, _07809_, _03132_);
  or (_07811_, _07810_, _07806_);
  and (_07812_, _03024_, _02511_);
  not (_07813_, _07812_);
  not (_07814_, _03132_);
  or (_07815_, _05771_, _07814_);
  and (_07816_, _07815_, _07813_);
  and (_07817_, _07816_, _07811_);
  nor (_07818_, _02768_, \oc8051_golden_model_1.ACC [7]);
  and (_07819_, _02768_, \oc8051_golden_model_1.ACC [7]);
  nor (_07820_, _07819_, _07818_);
  and (_07821_, _07812_, _07820_);
  or (_07822_, _07821_, _03021_);
  or (_07823_, _07822_, _07817_);
  and (_07824_, _07823_, _07271_);
  or (_07825_, _07824_, _03130_);
  or (_07826_, _07268_, _03131_);
  and (_07827_, _02532_, _02432_);
  not (_07828_, _07827_);
  and (_07829_, _07828_, _07826_);
  and (_07830_, _07829_, _07825_);
  and (_07831_, _07827_, _07219_);
  or (_07832_, _07831_, _03513_);
  or (_07833_, _07832_, _07830_);
  and (_07834_, _07833_, _07267_);
  or (_07835_, _07834_, _03141_);
  and (_07836_, _03024_, _02532_);
  not (_07837_, _07836_);
  not (_07838_, _03141_);
  or (_07839_, _05769_, _07838_);
  and (_07840_, _07839_, _07837_);
  and (_07841_, _07840_, _07835_);
  and (_07842_, _07836_, _07819_);
  or (_07843_, _07842_, _07841_);
  and (_07844_, _07843_, _05274_);
  or (_07845_, _07785_, _05770_);
  nor (_07846_, _07845_, _05274_);
  or (_07847_, _07846_, _07263_);
  or (_07848_, _07847_, _07844_);
  and (_07849_, _07848_, _07264_);
  and (_07850_, _02864_, _02537_);
  nor (_07851_, _07850_, _03523_);
  not (_07852_, _07851_);
  or (_07853_, _07852_, _07849_);
  not (_07854_, _03525_);
  nand (_07855_, _07852_, _07218_);
  and (_07856_, _07855_, _07854_);
  and (_07857_, _07856_, _07853_);
  and (_07858_, _02854_, _02537_);
  nor (_07859_, _07218_, _07854_);
  or (_07860_, _07859_, _07858_);
  or (_07861_, _07860_, _07857_);
  nand (_07862_, _07807_, _07858_);
  and (_07863_, _07862_, _03126_);
  and (_07864_, _07863_, _07861_);
  and (_07865_, _03024_, _02537_);
  nor (_07866_, _07865_, _03125_);
  not (_07867_, _07866_);
  not (_07868_, _07865_);
  nand (_07869_, _07868_, _05770_);
  and (_07870_, _07869_, _07867_);
  or (_07871_, _07870_, _07864_);
  nand (_07872_, _07865_, _07818_);
  and (_07873_, _07872_, _05781_);
  and (_07874_, _07873_, _07871_);
  nor (_07875_, _05312_, _07272_);
  nor (_07876_, _07875_, _07268_);
  nor (_07877_, _07876_, _05781_);
  and (_07878_, _02845_, _02530_);
  nor (_07879_, _07878_, _03535_);
  nor (_07880_, _02975_, _03537_);
  nor (_07881_, _07880_, _03310_);
  and (_07882_, _07881_, _07879_);
  not (_07883_, _07882_);
  or (_07884_, _07883_, _07877_);
  or (_07885_, _07884_, _07874_);
  and (_07886_, _02862_, _02530_);
  and (_07887_, _02864_, _02530_);
  nor (_07888_, _07887_, _07886_);
  and (_07889_, _07888_, _07882_);
  and (_07890_, _07528_, \oc8051_golden_model_1.ACC [6]);
  nor (_07891_, _07529_, _07530_);
  and (_07892_, _07533_, \oc8051_golden_model_1.ACC [5]);
  and (_07893_, _07540_, \oc8051_golden_model_1.ACC [4]);
  and (_07894_, _07549_, \oc8051_golden_model_1.ACC [3]);
  and (_07895_, _07554_, \oc8051_golden_model_1.ACC [2]);
  and (_07896_, _07561_, \oc8051_golden_model_1.ACC [1]);
  and (_07897_, _07565_, \oc8051_golden_model_1.ACC [0]);
  not (_07898_, _07897_);
  nor (_07899_, _07898_, _07575_);
  nor (_07900_, _07899_, _07896_);
  nor (_07901_, _07900_, _07557_);
  nor (_07902_, _07901_, _07895_);
  nor (_07903_, _07902_, _07552_);
  nor (_07904_, _07903_, _07894_);
  nor (_07905_, _07904_, _07543_);
  nor (_07906_, _07905_, _07893_);
  nor (_07907_, _07906_, _07536_);
  nor (_07908_, _07907_, _07892_);
  nor (_07909_, _07908_, _07891_);
  nor (_07910_, _07909_, _07890_);
  nor (_07911_, _07910_, _07525_);
  and (_07912_, _07910_, _07525_);
  nor (_07913_, _07912_, _07911_);
  and (_07914_, _07913_, _07888_);
  or (_07915_, _07914_, _07889_);
  and (_07916_, _07915_, _07885_);
  and (_07917_, _02854_, _02530_);
  not (_07918_, _07888_);
  and (_07919_, _07913_, _07918_);
  or (_07920_, _07919_, _07917_);
  or (_07921_, _07920_, _07916_);
  not (_07922_, _07917_);
  and (_07923_, _07357_, \oc8051_golden_model_1.ACC [6]);
  nor (_07924_, _07358_, _07359_);
  and (_07925_, _07361_, \oc8051_golden_model_1.ACC [5]);
  and (_07926_, _07367_, \oc8051_golden_model_1.ACC [4]);
  and (_07927_, _07379_, \oc8051_golden_model_1.ACC [3]);
  and (_07928_, _07384_, \oc8051_golden_model_1.ACC [2]);
  and (_07929_, _07391_, \oc8051_golden_model_1.ACC [1]);
  and (_07930_, _07395_, \oc8051_golden_model_1.ACC [0]);
  not (_07931_, _07930_);
  nor (_07932_, _07931_, _07405_);
  nor (_07933_, _07932_, _07929_);
  nor (_07934_, _07933_, _07387_);
  nor (_07935_, _07934_, _07928_);
  nor (_07936_, _07935_, _07382_);
  nor (_07937_, _07936_, _07927_);
  nor (_07938_, _07937_, _07373_);
  nor (_07939_, _07938_, _07926_);
  nor (_07940_, _07939_, _07371_);
  nor (_07941_, _07940_, _07925_);
  nor (_07942_, _07941_, _07924_);
  nor (_07943_, _07942_, _07923_);
  nor (_07944_, _07943_, _07351_);
  and (_07945_, _07943_, _07351_);
  nor (_07946_, _07945_, _07944_);
  or (_07947_, _07946_, _07922_);
  and (_07948_, _07947_, _03138_);
  and (_07949_, _07948_, _07921_);
  and (_07950_, _03024_, _02530_);
  not (_07951_, _07610_);
  not (_07952_, _07651_);
  not (_07953_, _07670_);
  not (_07954_, _07681_);
  nor (_07955_, _07700_, _07319_);
  and (_07956_, _07955_, _07954_);
  and (_07957_, _07956_, _07953_);
  and (_07958_, _07957_, _07952_);
  nor (_07959_, _07640_, _07624_);
  and (_07960_, _07959_, _07958_);
  and (_07961_, _07960_, _07951_);
  nor (_07962_, _07961_, _05528_);
  and (_07963_, _07961_, _05528_);
  nor (_07964_, _07963_, _07962_);
  and (_07965_, _07964_, \oc8051_golden_model_1.ACC [7]);
  nor (_07966_, _07964_, \oc8051_golden_model_1.ACC [7]);
  nor (_07967_, _07966_, _07965_);
  nor (_07968_, _07960_, _07951_);
  nor (_07969_, _07968_, _07961_);
  and (_07970_, _07969_, \oc8051_golden_model_1.ACC [6]);
  and (_07971_, _07969_, _06833_);
  nor (_07972_, _07969_, _06833_);
  nor (_07973_, _07972_, _07971_);
  not (_07974_, _07624_);
  not (_07975_, _07640_);
  and (_07976_, _07958_, _07975_);
  nor (_07977_, _07976_, _07974_);
  nor (_07978_, _07977_, _07960_);
  and (_07979_, _07978_, \oc8051_golden_model_1.ACC [5]);
  and (_07980_, _07978_, _06879_);
  nor (_07981_, _07978_, _06879_);
  nor (_07982_, _07981_, _07980_);
  nor (_07983_, _07958_, _07975_);
  nor (_07984_, _07983_, _07976_);
  and (_07985_, _07984_, \oc8051_golden_model_1.ACC [4]);
  nor (_07986_, _07984_, _06885_);
  and (_07987_, _07984_, _06885_);
  nor (_07988_, _07987_, _07986_);
  nor (_07989_, _07957_, _07952_);
  nor (_07990_, _07989_, _07958_);
  and (_07991_, _07990_, \oc8051_golden_model_1.ACC [3]);
  nor (_07992_, _07990_, _02701_);
  and (_07993_, _07990_, _02701_);
  nor (_07994_, _07993_, _07992_);
  nor (_07995_, _07956_, _07953_);
  nor (_07996_, _07995_, _07957_);
  and (_07997_, _07996_, \oc8051_golden_model_1.ACC [2]);
  nor (_07998_, _07996_, _06984_);
  and (_07999_, _07996_, _06984_);
  nor (_08000_, _07999_, _07998_);
  nor (_08001_, _07955_, _07954_);
  nor (_08002_, _08001_, _07956_);
  and (_08003_, _08002_, \oc8051_golden_model_1.ACC [1]);
  and (_08004_, _08002_, _02618_);
  nor (_08005_, _08002_, _02618_);
  nor (_08006_, _08005_, _08004_);
  and (_08007_, _07700_, _07319_);
  nor (_08008_, _08007_, _07955_);
  and (_08009_, _08008_, \oc8051_golden_model_1.ACC [0]);
  not (_08010_, _08009_);
  nor (_08011_, _08010_, _08006_);
  nor (_08012_, _08011_, _08003_);
  nor (_08013_, _08012_, _08000_);
  nor (_08014_, _08013_, _07997_);
  nor (_08015_, _08014_, _07994_);
  nor (_08016_, _08015_, _07991_);
  nor (_08017_, _08016_, _07988_);
  nor (_08018_, _08017_, _07985_);
  nor (_08019_, _08018_, _07982_);
  nor (_08020_, _08019_, _07979_);
  nor (_08021_, _08020_, _07973_);
  nor (_08022_, _08021_, _07970_);
  nor (_08023_, _08022_, _07967_);
  and (_08024_, _08022_, _07967_);
  nor (_08025_, _08024_, _08023_);
  and (_08026_, _08025_, _03137_);
  or (_08027_, _08026_, _07950_);
  or (_08028_, _08027_, _07949_);
  and (_08029_, _02547_, _02530_);
  not (_08030_, _08029_);
  not (_08031_, _07950_);
  and (_08032_, _07290_, \oc8051_golden_model_1.ACC [6]);
  and (_08033_, _07296_, \oc8051_golden_model_1.ACC [5]);
  and (_08034_, _07301_, \oc8051_golden_model_1.ACC [4]);
  and (_08035_, _07307_, \oc8051_golden_model_1.ACC [3]);
  and (_08036_, _07311_, \oc8051_golden_model_1.ACC [2]);
  and (_08037_, _07322_, \oc8051_golden_model_1.ACC [1]);
  nor (_08038_, _07323_, _07324_);
  nor (_08039_, _07327_, _02549_);
  not (_08040_, _08039_);
  nor (_08041_, _08040_, _08038_);
  nor (_08042_, _08041_, _08037_);
  nor (_08043_, _08042_, _07317_);
  nor (_08044_, _08043_, _08036_);
  nor (_08045_, _08044_, _07315_);
  nor (_08046_, _08045_, _08035_);
  nor (_08047_, _08046_, _07304_);
  nor (_08048_, _08047_, _08034_);
  nor (_08049_, _08048_, _07299_);
  nor (_08050_, _08049_, _08033_);
  nor (_08051_, _08050_, _07293_);
  nor (_08052_, _08051_, _08032_);
  nor (_08053_, _08052_, _07287_);
  and (_08054_, _08052_, _07287_);
  nor (_08055_, _08054_, _08053_);
  or (_08056_, _08055_, _08031_);
  and (_08057_, _08056_, _08030_);
  and (_08058_, _08057_, _08028_);
  and (_08059_, _08029_, \oc8051_golden_model_1.ACC [6]);
  or (_08060_, _08059_, _07258_);
  or (_08061_, _08060_, _08058_);
  and (_08062_, _08061_, _07260_);
  or (_08063_, _08062_, _07217_);
  not (_08064_, _07217_);
  and (_08065_, _05847_, \oc8051_golden_model_1.ACC [6]);
  nor (_08066_, _05847_, \oc8051_golden_model_1.ACC [6]);
  nor (_08067_, _08065_, _08066_);
  and (_08068_, _06180_, \oc8051_golden_model_1.ACC [5]);
  and (_08069_, _06076_, _06879_);
  and (_08070_, _06181_, \oc8051_golden_model_1.ACC [4]);
  and (_08071_, _06121_, _06885_);
  nor (_08072_, _08070_, _08071_);
  and (_08073_, _05984_, _02701_);
  not (_08074_, _08073_);
  and (_08075_, _06176_, \oc8051_golden_model_1.ACC [3]);
  not (_08076_, _08075_);
  and (_08077_, _06177_, \oc8051_golden_model_1.ACC [2]);
  and (_08078_, _06029_, _06984_);
  nor (_08079_, _08077_, _08078_);
  not (_08080_, _08079_);
  and (_08081_, _06173_, \oc8051_golden_model_1.ACC [1]);
  and (_08082_, _05893_, _02618_);
  nor (_08083_, _08081_, _08082_);
  and (_08084_, _06174_, \oc8051_golden_model_1.ACC [0]);
  and (_08085_, _08084_, _08083_);
  nor (_08086_, _08085_, _08081_);
  nor (_08087_, _08086_, _08080_);
  nor (_08088_, _08087_, _08077_);
  nand (_08089_, _08088_, _08076_);
  and (_08090_, _08089_, _08074_);
  and (_08091_, _08090_, _08072_);
  nor (_08092_, _08091_, _08070_);
  nor (_08093_, _08092_, _08069_);
  or (_08094_, _08093_, _08068_);
  and (_08095_, _08094_, _08067_);
  nor (_08096_, _08095_, _08065_);
  nor (_08097_, _08096_, _07808_);
  and (_08098_, _08096_, _07808_);
  or (_08099_, _08098_, _08097_);
  or (_08100_, _08099_, _08064_);
  and (_08101_, _08100_, _02901_);
  and (_08102_, _08101_, _08063_);
  and (_08103_, _03024_, _02535_);
  nor (_08104_, _08103_, _02899_);
  not (_08105_, _08104_);
  not (_08106_, _08103_);
  nor (_08107_, _07610_, _06833_);
  nor (_08108_, _07624_, _06879_);
  nor (_08109_, _07640_, _06885_);
  not (_08110_, _07711_);
  nor (_08111_, _07670_, _06984_);
  nor (_08112_, _07681_, _02618_);
  nor (_08113_, _07700_, _02549_);
  not (_08114_, _08113_);
  nor (_08115_, _08114_, _07732_);
  nor (_08116_, _08115_, _08112_);
  nor (_08117_, _08116_, _07705_);
  nor (_08118_, _08117_, _08111_);
  nor (_08119_, _08118_, _07651_);
  or (_08120_, _08119_, \oc8051_golden_model_1.ACC [3]);
  nand (_08121_, _08118_, _07651_);
  and (_08122_, _08121_, _08120_);
  and (_08123_, _08122_, _08110_);
  nor (_08124_, _08123_, _08109_);
  nor (_08125_, _08124_, _07724_);
  nor (_08126_, _08125_, _08108_);
  nor (_08127_, _08126_, _07613_);
  nor (_08128_, _08127_, _08107_);
  nor (_08129_, _08128_, _07600_);
  and (_08130_, _08128_, _07600_);
  nor (_08131_, _08130_, _08129_);
  nand (_08132_, _08131_, _08106_);
  and (_08133_, _08132_, _08105_);
  or (_08134_, _08133_, _08102_);
  and (_08135_, _02547_, _02535_);
  not (_08136_, _08135_);
  nor (_08137_, _02932_, _06833_);
  and (_08138_, _02932_, _06833_);
  nor (_08139_, _08138_, _08137_);
  nor (_08140_, _03215_, _06879_);
  and (_08141_, _03215_, _06879_);
  nor (_08142_, _08141_, _08140_);
  not (_08143_, _08142_);
  nor (_08144_, _03625_, _06885_);
  and (_08145_, _03625_, _06885_);
  or (_08146_, _08145_, _08144_);
  not (_08147_, _08146_);
  nor (_08148_, _02799_, _02701_);
  and (_08149_, _02799_, _02701_);
  nor (_08150_, _03260_, _06984_);
  and (_08151_, _03260_, _06984_);
  nor (_08152_, _08151_, _08150_);
  not (_08153_, _08152_);
  nor (_08154_, _03671_, _02618_);
  and (_08155_, _03671_, _02618_);
  nor (_08156_, _08155_, _08154_);
  nor (_08157_, _02832_, _02549_);
  and (_08158_, _08157_, _08156_);
  nor (_08159_, _08158_, _08154_);
  nor (_08160_, _08159_, _08153_);
  nor (_08161_, _08160_, _08150_);
  nor (_08162_, _08161_, _08149_);
  or (_08163_, _08162_, _08148_);
  and (_08164_, _08163_, _08147_);
  nor (_08165_, _08164_, _08144_);
  nor (_08166_, _08165_, _08143_);
  or (_08167_, _08166_, _08140_);
  and (_08168_, _08167_, _08139_);
  nor (_08169_, _08168_, _08137_);
  nor (_08170_, _08169_, _07820_);
  and (_08171_, _08169_, _07820_);
  or (_08172_, _08171_, _08170_);
  or (_08173_, _08172_, _08106_);
  and (_08174_, _08173_, _08136_);
  and (_08175_, _08174_, _08134_);
  and (_08176_, _08135_, \oc8051_golden_model_1.ACC [6]);
  or (_08177_, _08176_, _03166_);
  or (_08178_, _08177_, _08175_);
  and (_08179_, _03024_, _02370_);
  not (_08180_, _08179_);
  nand (_08181_, _07457_, _03166_);
  and (_08182_, _08181_, _08180_);
  and (_08183_, _08182_, _08178_);
  and (_08184_, _02547_, _02370_);
  nor (_08185_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08186_, _08185_, _06925_);
  and (_08187_, _08186_, _06849_);
  and (_08188_, _08187_, _06833_);
  nor (_08189_, _08188_, _05768_);
  and (_08190_, _08188_, _05768_);
  nor (_08191_, _08190_, _08189_);
  nor (_08192_, _08191_, _08180_);
  or (_08193_, _08192_, _08184_);
  or (_08194_, _08193_, _08183_);
  nand (_08195_, _08184_, _07319_);
  and (_08196_, _08195_, _02501_);
  and (_08197_, _08196_, _08194_);
  nor (_08198_, _07505_, _02501_);
  or (_08199_, _08198_, _03174_);
  or (_08200_, _08199_, _08197_);
  and (_08201_, _03024_, _02525_);
  not (_08202_, _08201_);
  and (_08203_, _05257_, _04712_);
  nor (_08204_, _08203_, _07268_);
  nand (_08205_, _08204_, _03174_);
  and (_08206_, _08205_, _08202_);
  and (_08207_, _08206_, _08200_);
  and (_08208_, _02547_, _02525_);
  and (_08209_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08210_, _08209_, _06926_);
  nor (_08211_, _08210_, _06885_);
  and (_08212_, _08211_, \oc8051_golden_model_1.ACC [5]);
  and (_08213_, _08212_, \oc8051_golden_model_1.ACC [6]);
  nor (_08214_, _08213_, \oc8051_golden_model_1.ACC [7]);
  and (_08215_, _08213_, \oc8051_golden_model_1.ACC [7]);
  nor (_08216_, _08215_, _08214_);
  and (_08217_, _08216_, _08201_);
  or (_08218_, _08217_, _08208_);
  or (_08219_, _08218_, _08207_);
  nand (_08220_, _08208_, _02549_);
  and (_08221_, _08220_, _34698_);
  and (_08222_, _08221_, _08219_);
  or (_08223_, _08222_, _07216_);
  and (_32486_, _08223_, _36029_);
  or (_08224_, _34698_, \oc8051_golden_model_1.DPL [7]);
  and (_08225_, _08224_, _36029_);
  not (_08226_, \oc8051_golden_model_1.DPL [7]);
  nor (_08227_, _04654_, _08226_);
  and (_08228_, _05771_, _04654_);
  or (_08229_, _08228_, _08227_);
  and (_08230_, _08229_, _03130_);
  not (_08231_, _04654_);
  nor (_08232_, _08231_, _04623_);
  or (_08233_, _08232_, _08227_);
  or (_08234_, _08233_, _06241_);
  not (_08235_, _03023_);
  and (_08236_, _05502_, _04654_);
  or (_08237_, _08236_, _08227_);
  or (_08238_, _08237_, _03821_);
  and (_08239_, _04654_, \oc8051_golden_model_1.ACC [7]);
  or (_08240_, _08239_, _08227_);
  and (_08241_, _08240_, _03825_);
  nor (_08242_, _03825_, _08226_);
  or (_08243_, _08242_, _02952_);
  or (_08244_, _08243_, _08241_);
  and (_08245_, _08244_, _03327_);
  and (_08246_, _08245_, _08238_);
  and (_08247_, _08233_, _02947_);
  or (_08248_, _08247_, _02950_);
  or (_08249_, _08248_, _08246_);
  and (_08250_, _02980_, _02547_);
  not (_08251_, _08250_);
  or (_08252_, _08240_, _02959_);
  and (_08253_, _08252_, _08251_);
  and (_08254_, _08253_, _08249_);
  and (_08255_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08256_, _08255_, \oc8051_golden_model_1.DPL [2]);
  and (_08257_, _08256_, \oc8051_golden_model_1.DPL [3]);
  and (_08258_, _08257_, \oc8051_golden_model_1.DPL [4]);
  and (_08259_, _08258_, \oc8051_golden_model_1.DPL [5]);
  and (_08260_, _08259_, \oc8051_golden_model_1.DPL [6]);
  nor (_08261_, _08260_, \oc8051_golden_model_1.DPL [7]);
  and (_08262_, _08260_, \oc8051_golden_model_1.DPL [7]);
  nor (_08263_, _08262_, _08261_);
  and (_08264_, _08263_, _08250_);
  or (_08265_, _08264_, _08254_);
  and (_08266_, _08265_, _08235_);
  nor (_08267_, _05311_, _08235_);
  or (_08268_, _08267_, _06793_);
  or (_08269_, _08268_, _08266_);
  and (_08270_, _08269_, _08234_);
  or (_08271_, _08270_, _02855_);
  and (_08272_, _05490_, _04654_);
  or (_08273_, _08227_, _02856_);
  or (_08274_, _08273_, _08272_);
  and (_08275_, _08274_, _02851_);
  and (_08276_, _08275_, _08271_);
  nor (_08277_, _05755_, _08231_);
  or (_08278_, _08277_, _08227_);
  and (_08279_, _08278_, _02576_);
  or (_08280_, _08279_, _03014_);
  or (_08281_, _08280_, _08276_);
  and (_08282_, _05563_, _04654_);
  or (_08283_, _08282_, _08227_);
  or (_08284_, _08283_, _03884_);
  and (_08285_, _08284_, _08281_);
  or (_08286_, _08285_, _03021_);
  and (_08287_, _05314_, _04654_);
  or (_08288_, _08227_, _05279_);
  or (_08289_, _08288_, _08287_);
  and (_08290_, _08289_, _03131_);
  and (_08291_, _08290_, _08286_);
  or (_08292_, _08291_, _08230_);
  and (_08293_, _08292_, _05274_);
  or (_08294_, _08227_, _04733_);
  and (_08295_, _08283_, _03020_);
  and (_08296_, _08295_, _08294_);
  or (_08297_, _08296_, _08293_);
  and (_08298_, _08297_, _03140_);
  and (_08299_, _08240_, _03139_);
  and (_08300_, _08299_, _08294_);
  or (_08301_, _08300_, _03036_);
  or (_08302_, _08301_, _08298_);
  nor (_08303_, _05312_, _08231_);
  or (_08304_, _08227_, _05781_);
  or (_08305_, _08304_, _08303_);
  and (_08306_, _08305_, _05786_);
  and (_08307_, _08306_, _08302_);
  nor (_08308_, _05770_, _08231_);
  or (_08309_, _08308_, _08227_);
  and (_08310_, _08309_, _03127_);
  or (_08311_, _08310_, _03166_);
  or (_08312_, _08311_, _08307_);
  or (_08313_, _08237_, _03563_);
  and (_08314_, _08313_, _03178_);
  and (_08315_, _08314_, _08312_);
  and (_08316_, _05257_, _04654_);
  or (_08317_, _08316_, _08227_);
  and (_08318_, _08317_, _03174_);
  or (_08319_, _08318_, _34702_);
  or (_08320_, _08319_, _08315_);
  and (_32487_, _08320_, _08225_);
  or (_08321_, _34698_, \oc8051_golden_model_1.DPH [7]);
  and (_08322_, _08321_, _36029_);
  not (_08323_, \oc8051_golden_model_1.DPH [7]);
  nor (_08324_, _05038_, _08323_);
  and (_08325_, _05771_, _04632_);
  or (_08326_, _08325_, _08324_);
  and (_08327_, _08326_, _03130_);
  not (_08328_, _04632_);
  nor (_08329_, _08328_, _04623_);
  or (_08330_, _08329_, _08324_);
  or (_08331_, _08330_, _06241_);
  and (_08332_, _05502_, _04632_);
  or (_08333_, _08332_, _08324_);
  or (_08334_, _08333_, _03821_);
  and (_08335_, _05038_, \oc8051_golden_model_1.ACC [7]);
  or (_08336_, _08335_, _08324_);
  and (_08337_, _08336_, _03825_);
  nor (_08338_, _03825_, _08323_);
  or (_08339_, _08338_, _02952_);
  or (_08340_, _08339_, _08337_);
  and (_08341_, _08340_, _03327_);
  and (_08342_, _08341_, _08334_);
  and (_08343_, _08330_, _02947_);
  or (_08344_, _08343_, _02950_);
  or (_08345_, _08344_, _08342_);
  or (_08346_, _08336_, _02959_);
  and (_08347_, _08346_, _08251_);
  and (_08348_, _08347_, _08345_);
  and (_08349_, _08262_, \oc8051_golden_model_1.DPH [0]);
  and (_08350_, _08349_, \oc8051_golden_model_1.DPH [1]);
  and (_08351_, _08350_, \oc8051_golden_model_1.DPH [2]);
  and (_08352_, _08351_, \oc8051_golden_model_1.DPH [3]);
  and (_08353_, _08352_, \oc8051_golden_model_1.DPH [4]);
  and (_08354_, _08353_, \oc8051_golden_model_1.DPH [5]);
  and (_08355_, _08354_, \oc8051_golden_model_1.DPH [6]);
  nand (_08356_, _08355_, \oc8051_golden_model_1.DPH [7]);
  or (_08357_, _08355_, \oc8051_golden_model_1.DPH [7]);
  and (_08358_, _08357_, _08250_);
  and (_08359_, _08358_, _08356_);
  or (_08360_, _08359_, _08348_);
  and (_08361_, _08360_, _08235_);
  and (_08362_, _03023_, _02768_);
  or (_08363_, _08362_, _06793_);
  or (_08364_, _08363_, _08361_);
  and (_08365_, _08364_, _08331_);
  or (_08366_, _08365_, _02855_);
  or (_08367_, _08324_, _02856_);
  and (_08368_, _05490_, _05038_);
  or (_08369_, _08368_, _08367_);
  and (_08370_, _08369_, _02851_);
  and (_08371_, _08370_, _08366_);
  not (_08372_, _05038_);
  nor (_08373_, _05755_, _08372_);
  or (_08374_, _08373_, _08324_);
  and (_08375_, _08374_, _02576_);
  or (_08376_, _08375_, _03014_);
  or (_08377_, _08376_, _08371_);
  and (_08378_, _05563_, _05038_);
  or (_08379_, _08378_, _08324_);
  or (_08380_, _08379_, _03884_);
  and (_08381_, _08380_, _08377_);
  or (_08382_, _08381_, _03021_);
  and (_08383_, _05314_, _04632_);
  or (_08384_, _08324_, _05279_);
  or (_08385_, _08384_, _08383_);
  and (_08386_, _08385_, _03131_);
  and (_08387_, _08386_, _08382_);
  or (_08388_, _08387_, _08327_);
  and (_08389_, _08388_, _05274_);
  or (_08390_, _08324_, _04733_);
  and (_08391_, _08379_, _03020_);
  and (_08392_, _08391_, _08390_);
  or (_08393_, _08392_, _08389_);
  and (_08394_, _08393_, _03140_);
  and (_08395_, _08336_, _03139_);
  and (_08396_, _08395_, _08390_);
  or (_08397_, _08396_, _03036_);
  or (_08398_, _08397_, _08394_);
  nor (_08399_, _05312_, _08328_);
  or (_08400_, _08324_, _05781_);
  or (_08401_, _08400_, _08399_);
  and (_08402_, _08401_, _05786_);
  and (_08403_, _08402_, _08398_);
  nor (_08404_, _05770_, _08328_);
  or (_08405_, _08404_, _08324_);
  and (_08406_, _08405_, _03127_);
  or (_08407_, _08406_, _03166_);
  or (_08408_, _08407_, _08403_);
  or (_08409_, _08333_, _03563_);
  and (_08410_, _08409_, _03178_);
  and (_08411_, _08410_, _08408_);
  and (_08412_, _05257_, _04632_);
  or (_08413_, _08412_, _08324_);
  and (_08414_, _08413_, _03174_);
  or (_08415_, _08414_, _34702_);
  or (_08416_, _08415_, _08411_);
  and (_32488_, _08416_, _08322_);
  and (_32489_, \oc8051_golden_model_1.IE [7], _36029_);
  and (_32490_, \oc8051_golden_model_1.IP [7], _36029_);
  not (_08417_, \oc8051_golden_model_1.P0 [7]);
  nor (_08418_, _34698_, _08417_);
  or (_08419_, _08418_, rst);
  nor (_08420_, _04716_, _08417_);
  and (_08421_, _05771_, _04716_);
  or (_08422_, _08421_, _08420_);
  and (_08423_, _08422_, _03130_);
  not (_08424_, _04716_);
  nor (_08425_, _08424_, _04623_);
  or (_08426_, _08425_, _08420_);
  or (_08427_, _08426_, _06241_);
  nor (_08428_, _04629_, _08417_);
  and (_08429_, _05380_, _04629_);
  or (_08430_, _08429_, _08428_);
  and (_08431_, _08430_, _02887_);
  and (_08432_, _05502_, _04716_);
  or (_08433_, _08432_, _08420_);
  or (_08434_, _08433_, _03821_);
  and (_08435_, _04716_, \oc8051_golden_model_1.ACC [7]);
  or (_08436_, _08435_, _08420_);
  and (_08437_, _08436_, _03825_);
  nor (_08438_, _03825_, _08417_);
  or (_08439_, _08438_, _02952_);
  or (_08440_, _08439_, _08437_);
  and (_08441_, _08440_, _02892_);
  and (_08442_, _08441_, _08434_);
  and (_08443_, _05385_, _04629_);
  or (_08444_, _08443_, _08428_);
  and (_08445_, _08444_, _02891_);
  or (_08446_, _08445_, _02947_);
  or (_08447_, _08446_, _08442_);
  or (_08448_, _08426_, _03327_);
  and (_08449_, _08448_, _08447_);
  or (_08450_, _08449_, _02950_);
  or (_08451_, _08436_, _02959_);
  and (_08452_, _08451_, _02888_);
  and (_08453_, _08452_, _08450_);
  or (_08454_, _08453_, _08431_);
  and (_08455_, _08454_, _02881_);
  or (_08456_, _08428_, _05533_);
  and (_08457_, _08456_, _02880_);
  and (_08458_, _08457_, _08444_);
  or (_08459_, _08458_, _08455_);
  and (_08460_, _08459_, _02875_);
  or (_08461_, _05380_, _05365_);
  and (_08462_, _08461_, _04629_);
  or (_08463_, _08462_, _08428_);
  and (_08464_, _08463_, _02874_);
  or (_08465_, _08464_, _06793_);
  or (_08466_, _08465_, _08460_);
  and (_08467_, _08466_, _08427_);
  or (_08468_, _08467_, _02855_);
  and (_08469_, _05490_, _04716_);
  or (_08470_, _08420_, _02856_);
  or (_08471_, _08470_, _08469_);
  and (_08472_, _08471_, _02851_);
  and (_08473_, _08472_, _08468_);
  and (_08474_, _05736_, \oc8051_golden_model_1.P0 [7]);
  and (_08475_, _05733_, \oc8051_golden_model_1.P1 [7]);
  and (_08476_, _05739_, \oc8051_golden_model_1.P2 [7]);
  and (_08477_, _05741_, \oc8051_golden_model_1.P3 [7]);
  or (_08478_, _08477_, _08476_);
  or (_08479_, _08478_, _08475_);
  nor (_08480_, _08479_, _08474_);
  and (_08481_, _08480_, _05751_);
  and (_08482_, _08481_, _05732_);
  nand (_08483_, _08482_, _05719_);
  or (_08484_, _08483_, _05564_);
  and (_08485_, _08484_, _04716_);
  or (_08486_, _08485_, _08420_);
  and (_08487_, _08486_, _02576_);
  or (_08488_, _08487_, _03014_);
  or (_08489_, _08488_, _08473_);
  and (_08490_, _05563_, _04716_);
  or (_08491_, _08490_, _08420_);
  or (_08492_, _08491_, _03884_);
  and (_08493_, _08492_, _08489_);
  or (_08494_, _08493_, _03021_);
  and (_08495_, _05314_, _04716_);
  or (_08496_, _08420_, _05279_);
  or (_08497_, _08496_, _08495_);
  and (_08498_, _08497_, _03131_);
  and (_08499_, _08498_, _08494_);
  or (_08500_, _08499_, _08423_);
  and (_08501_, _08500_, _05274_);
  or (_08502_, _08420_, _04733_);
  and (_08503_, _08491_, _03020_);
  and (_08504_, _08503_, _08502_);
  or (_08505_, _08504_, _08501_);
  and (_08506_, _08505_, _03140_);
  and (_08507_, _08436_, _03139_);
  and (_08508_, _08507_, _08502_);
  or (_08509_, _08508_, _03036_);
  or (_08510_, _08509_, _08506_);
  nor (_08511_, _05312_, _08424_);
  or (_08512_, _08420_, _05781_);
  or (_08513_, _08512_, _08511_);
  and (_08514_, _08513_, _05786_);
  and (_08515_, _08514_, _08510_);
  nor (_08516_, _05770_, _08424_);
  or (_08517_, _08516_, _08420_);
  and (_08518_, _08517_, _03127_);
  or (_08519_, _08518_, _03166_);
  or (_08520_, _08519_, _08515_);
  or (_08521_, _08433_, _03563_);
  and (_08522_, _08521_, _02501_);
  and (_08523_, _08522_, _08520_);
  and (_08524_, _08430_, _02500_);
  or (_08525_, _08524_, _03174_);
  or (_08526_, _08525_, _08523_);
  and (_08527_, _05257_, _04716_);
  or (_08528_, _08420_, _03178_);
  or (_08529_, _08528_, _08527_);
  and (_08530_, _08529_, _34698_);
  and (_08531_, _08530_, _08526_);
  or (_32491_, _08531_, _08419_);
  not (_08532_, \oc8051_golden_model_1.P1 [7]);
  nor (_08533_, _34698_, _08532_);
  or (_08534_, _08533_, rst);
  nor (_08535_, _04719_, _08532_);
  and (_08536_, _05771_, _04719_);
  or (_08537_, _08536_, _08535_);
  and (_08538_, _08537_, _03130_);
  not (_08539_, _04719_);
  nor (_08540_, _08539_, _04623_);
  or (_08541_, _08540_, _08535_);
  or (_08542_, _08541_, _06241_);
  nor (_08543_, _05344_, _08532_);
  and (_08544_, _05380_, _05344_);
  or (_08545_, _08544_, _08543_);
  and (_08546_, _08545_, _02887_);
  and (_08547_, _05502_, _04719_);
  or (_08548_, _08547_, _08535_);
  or (_08549_, _08548_, _03821_);
  and (_08550_, _04719_, \oc8051_golden_model_1.ACC [7]);
  or (_08551_, _08550_, _08535_);
  and (_08552_, _08551_, _03825_);
  nor (_08553_, _03825_, _08532_);
  or (_08554_, _08553_, _02952_);
  or (_08555_, _08554_, _08552_);
  and (_08556_, _08555_, _02892_);
  and (_08557_, _08556_, _08549_);
  and (_08558_, _05385_, _05344_);
  or (_08559_, _08558_, _08543_);
  and (_08560_, _08559_, _02891_);
  or (_08561_, _08560_, _02947_);
  or (_08562_, _08561_, _08557_);
  or (_08563_, _08541_, _03327_);
  and (_08564_, _08563_, _08562_);
  or (_08565_, _08564_, _02950_);
  or (_08566_, _08551_, _02959_);
  and (_08567_, _08566_, _02888_);
  and (_08568_, _08567_, _08565_);
  or (_08569_, _08568_, _08546_);
  and (_08570_, _08569_, _02881_);
  and (_08571_, _05534_, _05344_);
  or (_08572_, _08571_, _08543_);
  and (_08573_, _08572_, _02880_);
  or (_08574_, _08573_, _08570_);
  and (_08575_, _08574_, _02875_);
  and (_08576_, _08461_, _05344_);
  or (_08577_, _08576_, _08543_);
  and (_08578_, _08577_, _02874_);
  or (_08579_, _08578_, _06793_);
  or (_08580_, _08579_, _08575_);
  and (_08581_, _08580_, _08542_);
  or (_08582_, _08581_, _02855_);
  and (_08583_, _05490_, _04719_);
  or (_08584_, _08535_, _02856_);
  or (_08585_, _08584_, _08583_);
  and (_08586_, _08585_, _02851_);
  and (_08587_, _08586_, _08582_);
  and (_08588_, _08484_, _04719_);
  or (_08589_, _08588_, _08535_);
  and (_08590_, _08589_, _02576_);
  or (_08591_, _08590_, _03014_);
  or (_08592_, _08591_, _08587_);
  and (_08593_, _05563_, _04719_);
  or (_08594_, _08593_, _08535_);
  or (_08595_, _08594_, _03884_);
  and (_08596_, _08595_, _08592_);
  or (_08597_, _08596_, _03021_);
  and (_08598_, _05314_, _04719_);
  or (_08599_, _08535_, _05279_);
  or (_08600_, _08599_, _08598_);
  and (_08601_, _08600_, _03131_);
  and (_08602_, _08601_, _08597_);
  or (_08603_, _08602_, _08538_);
  and (_08604_, _08603_, _05274_);
  or (_08605_, _08535_, _04733_);
  and (_08606_, _08594_, _03020_);
  and (_08607_, _08606_, _08605_);
  or (_08608_, _08607_, _08604_);
  and (_08609_, _08608_, _03140_);
  and (_08610_, _08551_, _03139_);
  and (_08611_, _08610_, _08605_);
  or (_08612_, _08611_, _03036_);
  or (_08613_, _08612_, _08609_);
  nor (_08614_, _05312_, _08539_);
  or (_08615_, _08535_, _05781_);
  or (_08616_, _08615_, _08614_);
  and (_08617_, _08616_, _05786_);
  and (_08618_, _08617_, _08613_);
  nor (_08619_, _05770_, _08539_);
  or (_08620_, _08619_, _08535_);
  and (_08621_, _08620_, _03127_);
  or (_08622_, _08621_, _03166_);
  or (_08623_, _08622_, _08618_);
  or (_08624_, _08548_, _03563_);
  and (_08625_, _08624_, _02501_);
  and (_08626_, _08625_, _08623_);
  and (_08627_, _08545_, _02500_);
  or (_08628_, _08627_, _03174_);
  or (_08629_, _08628_, _08626_);
  and (_08630_, _05257_, _04719_);
  or (_08631_, _08535_, _03178_);
  or (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _34698_);
  and (_08634_, _08633_, _08629_);
  or (_32492_, _08634_, _08534_);
  not (_08635_, \oc8051_golden_model_1.P2 [7]);
  nor (_08636_, _34698_, _08635_);
  or (_08637_, _08636_, rst);
  nor (_08638_, _04722_, _08635_);
  and (_08639_, _05771_, _04722_);
  or (_08640_, _08639_, _08638_);
  and (_08641_, _08640_, _03130_);
  not (_08642_, _04722_);
  nor (_08643_, _08642_, _04623_);
  or (_08644_, _08643_, _08638_);
  or (_08645_, _08644_, _06241_);
  nor (_08646_, _05346_, _08635_);
  and (_08647_, _05380_, _05346_);
  or (_08648_, _08647_, _08646_);
  and (_08649_, _08648_, _02887_);
  and (_08650_, _05502_, _04722_);
  or (_08651_, _08650_, _08638_);
  or (_08652_, _08651_, _03821_);
  and (_08653_, _04722_, \oc8051_golden_model_1.ACC [7]);
  or (_08654_, _08653_, _08638_);
  and (_08655_, _08654_, _03825_);
  nor (_08656_, _03825_, _08635_);
  or (_08657_, _08656_, _02952_);
  or (_08658_, _08657_, _08655_);
  and (_08659_, _08658_, _02892_);
  and (_08660_, _08659_, _08652_);
  and (_08661_, _05385_, _05346_);
  or (_08662_, _08661_, _08646_);
  and (_08663_, _08662_, _02891_);
  or (_08664_, _08663_, _02947_);
  or (_08665_, _08664_, _08660_);
  or (_08666_, _08644_, _03327_);
  and (_08667_, _08666_, _08665_);
  or (_08668_, _08667_, _02950_);
  or (_08669_, _08654_, _02959_);
  and (_08670_, _08669_, _02888_);
  and (_08671_, _08670_, _08668_);
  or (_08672_, _08671_, _08649_);
  and (_08673_, _08672_, _02881_);
  or (_08674_, _08646_, _05533_);
  and (_08675_, _08674_, _02880_);
  and (_08676_, _08675_, _08662_);
  or (_08677_, _08676_, _08673_);
  and (_08678_, _08677_, _02875_);
  and (_08679_, _08461_, _05346_);
  or (_08680_, _08679_, _08646_);
  and (_08681_, _08680_, _02874_);
  or (_08682_, _08681_, _06793_);
  or (_08683_, _08682_, _08678_);
  and (_08684_, _08683_, _08645_);
  or (_08685_, _08684_, _02855_);
  and (_08686_, _05490_, _04722_);
  or (_08687_, _08638_, _02856_);
  or (_08688_, _08687_, _08686_);
  and (_08689_, _08688_, _02851_);
  and (_08690_, _08689_, _08685_);
  and (_08691_, _08484_, _04722_);
  or (_08692_, _08691_, _08638_);
  and (_08693_, _08692_, _02576_);
  or (_08694_, _08693_, _03014_);
  or (_08695_, _08694_, _08690_);
  and (_08696_, _05563_, _04722_);
  or (_08697_, _08696_, _08638_);
  or (_08698_, _08697_, _03884_);
  and (_08699_, _08698_, _08695_);
  or (_08700_, _08699_, _03021_);
  and (_08701_, _05314_, _04722_);
  or (_08702_, _08638_, _05279_);
  or (_08703_, _08702_, _08701_);
  and (_08704_, _08703_, _03131_);
  and (_08705_, _08704_, _08700_);
  or (_08706_, _08705_, _08641_);
  and (_08707_, _08706_, _05274_);
  or (_08708_, _08638_, _04733_);
  and (_08709_, _08697_, _03020_);
  and (_08710_, _08709_, _08708_);
  or (_08711_, _08710_, _08707_);
  and (_08712_, _08711_, _03140_);
  and (_08713_, _08654_, _03139_);
  and (_08714_, _08713_, _08708_);
  or (_08715_, _08714_, _03036_);
  or (_08716_, _08715_, _08712_);
  nor (_08717_, _05312_, _08642_);
  or (_08718_, _08638_, _05781_);
  or (_08719_, _08718_, _08717_);
  and (_08720_, _08719_, _05786_);
  and (_08721_, _08720_, _08716_);
  nor (_08722_, _05770_, _08642_);
  or (_08723_, _08722_, _08638_);
  and (_08724_, _08723_, _03127_);
  or (_08725_, _08724_, _03166_);
  or (_08726_, _08725_, _08721_);
  or (_08727_, _08651_, _03563_);
  and (_08728_, _08727_, _02501_);
  and (_08729_, _08728_, _08726_);
  and (_08730_, _08648_, _02500_);
  or (_08731_, _08730_, _03174_);
  or (_08732_, _08731_, _08729_);
  and (_08733_, _05257_, _04722_);
  or (_08734_, _08638_, _03178_);
  or (_08735_, _08734_, _08733_);
  and (_08736_, _08735_, _34698_);
  and (_08737_, _08736_, _08732_);
  or (_32493_, _08737_, _08637_);
  not (_08738_, \oc8051_golden_model_1.P3 [7]);
  nor (_08739_, _34698_, _08738_);
  or (_08740_, _08739_, rst);
  nor (_08741_, _04724_, _08738_);
  and (_08742_, _05771_, _04724_);
  or (_08743_, _08742_, _08741_);
  and (_08744_, _08743_, _03130_);
  not (_08745_, _04724_);
  nor (_08746_, _08745_, _04623_);
  or (_08747_, _08746_, _08741_);
  or (_08748_, _08747_, _06241_);
  nor (_08749_, _05357_, _08738_);
  and (_08750_, _05380_, _05357_);
  or (_08751_, _08750_, _08749_);
  and (_08752_, _08751_, _02887_);
  and (_08753_, _05502_, _04724_);
  or (_08754_, _08753_, _08741_);
  or (_08755_, _08754_, _03821_);
  and (_08756_, _04724_, \oc8051_golden_model_1.ACC [7]);
  or (_08757_, _08756_, _08741_);
  and (_08758_, _08757_, _03825_);
  nor (_08759_, _03825_, _08738_);
  or (_08760_, _08759_, _02952_);
  or (_08761_, _08760_, _08758_);
  and (_08762_, _08761_, _02892_);
  and (_08763_, _08762_, _08755_);
  and (_08764_, _05385_, _05357_);
  or (_08765_, _08764_, _08749_);
  and (_08766_, _08765_, _02891_);
  or (_08767_, _08766_, _02947_);
  or (_08768_, _08767_, _08763_);
  or (_08769_, _08747_, _03327_);
  and (_08770_, _08769_, _08768_);
  or (_08771_, _08770_, _02950_);
  or (_08772_, _08757_, _02959_);
  and (_08773_, _08772_, _02888_);
  and (_08774_, _08773_, _08771_);
  or (_08775_, _08774_, _08752_);
  and (_08776_, _08775_, _02881_);
  and (_08777_, _05534_, _05357_);
  or (_08778_, _08777_, _08749_);
  and (_08779_, _08778_, _02880_);
  or (_08780_, _08779_, _08776_);
  and (_08781_, _08780_, _02875_);
  and (_08782_, _08461_, _05357_);
  or (_08783_, _08782_, _08749_);
  and (_08784_, _08783_, _02874_);
  or (_08785_, _08784_, _06793_);
  or (_08786_, _08785_, _08781_);
  and (_08787_, _08786_, _08748_);
  or (_08788_, _08787_, _02855_);
  and (_08789_, _05490_, _04724_);
  or (_08790_, _08741_, _02856_);
  or (_08791_, _08790_, _08789_);
  and (_08792_, _08791_, _02851_);
  and (_08793_, _08792_, _08788_);
  and (_08794_, _08484_, _04724_);
  or (_08795_, _08794_, _08741_);
  and (_08796_, _08795_, _02576_);
  or (_08797_, _08796_, _03014_);
  or (_08798_, _08797_, _08793_);
  and (_08799_, _05563_, _04724_);
  or (_08800_, _08799_, _08741_);
  or (_08801_, _08800_, _03884_);
  and (_08802_, _08801_, _08798_);
  or (_08803_, _08802_, _03021_);
  and (_08804_, _05314_, _04724_);
  or (_08805_, _08741_, _05279_);
  or (_08806_, _08805_, _08804_);
  and (_08807_, _08806_, _03131_);
  and (_08808_, _08807_, _08803_);
  or (_08809_, _08808_, _08744_);
  and (_08810_, _08809_, _05274_);
  or (_08811_, _08741_, _04733_);
  and (_08812_, _08800_, _03020_);
  and (_08813_, _08812_, _08811_);
  or (_08814_, _08813_, _08810_);
  and (_08815_, _08814_, _03140_);
  and (_08816_, _08757_, _03139_);
  and (_08817_, _08816_, _08811_);
  or (_08818_, _08817_, _03036_);
  or (_08819_, _08818_, _08815_);
  nor (_08820_, _05312_, _08745_);
  or (_08821_, _08741_, _05781_);
  or (_08822_, _08821_, _08820_);
  and (_08823_, _08822_, _05786_);
  and (_08824_, _08823_, _08819_);
  nor (_08825_, _05770_, _08745_);
  or (_08826_, _08825_, _08741_);
  and (_08827_, _08826_, _03127_);
  or (_08828_, _08827_, _03166_);
  or (_08829_, _08828_, _08824_);
  or (_08830_, _08754_, _03563_);
  and (_08831_, _08830_, _02501_);
  and (_08832_, _08831_, _08829_);
  and (_08833_, _08751_, _02500_);
  or (_08834_, _08833_, _03174_);
  or (_08835_, _08834_, _08832_);
  and (_08836_, _05257_, _04724_);
  or (_08837_, _08741_, _03178_);
  or (_08838_, _08837_, _08836_);
  and (_08839_, _08838_, _34698_);
  and (_08840_, _08839_, _08835_);
  or (_32495_, _08840_, _08740_);
  and (_08841_, _05390_, _02233_);
  and (_08842_, _08841_, \oc8051_golden_model_1.PC [7]);
  and (_08843_, _08842_, _06197_);
  and (_08844_, _08843_, \oc8051_golden_model_1.PC [11]);
  and (_08845_, _08844_, \oc8051_golden_model_1.PC [12]);
  and (_08846_, _08845_, \oc8051_golden_model_1.PC [13]);
  and (_08847_, _08846_, \oc8051_golden_model_1.PC [14]);
  nor (_08848_, _08847_, \oc8051_golden_model_1.PC [15]);
  and (_08849_, _08842_, \oc8051_golden_model_1.PC [8]);
  and (_08850_, _08849_, \oc8051_golden_model_1.PC [9]);
  and (_08851_, _08850_, \oc8051_golden_model_1.PC [10]);
  and (_08852_, _08851_, \oc8051_golden_model_1.PC [11]);
  and (_08853_, _08852_, \oc8051_golden_model_1.PC [12]);
  and (_08854_, _08853_, \oc8051_golden_model_1.PC [13]);
  and (_08855_, _08854_, \oc8051_golden_model_1.PC [14]);
  and (_08856_, _08855_, \oc8051_golden_model_1.PC [15]);
  nor (_08857_, _08856_, _08848_);
  nor (_08858_, _07258_, _07217_);
  or (_08859_, _08858_, _08857_);
  nor (_08860_, _07950_, _03137_);
  not (_08861_, _08860_);
  and (_08862_, _07889_, _07922_);
  or (_08863_, _08862_, _08857_);
  and (_08864_, _02537_, _02499_);
  not (_08865_, _08864_);
  nor (_08866_, _03127_, _02538_);
  or (_08867_, _08866_, _06227_);
  and (_08868_, _08867_, _08865_);
  not (_08869_, _07858_);
  nor (_08870_, _07850_, _03525_);
  nor (_08871_, _03715_, _03360_);
  and (_08872_, _08871_, _08870_);
  and (_08873_, _08872_, _08869_);
  or (_08874_, _08873_, _08857_);
  and (_08875_, _02532_, _02499_);
  not (_08876_, _08875_);
  nor (_08877_, _03139_, _02533_);
  or (_08878_, _08877_, _06227_);
  and (_08879_, _08878_, _08876_);
  not (_08880_, _08190_);
  nor (_08881_, _06216_, \oc8051_golden_model_1.PC [14]);
  nor (_08882_, _08881_, _06217_);
  and (_08883_, _08882_, _02768_);
  nor (_08884_, _08882_, _02768_);
  nor (_08885_, _08884_, _08883_);
  not (_08886_, _08885_);
  not (_08887_, \oc8051_golden_model_1.PC [13]);
  and (_08888_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_08889_, _08888_, _06196_);
  and (_08890_, _08889_, _05392_);
  and (_08891_, _08890_, \oc8051_golden_model_1.PC [12]);
  nor (_08892_, _08891_, _08887_);
  and (_08893_, _08891_, _08887_);
  or (_08894_, _08893_, _08892_);
  nor (_08895_, _08894_, _02768_);
  and (_08896_, _08894_, _02768_);
  not (_08897_, _08896_);
  nor (_08898_, _06214_, \oc8051_golden_model_1.PC [12]);
  nor (_08899_, _08898_, _06215_);
  and (_08900_, _08899_, _02768_);
  not (_08901_, \oc8051_golden_model_1.PC [11]);
  nor (_08902_, _06213_, _08901_);
  and (_08903_, _06213_, _08901_);
  or (_08904_, _08903_, _08902_);
  and (_08905_, _08904_, _02768_);
  nor (_08906_, _08904_, _02768_);
  nor (_08907_, _06220_, \oc8051_golden_model_1.PC [10]);
  nor (_08908_, _08907_, _06213_);
  and (_08909_, _08908_, _02768_);
  nor (_08910_, _08908_, _02768_);
  nor (_08911_, _08910_, _08909_);
  nor (_08912_, _06219_, \oc8051_golden_model_1.PC [9]);
  nor (_08913_, _08912_, _06220_);
  and (_08914_, _08913_, _02768_);
  nor (_08915_, _08913_, _02768_);
  nor (_08916_, _05392_, \oc8051_golden_model_1.PC [8]);
  nor (_08917_, _08916_, _06219_);
  and (_08918_, _08917_, _02768_);
  and (_08919_, _05394_, _02768_);
  nor (_08920_, _05394_, _02768_);
  and (_08921_, _05389_, _02674_);
  nor (_08922_, _08921_, \oc8051_golden_model_1.PC [6]);
  nor (_08923_, _08922_, _05391_);
  not (_08924_, _08923_);
  nor (_08925_, _08924_, _02932_);
  and (_08926_, _08924_, _02932_);
  nor (_08927_, _08926_, _08925_);
  not (_08928_, _08927_);
  and (_08929_, _02674_, \oc8051_golden_model_1.PC [4]);
  nor (_08930_, _08929_, \oc8051_golden_model_1.PC [5]);
  nor (_08931_, _08930_, _08921_);
  not (_08932_, _08931_);
  nor (_08933_, _08932_, _03215_);
  and (_08934_, _08932_, _03215_);
  nor (_08935_, _02674_, \oc8051_golden_model_1.PC [4]);
  nor (_08936_, _08935_, _08929_);
  not (_08937_, _08936_);
  nor (_08938_, _08937_, _03625_);
  nor (_08939_, _02799_, _02677_);
  and (_08940_, _02799_, _02677_);
  nor (_08941_, _03260_, _02634_);
  nor (_08942_, _03671_, \oc8051_golden_model_1.PC [1]);
  nor (_08943_, _02832_, _02247_);
  and (_08944_, _03671_, \oc8051_golden_model_1.PC [1]);
  nor (_08945_, _08944_, _08942_);
  and (_08946_, _08945_, _08943_);
  nor (_08947_, _08946_, _08942_);
  and (_08948_, _03260_, _02634_);
  nor (_08949_, _08948_, _08941_);
  not (_08950_, _08949_);
  nor (_08951_, _08950_, _08947_);
  nor (_08952_, _08951_, _08941_);
  nor (_08953_, _08952_, _08940_);
  nor (_08954_, _08953_, _08939_);
  and (_08955_, _08937_, _03625_);
  nor (_08956_, _08955_, _08938_);
  not (_08957_, _08956_);
  nor (_08958_, _08957_, _08954_);
  nor (_08959_, _08958_, _08938_);
  nor (_08960_, _08959_, _08934_);
  nor (_08961_, _08960_, _08933_);
  nor (_08962_, _08961_, _08928_);
  nor (_08963_, _08962_, _08925_);
  nor (_08964_, _08963_, _08920_);
  or (_08965_, _08964_, _08919_);
  nor (_08966_, _08917_, _02768_);
  nor (_08967_, _08966_, _08918_);
  and (_08968_, _08967_, _08965_);
  nor (_08969_, _08968_, _08918_);
  nor (_08970_, _08969_, _08915_);
  nor (_08971_, _08970_, _08914_);
  not (_08972_, _08971_);
  and (_08974_, _08972_, _08911_);
  nor (_08975_, _08974_, _08909_);
  nor (_08976_, _08975_, _08906_);
  or (_08977_, _08976_, _08905_);
  nor (_08978_, _08899_, _02768_);
  nor (_08979_, _08978_, _08900_);
  and (_08980_, _08979_, _08977_);
  nor (_08981_, _08980_, _08900_);
  and (_08982_, _08981_, _08897_);
  or (_08983_, _08982_, _08895_);
  nor (_08985_, _08983_, _08886_);
  nor (_08986_, _08985_, _08883_);
  nor (_08987_, _06227_, _02768_);
  and (_08988_, _06227_, _02768_);
  nor (_08989_, _08988_, _08987_);
  and (_08990_, _08989_, _08986_);
  nor (_08991_, _08989_, _08986_);
  or (_08992_, _08991_, _08990_);
  or (_08993_, _08992_, _08880_);
  and (_08994_, _02511_, _02499_);
  or (_08996_, _08190_, _06227_);
  and (_08997_, _08996_, _08994_);
  and (_08998_, _08997_, _08993_);
  or (_08999_, _08992_, _08190_);
  and (_09000_, _02516_, _02499_);
  or (_09001_, _08880_, _06227_);
  and (_09002_, _09001_, _09000_);
  and (_09003_, _09002_, _08999_);
  and (_09004_, _06211_, _02576_);
  and (_09005_, _07426_, _07344_);
  or (_09007_, _09005_, _08857_);
  not (_09008_, _08857_);
  and (_09009_, _02575_, _02980_);
  not (_09010_, _09009_);
  nor (_09011_, _08250_, _06271_);
  and (_09012_, _09011_, _09010_);
  nor (_09013_, _09012_, _09008_);
  nor (_09014_, _06201_, \oc8051_golden_model_1.PC [14]);
  nor (_09015_, _09014_, _06202_);
  and (_09016_, _09015_, _05563_);
  nor (_09018_, _09015_, _05563_);
  nor (_09019_, _09018_, _09016_);
  not (_09020_, _09019_);
  nor (_09021_, _06207_, \oc8051_golden_model_1.PC [13]);
  nor (_09022_, _09021_, _06208_);
  not (_09023_, _09022_);
  nor (_09024_, _09023_, _05311_);
  and (_09025_, _09023_, _05311_);
  nor (_09026_, _06199_, \oc8051_golden_model_1.PC [12]);
  nor (_09027_, _09026_, _06200_);
  and (_09029_, _09027_, _05563_);
  nor (_09030_, _06198_, _08901_);
  and (_09031_, _06198_, _08901_);
  or (_09032_, _09031_, _09030_);
  not (_09033_, _09032_);
  nor (_09034_, _09033_, _05311_);
  and (_09035_, _09033_, _05311_);
  nor (_09036_, _09035_, _09034_);
  nor (_09037_, _06204_, \oc8051_golden_model_1.PC [10]);
  nor (_09038_, _09037_, _06205_);
  not (_09040_, _09038_);
  nor (_09041_, _09040_, _05311_);
  and (_09042_, _09040_, _05311_);
  nor (_09043_, _09042_, _09041_);
  and (_09044_, _09043_, _09036_);
  and (_09045_, _06136_, \oc8051_golden_model_1.PC [8]);
  nor (_09046_, _09045_, \oc8051_golden_model_1.PC [9]);
  nor (_09047_, _09046_, _06204_);
  not (_09048_, _09047_);
  nor (_09049_, _09048_, _05311_);
  and (_09050_, _09048_, _05311_);
  nor (_09051_, _09050_, _09049_);
  nor (_09052_, _06139_, _05311_);
  and (_09053_, _06139_, _05311_);
  and (_09054_, _06134_, _05389_);
  nor (_09055_, _09054_, \oc8051_golden_model_1.PC [6]);
  nor (_09056_, _09055_, _06135_);
  not (_09057_, _09056_);
  nor (_09058_, _09057_, _05598_);
  and (_09059_, _09057_, _05598_);
  nor (_09060_, _09059_, _09058_);
  not (_09061_, _09060_);
  and (_09062_, _06134_, \oc8051_golden_model_1.PC [4]);
  nor (_09063_, _09062_, \oc8051_golden_model_1.PC [5]);
  nor (_09064_, _09063_, _09054_);
  not (_09065_, _09064_);
  nor (_09066_, _09065_, _05661_);
  and (_09067_, _09065_, _05661_);
  nor (_09068_, _06134_, \oc8051_golden_model_1.PC [4]);
  nor (_09069_, _09068_, _09062_);
  not (_09070_, _09069_);
  nor (_09071_, _09070_, _05630_);
  and (_09072_, _02251_, \oc8051_golden_model_1.PC [2]);
  nor (_09073_, _09072_, \oc8051_golden_model_1.PC [3]);
  nor (_09074_, _09073_, _06134_);
  not (_09075_, _09074_);
  nor (_09076_, _09075_, _03120_);
  and (_09077_, _09075_, _03120_);
  nor (_09078_, _02251_, \oc8051_golden_model_1.PC [2]);
  nor (_09079_, _09078_, _09072_);
  not (_09080_, _09079_);
  nor (_09081_, _09080_, _03302_);
  not (_09082_, _02602_);
  nor (_09083_, _03705_, _09082_);
  nor (_09084_, _03492_, \oc8051_golden_model_1.PC [0]);
  and (_09085_, _03705_, _09082_);
  nor (_09086_, _09085_, _09083_);
  and (_09087_, _09086_, _09084_);
  nor (_09088_, _09087_, _09083_);
  and (_09089_, _09080_, _03302_);
  nor (_09090_, _09089_, _09081_);
  not (_09091_, _09090_);
  nor (_09092_, _09091_, _09088_);
  nor (_09093_, _09092_, _09081_);
  nor (_09094_, _09093_, _09077_);
  nor (_09095_, _09094_, _09076_);
  and (_09096_, _09070_, _05630_);
  nor (_09097_, _09096_, _09071_);
  not (_09098_, _09097_);
  nor (_09099_, _09098_, _09095_);
  nor (_09100_, _09099_, _09071_);
  nor (_09101_, _09100_, _09067_);
  nor (_09102_, _09101_, _09066_);
  nor (_09103_, _09102_, _09061_);
  nor (_09104_, _09103_, _09058_);
  nor (_09105_, _09104_, _09053_);
  or (_09106_, _09105_, _09052_);
  nor (_09107_, _06136_, \oc8051_golden_model_1.PC [8]);
  nor (_09108_, _09107_, _09045_);
  not (_09109_, _09108_);
  nor (_09110_, _09109_, _05311_);
  and (_09111_, _09109_, _05311_);
  nor (_09112_, _09111_, _09110_);
  and (_09113_, _09112_, _09106_);
  and (_09114_, _09113_, _09051_);
  and (_09115_, _09114_, _09044_);
  nor (_09116_, _09110_, _09049_);
  not (_09117_, _09116_);
  and (_09118_, _09117_, _09044_);
  or (_09119_, _09118_, _09041_);
  or (_09120_, _09119_, _09115_);
  nor (_09121_, _09120_, _09034_);
  nor (_09122_, _09027_, _05563_);
  nor (_09123_, _09122_, _09029_);
  not (_09124_, _09123_);
  nor (_09125_, _09124_, _09121_);
  nor (_09126_, _09125_, _09029_);
  nor (_09127_, _09126_, _09025_);
  nor (_09128_, _09127_, _09024_);
  nor (_09129_, _09128_, _09020_);
  nor (_09130_, _09129_, _09016_);
  not (_09131_, _06211_);
  and (_09132_, _09131_, _05311_);
  nor (_09133_, _09131_, _05311_);
  nor (_09134_, _09133_, _09132_);
  and (_09135_, _09134_, _09130_);
  nor (_09136_, _09134_, _09130_);
  or (_09137_, _09136_, _09135_);
  and (_09138_, _05984_, _02934_);
  and (_09139_, _06176_, _02799_);
  nor (_09140_, _09139_, _09138_);
  and (_09141_, _06029_, _03261_);
  and (_09142_, _06177_, _03260_);
  nor (_09143_, _09142_, _09141_);
  and (_09144_, _09143_, _09140_);
  and (_09145_, _06174_, _02832_);
  not (_09146_, _09145_);
  and (_09147_, _05893_, _03672_);
  and (_09148_, _06173_, _03671_);
  nor (_09149_, _09148_, _09147_);
  and (_09150_, _09149_, _09146_);
  and (_09151_, _09150_, _09144_);
  and (_09152_, _05938_, _02833_);
  not (_09153_, _09152_);
  nor (_09154_, _05490_, _02858_);
  nor (_09155_, _09154_, _05544_);
  nor (_09156_, _05847_, _02932_);
  and (_09157_, _05847_, _02932_);
  nor (_09158_, _09157_, _09156_);
  and (_09159_, _09158_, _09155_);
  and (_09160_, _06180_, _03215_);
  and (_09161_, _06076_, _04669_);
  nor (_09162_, _09161_, _09160_);
  and (_09163_, _06181_, _03625_);
  and (_09164_, _06121_, _04662_);
  nor (_09165_, _09164_, _09163_);
  and (_09166_, _09165_, _09162_);
  and (_09167_, _09166_, _09159_);
  and (_09168_, _09167_, _09153_);
  and (_09169_, _09168_, _09151_);
  not (_09170_, _09169_);
  and (_09171_, _09170_, _09137_);
  not (_09172_, _03038_);
  and (_09173_, _09169_, _06211_);
  or (_09174_, _09173_, _09172_);
  or (_09175_, _09174_, _09171_);
  and (_09176_, _06227_, _02950_);
  and (_09177_, _02951_, _02556_);
  or (_09178_, _09177_, _06227_);
  and (_09179_, _02890_, _02547_);
  nor (_09180_, _09179_, _07455_);
  and (_09181_, _04837_, _04732_);
  and (_09182_, _09181_, _05494_);
  not (_09183_, _05044_);
  and (_09184_, _05095_, _09183_);
  and (_09185_, _05496_, _09184_);
  nand (_09186_, _09185_, _09182_);
  or (_09187_, _09186_, _06211_);
  not (_09188_, _09186_);
  or (_09189_, _09188_, _09137_);
  and (_09190_, _09189_, _02952_);
  and (_09191_, _09190_, _09187_);
  and (_09192_, _05262_, _05260_);
  and (_09193_, _04038_, _03817_);
  and (_09194_, _04787_, _04623_);
  and (_09195_, _09194_, _09193_);
  and (_09196_, _09195_, _09192_);
  and (_09197_, _09196_, _06227_);
  nand (_09198_, _09195_, _09192_);
  and (_09199_, _09198_, _08992_);
  or (_09200_, _09199_, _05387_);
  or (_09201_, _09200_, _09197_);
  not (_09202_, _07452_);
  and (_09203_, _07440_, _07436_);
  not (_09204_, _07442_);
  nor (_09205_, _02854_, _02432_);
  or (_09206_, _09205_, _02557_);
  and (_09207_, _09206_, _09204_);
  and (_09208_, _09207_, _09203_);
  nand (_09209_, _09208_, _09202_);
  nand (_09210_, _09209_, _09008_);
  nor (_09211_, _02954_, \oc8051_golden_model_1.PC [15]);
  and (_09212_, _09211_, _09204_);
  nor (_09213_, _03825_, _03824_);
  and (_09214_, _09213_, _09206_);
  and (_09215_, _09214_, _09212_);
  nor (_09216_, _09213_, _06227_);
  or (_09217_, _09216_, _09215_);
  nand (_09218_, _09217_, _09203_);
  or (_09219_, _06227_, _07433_);
  and (_09220_, _09219_, _09218_);
  or (_09221_, _09220_, _07452_);
  and (_09222_, _09221_, _02563_);
  and (_09223_, _09222_, _09210_);
  not (_09224_, _02563_);
  nand (_09225_, _06227_, _09224_);
  nand (_09226_, _09225_, _05387_);
  or (_09227_, _09226_, _09223_);
  nor (_09228_, _03818_, _02952_);
  and (_09229_, _09228_, _09227_);
  and (_09230_, _09229_, _09201_);
  or (_09231_, _09230_, _09191_);
  and (_09232_, _09231_, _09180_);
  not (_09233_, _09177_);
  and (_09234_, _09180_, _05402_);
  nor (_09235_, _09234_, _09008_);
  or (_09236_, _09235_, _09233_);
  or (_09237_, _09236_, _09232_);
  and (_09238_, _09237_, _09178_);
  and (_09239_, _07430_, _03849_);
  not (_09240_, _09239_);
  or (_09241_, _09240_, _09238_);
  or (_09242_, _09239_, _08857_);
  and (_09243_, _09242_, _02959_);
  and (_09244_, _09243_, _09241_);
  or (_09245_, _09244_, _09176_);
  and (_09246_, _02885_, _02547_);
  nor (_09247_, _09246_, _07497_);
  and (_09248_, _09247_, _09245_);
  not (_09249_, _09247_);
  and (_09250_, _09249_, _08857_);
  not (_09251_, _02568_);
  nor (_09252_, _02886_, _09251_);
  and (_09253_, _09252_, _02888_);
  not (_09254_, _09253_);
  or (_09255_, _09254_, _09250_);
  or (_09256_, _09255_, _09248_);
  or (_09257_, _09253_, _06227_);
  not (_09258_, _03012_);
  nor (_09259_, _02975_, _02560_);
  and (_09260_, _02842_, _02497_);
  and (_09261_, _09260_, _02879_);
  nor (_09262_, _09261_, _09259_);
  and (_09263_, _09262_, _09258_);
  and (_09264_, _09263_, _09257_);
  and (_09265_, _09264_, _09256_);
  nor (_09266_, _03817_, _02832_);
  not (_09267_, _09266_);
  and (_09268_, _04623_, _02768_);
  nor (_09269_, _09268_, _04624_);
  nor (_09270_, _04787_, _04352_);
  and (_09271_, _04787_, _04352_);
  nor (_09272_, _09271_, _09270_);
  and (_09273_, _09272_, _09269_);
  nor (_09274_, _04896_, _04669_);
  and (_09275_, _04896_, _04669_);
  nor (_09276_, _09275_, _09274_);
  and (_09277_, _05202_, _04662_);
  nor (_09278_, _05202_, _04662_);
  nor (_09279_, _09278_, _09277_);
  and (_09280_, _09279_, _09276_);
  and (_09281_, _09280_, _09273_);
  and (_09282_, _04242_, _02934_);
  nor (_09283_, _04242_, _02934_);
  nor (_09284_, _09283_, _09282_);
  and (_09285_, _04440_, _03261_);
  nor (_09286_, _04440_, _03261_);
  nor (_09287_, _09286_, _09285_);
  and (_09288_, _09287_, _09284_);
  and (_09289_, _03817_, _02832_);
  not (_09290_, _09289_);
  and (_09291_, _04038_, _03672_);
  and (_09292_, _04005_, _03671_);
  nor (_09293_, _09292_, _09291_);
  and (_09294_, _09293_, _09290_);
  and (_09295_, _09294_, _09288_);
  and (_09296_, _09295_, _09281_);
  and (_09297_, _09296_, _09267_);
  nand (_09298_, _09297_, _09131_);
  not (_09299_, _09263_);
  or (_09300_, _09297_, _09137_);
  and (_09301_, _09300_, _09299_);
  and (_09302_, _09301_, _09298_);
  or (_09303_, _09302_, _03038_);
  or (_09304_, _09303_, _09265_);
  and (_09305_, _02879_, _02547_);
  not (_09306_, _09305_);
  nor (_09307_, _03025_, _02966_);
  and (_09308_, _09307_, _09306_);
  and (_09309_, _09308_, _09304_);
  and (_09310_, _09309_, _09175_);
  nand (_09311_, _09305_, _08857_);
  nor (_09312_, _03867_, _04125_);
  and (_09313_, _09312_, _02943_);
  and (_09314_, _09313_, _02983_);
  nand (_09315_, _09314_, _09311_);
  and (_09316_, _02832_, _02549_);
  nor (_09317_, _09316_, _08157_);
  nor (_09318_, _09317_, _08156_);
  nor (_09319_, _08148_, _08149_);
  nor (_09320_, _09319_, _08152_);
  and (_09321_, _08143_, _08146_);
  nor (_09322_, _08139_, _07820_);
  and (_09323_, _09322_, _09321_);
  and (_09324_, _09323_, _09320_);
  and (_09325_, _09324_, _09318_);
  or (_09326_, _09325_, _09137_);
  nand (_09327_, _09325_, _09131_);
  and (_09328_, _09327_, _03025_);
  and (_09329_, _09328_, _09326_);
  and (_09330_, _07724_, _07711_);
  not (_09331_, _07600_);
  and (_09332_, _07613_, _09331_);
  and (_09333_, _09332_, _09330_);
  and (_09334_, _09333_, _07736_);
  or (_09335_, _09334_, _09137_);
  nand (_09336_, _09334_, _09131_);
  and (_09337_, _09336_, _02966_);
  and (_09338_, _09337_, _09335_);
  or (_09339_, _09338_, _09329_);
  or (_09340_, _09339_, _09315_);
  or (_09341_, _09340_, _09310_);
  or (_09342_, _09314_, _06227_);
  and (_09343_, _09342_, _09012_);
  and (_09344_, _09343_, _09341_);
  or (_09345_, _09344_, _09013_);
  not (_09346_, _02987_);
  not (_09347_, _02566_);
  nor (_09348_, _02986_, _09347_);
  and (_09349_, _09348_, _09346_);
  and (_09350_, _09349_, _09345_);
  not (_09351_, _06227_);
  or (_09352_, _09349_, _09351_);
  nand (_09353_, _09352_, _09005_);
  or (_09354_, _09353_, _09350_);
  and (_09355_, _09354_, _09007_);
  or (_09356_, _09355_, _07597_);
  or (_09357_, _07596_, _06227_);
  and (_09358_, _09357_, _02586_);
  and (_09359_, _09358_, _09356_);
  and (_09360_, _08857_, _02585_);
  nor (_09361_, _02874_, _02578_);
  not (_09362_, _09361_);
  or (_09363_, _09362_, _09360_);
  or (_09364_, _09363_, _09359_);
  or (_09365_, _09361_, _06227_);
  and (_09366_, _09365_, _08235_);
  and (_09367_, _09366_, _09364_);
  nand (_09368_, _06211_, _03023_);
  and (_09369_, _06241_, _02856_);
  nand (_09370_, _09369_, _09368_);
  or (_09371_, _09370_, _09367_);
  or (_09372_, _09369_, _06227_);
  and (_09373_, _09372_, _02851_);
  and (_09374_, _09373_, _09371_);
  or (_09375_, _09374_, _09004_);
  nor (_09376_, _06807_, _02548_);
  and (_09377_, _09376_, _09375_);
  not (_09378_, _09376_);
  and (_09379_, _09378_, _08857_);
  nor (_09380_, _02938_, _02521_);
  not (_09381_, _09380_);
  or (_09382_, _09381_, _09379_);
  or (_09383_, _09382_, _09377_);
  and (_09384_, _02520_, _02499_);
  not (_09385_, _09384_);
  or (_09386_, _09380_, _06227_);
  and (_09387_, _09386_, _09385_);
  and (_09388_, _09387_, _09383_);
  and (_09389_, _09384_, _08992_);
  or (_09390_, _09389_, _05562_);
  or (_09391_, _09390_, _09388_);
  or (_09392_, _06227_, _05322_);
  and (_09393_, _09392_, _09391_);
  or (_09394_, _09393_, _03014_);
  or (_09395_, _06211_, _03884_);
  and (_09396_, _09395_, _07783_);
  and (_09397_, _09396_, _09394_);
  and (_09398_, _07782_, _06227_);
  or (_09399_, _09398_, _09397_);
  and (_09400_, _02547_, _02516_);
  not (_09401_, _09400_);
  and (_09402_, _09401_, _09399_);
  not (_09403_, \oc8051_golden_model_1.DPH [0]);
  and (_09404_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_09405_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_09406_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09407_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09408_, _09407_, _09406_);
  not (_09409_, _09408_);
  and (_09410_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09411_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09412_, _09411_, _09410_);
  not (_09413_, _09412_);
  and (_09414_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09415_, _02685_, _02681_);
  nor (_09416_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09417_, _09416_, _09414_);
  not (_09418_, _09417_);
  nor (_09419_, _09418_, _09415_);
  nor (_09420_, _09419_, _09414_);
  nor (_09421_, _09420_, _09413_);
  nor (_09422_, _09421_, _09410_);
  nor (_09423_, _09422_, _09409_);
  nor (_09424_, _09423_, _09406_);
  nor (_09425_, _09424_, _09405_);
  nor (_09426_, _09425_, _09404_);
  nor (_09427_, _09426_, _09403_);
  and (_09428_, _09427_, \oc8051_golden_model_1.DPH [1]);
  and (_09429_, _09428_, \oc8051_golden_model_1.DPH [2]);
  and (_09430_, _09429_, \oc8051_golden_model_1.DPH [3]);
  and (_09431_, _09430_, \oc8051_golden_model_1.DPH [4]);
  and (_09432_, _09431_, \oc8051_golden_model_1.DPH [5]);
  and (_09433_, _09432_, \oc8051_golden_model_1.DPH [6]);
  or (_09434_, _09433_, \oc8051_golden_model_1.DPH [7]);
  nand (_09435_, _09433_, \oc8051_golden_model_1.DPH [7]);
  and (_09436_, _09435_, _09434_);
  and (_09437_, _09436_, _09400_);
  nor (_09438_, _02937_, _02517_);
  not (_09439_, _09438_);
  or (_09440_, _09439_, _09437_);
  or (_09441_, _09440_, _09402_);
  not (_09442_, _09000_);
  or (_09443_, _09438_, _06227_);
  and (_09444_, _09443_, _09442_);
  and (_09445_, _09444_, _09441_);
  or (_09446_, _09445_, _09003_);
  nor (_09447_, _07791_, _07802_);
  and (_09448_, _09447_, _07797_);
  and (_09449_, _09448_, _09446_);
  nor (_09450_, _07812_, _03132_);
  not (_09451_, _09450_);
  nor (_09452_, _09448_, _09008_);
  or (_09453_, _09452_, _09451_);
  or (_09454_, _09453_, _09449_);
  or (_09455_, _09450_, _06227_);
  and (_09456_, _09455_, _05279_);
  and (_09457_, _09456_, _09454_);
  nand (_09458_, _06211_, _03021_);
  nor (_09459_, _03130_, _02512_);
  nand (_09460_, _09459_, _09458_);
  or (_09461_, _09460_, _09457_);
  not (_09462_, _08994_);
  or (_09463_, _09459_, _06227_);
  and (_09464_, _09463_, _09462_);
  and (_09465_, _09464_, _09461_);
  or (_09466_, _09465_, _08998_);
  nor (_09467_, _03011_, _03509_);
  nor (_09468_, _02975_, _03509_);
  nor (_09469_, _09468_, _09467_);
  and (_09470_, _02864_, _02532_);
  nor (_09471_, _09470_, _03512_);
  and (_09472_, _09471_, _07265_);
  and (_09473_, _09472_, _09469_);
  and (_09474_, _09473_, _09466_);
  nor (_09475_, _07836_, _03141_);
  not (_09476_, _09475_);
  nor (_09477_, _09473_, _09008_);
  or (_09478_, _09477_, _09476_);
  or (_09479_, _09478_, _09474_);
  or (_09480_, _09475_, _06227_);
  and (_09481_, _09480_, _05274_);
  and (_09482_, _09481_, _09479_);
  nand (_09483_, _06211_, _03020_);
  nand (_09484_, _09483_, _08877_);
  or (_09485_, _09484_, _09482_);
  and (_09486_, _09485_, _08879_);
  not (_09487_, _08873_);
  or (_09488_, _08992_, \oc8051_golden_model_1.PSW [7]);
  or (_09489_, _06227_, _07319_);
  and (_09490_, _09489_, _08875_);
  and (_09491_, _09490_, _09488_);
  or (_09492_, _09491_, _09487_);
  or (_09493_, _09492_, _09486_);
  and (_09494_, _09493_, _08874_);
  or (_09495_, _09494_, _07867_);
  or (_09496_, _07866_, _06227_);
  and (_09497_, _09496_, _05781_);
  and (_09498_, _09497_, _09495_);
  nand (_09499_, _06211_, _03036_);
  nand (_09500_, _09499_, _08866_);
  or (_09501_, _09500_, _09498_);
  and (_09502_, _09501_, _08868_);
  not (_09503_, _08862_);
  or (_09504_, _08992_, _07319_);
  or (_09505_, _06227_, \oc8051_golden_model_1.PSW [7]);
  and (_09506_, _09505_, _08864_);
  and (_09507_, _09506_, _09504_);
  or (_09508_, _09507_, _09503_);
  or (_09509_, _09508_, _09502_);
  and (_09510_, _09509_, _08863_);
  or (_09511_, _09510_, _08861_);
  or (_09512_, _08860_, _06227_);
  and (_09513_, _09512_, _08030_);
  and (_09514_, _09513_, _09511_);
  and (_09515_, _08857_, _08029_);
  or (_09516_, _09515_, _03148_);
  or (_09517_, _09516_, _09514_);
  nand (_09518_, _04623_, _03148_);
  and (_09519_, _09518_, _09517_);
  or (_09520_, _09519_, _02531_);
  or (_09521_, _06227_, _05792_);
  and (_09522_, _09521_, _03152_);
  and (_09523_, _09522_, _09520_);
  not (_09524_, _08858_);
  and (_09525_, _04652_, _03261_);
  not (_09526_, _09525_);
  and (_09527_, _05355_, \oc8051_golden_model_1.TCON [6]);
  and (_09528_, _05338_, \oc8051_golden_model_1.B [6]);
  nor (_09529_, _09528_, _09527_);
  and (_09530_, _05329_, \oc8051_golden_model_1.PSW [6]);
  not (_09531_, _09530_);
  and (_09532_, _05336_, \oc8051_golden_model_1.IP [6]);
  and (_09533_, _05331_, \oc8051_golden_model_1.ACC [6]);
  nor (_09534_, _09533_, _09532_);
  and (_09535_, _09534_, _09531_);
  and (_09536_, _09535_, _09529_);
  and (_09537_, _05350_, \oc8051_golden_model_1.SCON [6]);
  and (_09538_, _05352_, \oc8051_golden_model_1.IE [6]);
  nor (_09539_, _09538_, _09537_);
  and (_09540_, _04629_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09541_, _05346_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_09542_, _09541_, _09540_);
  and (_09543_, _05344_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09544_, _05357_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09545_, _09544_, _09543_);
  and (_09546_, _09545_, _09542_);
  and (_09547_, _09546_, _09539_);
  and (_09548_, _09547_, _09536_);
  and (_09549_, _09548_, _04788_);
  nor (_09550_, _09549_, _09526_);
  not (_09551_, _04631_);
  and (_09552_, _05350_, \oc8051_golden_model_1.SCON [3]);
  not (_09553_, _09552_);
  and (_09554_, _05352_, \oc8051_golden_model_1.IE [3]);
  and (_09555_, _05338_, \oc8051_golden_model_1.B [3]);
  nor (_09556_, _09555_, _09554_);
  and (_09557_, _09556_, _09553_);
  and (_09558_, _05329_, \oc8051_golden_model_1.PSW [3]);
  and (_09559_, _05331_, \oc8051_golden_model_1.ACC [3]);
  nor (_09560_, _09559_, _09558_);
  and (_09561_, _05355_, \oc8051_golden_model_1.TCON [3]);
  and (_09562_, _05336_, \oc8051_golden_model_1.IP [3]);
  nor (_09563_, _09562_, _09561_);
  and (_09564_, _09563_, _09560_);
  and (_09565_, _09564_, _09557_);
  and (_09566_, _04629_, \oc8051_golden_model_1.P0INREG [3]);
  and (_09567_, _05346_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09568_, _09567_, _09566_);
  and (_09569_, _05344_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09570_, _05357_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_09571_, _09570_, _09569_);
  and (_09572_, _09571_, _09568_);
  and (_09573_, _09572_, _09565_);
  and (_09574_, _09573_, _04945_);
  nor (_09575_, _09574_, _09551_);
  nor (_09576_, _09575_, _09550_);
  and (_09577_, _04647_, _03261_);
  not (_09578_, _09577_);
  and (_09579_, _05336_, \oc8051_golden_model_1.IP [5]);
  and (_09580_, _05331_, \oc8051_golden_model_1.ACC [5]);
  nor (_09581_, _09580_, _09579_);
  and (_09582_, _05329_, \oc8051_golden_model_1.PSW [5]);
  and (_09583_, _05338_, \oc8051_golden_model_1.B [5]);
  nor (_09584_, _09583_, _09582_);
  and (_09585_, _09584_, _09581_);
  and (_09586_, _05350_, \oc8051_golden_model_1.SCON [5]);
  and (_09587_, _05352_, \oc8051_golden_model_1.IE [5]);
  nor (_09588_, _09587_, _09586_);
  and (_09589_, _05355_, \oc8051_golden_model_1.TCON [5]);
  and (_09591_, _05357_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09592_, _09591_, _09589_);
  and (_09593_, _09592_, _09588_);
  and (_09594_, _05344_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09595_, _05346_, \oc8051_golden_model_1.P2INREG [5]);
  and (_09596_, _04629_, \oc8051_golden_model_1.P0INREG [5]);
  or (_09597_, _09596_, _09595_);
  nor (_09598_, _09597_, _09594_);
  and (_09599_, _09598_, _09593_);
  and (_09600_, _09599_, _09585_);
  and (_09601_, _09600_, _04897_);
  nor (_09602_, _09601_, _09578_);
  not (_09603_, _04649_);
  and (_09604_, _05355_, \oc8051_golden_model_1.TCON [1]);
  and (_09605_, _05331_, \oc8051_golden_model_1.ACC [1]);
  nor (_09606_, _09605_, _09604_);
  and (_09607_, _05336_, \oc8051_golden_model_1.IP [1]);
  not (_09608_, _09607_);
  and (_09609_, _05329_, \oc8051_golden_model_1.PSW [1]);
  and (_09610_, _05338_, \oc8051_golden_model_1.B [1]);
  nor (_09612_, _09610_, _09609_);
  and (_09613_, _09612_, _09608_);
  and (_09614_, _09613_, _09606_);
  and (_09615_, _05350_, \oc8051_golden_model_1.SCON [1]);
  and (_09616_, _05352_, \oc8051_golden_model_1.IE [1]);
  nor (_09617_, _09616_, _09615_);
  and (_09618_, _04629_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09619_, _05346_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09620_, _09619_, _09618_);
  and (_09621_, _05344_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09622_, _05357_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09623_, _09622_, _09621_);
  and (_09624_, _09623_, _09620_);
  and (_09625_, _09624_, _09617_);
  and (_09626_, _09625_, _09614_);
  and (_09627_, _09626_, _05045_);
  nor (_09628_, _09627_, _09603_);
  nor (_09629_, _09628_, _09602_);
  and (_09630_, _09629_, _09576_);
  not (_09631_, _04653_);
  and (_09632_, _05355_, \oc8051_golden_model_1.TCON [2]);
  and (_09633_, _05338_, \oc8051_golden_model_1.B [2]);
  nor (_09634_, _09633_, _09632_);
  and (_09635_, _05336_, \oc8051_golden_model_1.IP [2]);
  not (_09636_, _09635_);
  and (_09637_, _05329_, \oc8051_golden_model_1.PSW [2]);
  and (_09638_, _05331_, \oc8051_golden_model_1.ACC [2]);
  nor (_09639_, _09638_, _09637_);
  and (_09640_, _09639_, _09636_);
  and (_09641_, _09640_, _09634_);
  and (_09642_, _05350_, \oc8051_golden_model_1.SCON [2]);
  and (_09643_, _05352_, \oc8051_golden_model_1.IE [2]);
  nor (_09644_, _09643_, _09642_);
  and (_09645_, _04629_, \oc8051_golden_model_1.P0INREG [2]);
  and (_09646_, _05346_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_09647_, _09646_, _09645_);
  and (_09648_, _05344_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09649_, _05357_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_09650_, _09649_, _09648_);
  and (_09651_, _09650_, _09647_);
  and (_09652_, _09651_, _09644_);
  and (_09653_, _09652_, _09641_);
  and (_09654_, _09653_, _05097_);
  nor (_09655_, _09654_, _09631_);
  nor (_09656_, _05363_, _05384_);
  nor (_09657_, _09656_, _09655_);
  not (_09658_, _04667_);
  and (_09659_, _05350_, \oc8051_golden_model_1.SCON [0]);
  and (_09660_, _05352_, \oc8051_golden_model_1.IE [0]);
  nor (_09661_, _09660_, _09659_);
  and (_09662_, _05355_, \oc8051_golden_model_1.TCON [0]);
  and (_09663_, _05357_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09664_, _09663_, _09662_);
  and (_09665_, _09664_, _09661_);
  and (_09666_, _05336_, \oc8051_golden_model_1.IP [0]);
  and (_09667_, _05331_, \oc8051_golden_model_1.ACC [0]);
  nor (_09668_, _09667_, _09666_);
  and (_09669_, _05329_, \oc8051_golden_model_1.PSW [0]);
  and (_09670_, _05338_, \oc8051_golden_model_1.B [0]);
  nor (_09671_, _09670_, _09669_);
  and (_09672_, _09671_, _09668_);
  and (_09673_, _05344_, \oc8051_golden_model_1.P1INREG [0]);
  and (_09674_, _05346_, \oc8051_golden_model_1.P2INREG [0]);
  and (_09675_, _04629_, \oc8051_golden_model_1.P0INREG [0]);
  or (_09676_, _09675_, _09674_);
  nor (_09677_, _09676_, _09673_);
  and (_09678_, _09677_, _09672_);
  and (_09679_, _09678_, _09665_);
  and (_09680_, _09679_, _04997_);
  nor (_09681_, _09680_, _09658_);
  and (_09682_, _04635_, _03261_);
  not (_09683_, _09682_);
  and (_09684_, _05350_, \oc8051_golden_model_1.SCON [4]);
  and (_09685_, _05352_, \oc8051_golden_model_1.IE [4]);
  nor (_09686_, _09685_, _09684_);
  and (_09687_, _05355_, \oc8051_golden_model_1.TCON [4]);
  and (_09688_, _05357_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_09689_, _09688_, _09687_);
  and (_09690_, _09689_, _09686_);
  and (_09691_, _05336_, \oc8051_golden_model_1.IP [4]);
  and (_09692_, _05338_, \oc8051_golden_model_1.B [4]);
  nor (_09693_, _09692_, _09691_);
  and (_09694_, _05329_, \oc8051_golden_model_1.PSW [4]);
  and (_09695_, _05331_, \oc8051_golden_model_1.ACC [4]);
  nor (_09696_, _09695_, _09694_);
  and (_09697_, _09696_, _09693_);
  and (_09698_, _05344_, \oc8051_golden_model_1.P1INREG [4]);
  and (_09699_, _05346_, \oc8051_golden_model_1.P2INREG [4]);
  and (_09700_, _04629_, \oc8051_golden_model_1.P0INREG [4]);
  or (_09701_, _09700_, _09699_);
  nor (_09702_, _09701_, _09698_);
  and (_09703_, _09702_, _09697_);
  and (_09704_, _09703_, _09690_);
  and (_09705_, _09704_, _05203_);
  nor (_09706_, _09705_, _09683_);
  nor (_09707_, _09706_, _09681_);
  and (_09708_, _09707_, _09657_);
  and (_09709_, _09708_, _09630_);
  not (_09710_, _09709_);
  or (_09711_, _09710_, _09137_);
  or (_09712_, _09709_, _06211_);
  and (_09713_, _09712_, _03035_);
  and (_09714_, _09713_, _09711_);
  or (_09715_, _09714_, _09524_);
  or (_09716_, _09715_, _09523_);
  and (_09717_, _09716_, _08859_);
  or (_09718_, _09717_, _08105_);
  or (_09719_, _08104_, _06227_);
  and (_09720_, _09719_, _08136_);
  and (_09721_, _09720_, _09718_);
  and (_09722_, _08857_, _08135_);
  or (_09723_, _09722_, _02897_);
  or (_09724_, _09723_, _09721_);
  nand (_09725_, _04623_, _02897_);
  and (_09726_, _09725_, _09724_);
  or (_09727_, _09726_, _02536_);
  not (_09728_, _02536_);
  or (_09729_, _06227_, _09728_);
  and (_09730_, _09729_, _02896_);
  and (_09731_, _09730_, _09727_);
  or (_09732_, _09709_, _09137_);
  nand (_09733_, _09709_, _09131_);
  and (_09734_, _09733_, _09732_);
  and (_09735_, _09734_, _02895_);
  and (_09736_, _05271_, _03910_);
  not (_09737_, _09736_);
  or (_09738_, _09737_, _09735_);
  or (_09739_, _09738_, _09731_);
  or (_09740_, _09736_, _08857_);
  and (_09741_, _09740_, _03563_);
  and (_09742_, _09741_, _09739_);
  nor (_09743_, _08184_, _08179_);
  not (_09744_, _09743_);
  and (_09745_, _06227_, _03166_);
  or (_09746_, _09745_, _09744_);
  or (_09747_, _09746_, _09742_);
  or (_09748_, _08857_, _09743_);
  and (_09749_, _09748_, _06195_);
  and (_09750_, _09749_, _09747_);
  and (_09751_, _03004_, _02768_);
  or (_09752_, _09751_, _02528_);
  or (_09753_, _09752_, _09750_);
  or (_09754_, _06227_, _02529_);
  and (_09755_, _09754_, _02501_);
  and (_09756_, _09755_, _09753_);
  and (_09757_, _09734_, _02500_);
  and (_09758_, _06154_, _03927_);
  not (_09759_, _09758_);
  or (_09760_, _09759_, _09757_);
  or (_09761_, _09760_, _09756_);
  or (_09762_, _09758_, _08857_);
  and (_09763_, _09762_, _03178_);
  and (_09764_, _09763_, _09761_);
  nor (_09765_, _08208_, _08201_);
  not (_09766_, _09765_);
  and (_09767_, _06227_, _03174_);
  or (_09768_, _09767_, _09766_);
  or (_09769_, _09768_, _09764_);
  not (_09770_, _03006_);
  or (_09771_, _08857_, _09765_);
  and (_09772_, _09771_, _09770_);
  and (_09773_, _09772_, _09769_);
  and (_09774_, _03006_, _02768_);
  or (_09775_, _09774_, _02526_);
  or (_09776_, _09775_, _09773_);
  and (_09777_, _02525_, _02499_);
  not (_09778_, _09777_);
  or (_09779_, _06227_, _02527_);
  and (_09780_, _09779_, _09778_);
  and (_09781_, _09780_, _09776_);
  and (_09782_, _09777_, _08857_);
  or (_09783_, _09782_, _09781_);
  or (_09784_, _09783_, _34702_);
  or (_09785_, _34698_, \oc8051_golden_model_1.PC [15]);
  and (_09786_, _09785_, _36029_);
  and (_32496_, _09786_, _09784_);
  not (_09787_, _08184_);
  or (_09788_, _08169_, _07818_);
  nor (_09789_, _08106_, _07819_);
  and (_09790_, _09789_, _09788_);
  nor (_09791_, _04787_, _04623_);
  and (_09792_, _09791_, _07526_);
  nor (_09793_, _07522_, _05768_);
  or (_09794_, _09793_, _07911_);
  or (_09795_, _09794_, _09792_);
  nor (_09796_, _09795_, _07889_);
  nor (_09797_, _04709_, _07319_);
  and (_09798_, _05771_, _04709_);
  nor (_09799_, _09798_, _09797_);
  nor (_09800_, _09799_, _03131_);
  not (_09801_, _02938_);
  not (_09802_, _04709_);
  nor (_09803_, _05755_, _09802_);
  nor (_09804_, _09803_, _09797_);
  nor (_09805_, _09804_, _02851_);
  nor (_09806_, _09802_, _04623_);
  nor (_09807_, _09806_, _09797_);
  and (_09808_, _09807_, _06793_);
  not (_09809_, _02986_);
  and (_09810_, _05346_, \oc8051_golden_model_1.P2 [2]);
  and (_09811_, _05357_, \oc8051_golden_model_1.P3 [2]);
  nor (_09812_, _09811_, _09810_);
  and (_09813_, _04629_, \oc8051_golden_model_1.P0 [2]);
  and (_09814_, _05344_, \oc8051_golden_model_1.P1 [2]);
  nor (_09815_, _09814_, _09813_);
  and (_09816_, _09815_, _09812_);
  and (_09817_, _09816_, _09644_);
  and (_09818_, _09817_, _09641_);
  and (_09819_, _09818_, _05097_);
  nor (_09820_, _09819_, _09631_);
  and (_09821_, _05346_, \oc8051_golden_model_1.P2 [1]);
  and (_09822_, _05357_, \oc8051_golden_model_1.P3 [1]);
  nor (_09823_, _09822_, _09821_);
  and (_09824_, _04629_, \oc8051_golden_model_1.P0 [1]);
  and (_09825_, _05344_, \oc8051_golden_model_1.P1 [1]);
  nor (_09826_, _09825_, _09824_);
  and (_09827_, _09826_, _09823_);
  and (_09828_, _09827_, _09617_);
  and (_09829_, _09828_, _09614_);
  and (_09830_, _09829_, _05045_);
  nor (_09831_, _09830_, _09603_);
  nor (_09832_, _09831_, _09820_);
  and (_09833_, _04629_, \oc8051_golden_model_1.P0 [4]);
  and (_09834_, _05344_, \oc8051_golden_model_1.P1 [4]);
  nor (_09835_, _09834_, _09833_);
  and (_09836_, _05357_, \oc8051_golden_model_1.P3 [4]);
  and (_09837_, _05346_, \oc8051_golden_model_1.P2 [4]);
  or (_09838_, _09837_, _09836_);
  nor (_09839_, _09838_, _09687_);
  and (_09840_, _09839_, _09697_);
  and (_09841_, _09840_, _09686_);
  and (_09842_, _09841_, _09835_);
  and (_09843_, _09842_, _05203_);
  nor (_09844_, _09683_, _09843_);
  nor (_09845_, _09844_, _05532_);
  and (_09846_, _09845_, _09832_);
  and (_09847_, _04629_, \oc8051_golden_model_1.P0 [0]);
  and (_09848_, _05344_, \oc8051_golden_model_1.P1 [0]);
  nor (_09849_, _09848_, _09847_);
  and (_09850_, _05357_, \oc8051_golden_model_1.P3 [0]);
  and (_09851_, _05346_, \oc8051_golden_model_1.P2 [0]);
  or (_09852_, _09851_, _09850_);
  nor (_09853_, _09852_, _09662_);
  and (_09854_, _09853_, _09672_);
  and (_09855_, _09854_, _09661_);
  and (_09856_, _09855_, _09849_);
  and (_09857_, _09856_, _04997_);
  nor (_09858_, _09857_, _09658_);
  and (_09859_, _05346_, \oc8051_golden_model_1.P2 [6]);
  and (_09860_, _05357_, \oc8051_golden_model_1.P3 [6]);
  nor (_09861_, _09860_, _09859_);
  and (_09862_, _04629_, \oc8051_golden_model_1.P0 [6]);
  and (_09863_, _05344_, \oc8051_golden_model_1.P1 [6]);
  nor (_09864_, _09863_, _09862_);
  and (_09865_, _09864_, _09861_);
  and (_09866_, _09865_, _09539_);
  and (_09867_, _09866_, _09536_);
  and (_09868_, _09867_, _04788_);
  nor (_09869_, _09526_, _09868_);
  nor (_09870_, _09869_, _09858_);
  and (_09871_, _04629_, \oc8051_golden_model_1.P0 [3]);
  and (_09872_, _05357_, \oc8051_golden_model_1.P3 [3]);
  nor (_09873_, _09872_, _09871_);
  and (_09874_, _05344_, \oc8051_golden_model_1.P1 [3]);
  and (_09875_, _05346_, \oc8051_golden_model_1.P2 [3]);
  nor (_09876_, _09875_, _09874_);
  and (_09877_, _09876_, _09873_);
  and (_09878_, _09877_, _09565_);
  and (_09879_, _09878_, _04945_);
  nor (_09880_, _09879_, _09551_);
  and (_09881_, _05357_, \oc8051_golden_model_1.P3 [5]);
  not (_09882_, _09881_);
  and (_09883_, _05346_, \oc8051_golden_model_1.P2 [5]);
  nor (_09884_, _09883_, _09589_);
  and (_09885_, _09884_, _09882_);
  and (_09886_, _04629_, \oc8051_golden_model_1.P0 [5]);
  and (_09887_, _05344_, \oc8051_golden_model_1.P1 [5]);
  nor (_09888_, _09887_, _09886_);
  and (_09889_, _09888_, _09588_);
  and (_09890_, _09889_, _09885_);
  and (_09891_, _09890_, _09585_);
  and (_09892_, _09891_, _04897_);
  nor (_09893_, _09578_, _09892_);
  nor (_09894_, _09893_, _09880_);
  and (_09895_, _09894_, _09870_);
  and (_09896_, _09895_, _09846_);
  nor (_09897_, _09896_, \oc8051_golden_model_1.PSW [7]);
  nor (_09898_, _09897_, _09809_);
  nor (_09899_, _09709_, _09346_);
  not (_09900_, _09308_);
  and (_09901_, _05502_, _04709_);
  nor (_09902_, _09901_, _09797_);
  and (_09903_, _09902_, _02952_);
  and (_09904_, _04709_, \oc8051_golden_model_1.ACC [7]);
  nor (_09905_, _09904_, _09797_);
  nor (_09906_, _09905_, _03826_);
  nor (_09907_, _03825_, _07319_);
  or (_09908_, _09907_, _02952_);
  nor (_09909_, _09908_, _09906_);
  nor (_09910_, _09909_, _07455_);
  not (_09911_, _09910_);
  nor (_09912_, _09911_, _09903_);
  nor (_09913_, _07465_, \oc8051_golden_model_1.PSW [7]);
  not (_09914_, _09913_);
  nor (_09915_, _09914_, _07475_);
  not (_09916_, _09915_);
  and (_09917_, _09916_, _07455_);
  not (_09918_, _02951_);
  or (_09919_, _09179_, _09918_);
  or (_09920_, _09919_, _09917_);
  or (_09921_, _09920_, _09912_);
  nor (_09922_, _05329_, _07319_);
  and (_09923_, _05385_, _05329_);
  nor (_09924_, _09923_, _09922_);
  and (_09925_, _09924_, _02891_);
  and (_09926_, _09807_, _02947_);
  nor (_09927_, _09926_, _09925_);
  and (_09928_, _09927_, _09921_);
  nand (_09929_, _09928_, _02959_);
  or (_09930_, _09905_, _02959_);
  and (_09931_, _09930_, _09929_);
  nor (_09932_, _09931_, _09246_);
  and (_09933_, _09932_, _02888_);
  and (_09934_, _05380_, _05329_);
  nor (_09935_, _09934_, _09922_);
  nor (_09936_, _09935_, _02888_);
  nor (_09937_, _09936_, _09299_);
  not (_09938_, _09937_);
  nor (_09939_, _09938_, _09933_);
  nor (_09940_, _09271_, _09268_);
  nor (_09941_, _09940_, _04624_);
  nor (_09942_, _09275_, _09277_);
  nor (_09943_, _09942_, _09274_);
  and (_09944_, _09943_, _09273_);
  or (_09945_, _09944_, _09941_);
  and (_09946_, _09291_, _09288_);
  and (_09947_, _09284_, _09285_);
  nor (_09948_, _09947_, _09282_);
  not (_09949_, _09948_);
  or (_09950_, _09949_, _09295_);
  or (_09951_, _09950_, _09946_);
  and (_09952_, _09951_, _09281_);
  nor (_09953_, _09952_, _09945_);
  nor (_09954_, _09953_, _09297_);
  nor (_09955_, _09954_, _09263_);
  nor (_09956_, _09955_, _03038_);
  not (_09957_, _09956_);
  nor (_09958_, _09957_, _09939_);
  not (_09959_, _09167_);
  nand (_09960_, _09147_, _09144_);
  and (_09961_, _09140_, _09141_);
  nor (_09962_, _09961_, _09138_);
  not (_09963_, _09962_);
  nor (_09964_, _09963_, _09151_);
  and (_09965_, _09964_, _09960_);
  nor (_09966_, _09965_, _09959_);
  nor (_09967_, _09154_, _09156_);
  nor (_09968_, _09967_, _05544_);
  and (_09969_, _09162_, _09164_);
  or (_09970_, _09969_, _09161_);
  and (_09971_, _09970_, _09159_);
  nor (_09972_, _09971_, _09968_);
  not (_09973_, _09972_);
  nor (_09974_, _09973_, _09966_);
  nor (_09975_, _09169_, _09172_);
  not (_09976_, _09975_);
  nor (_09977_, _09976_, _09974_);
  nor (_09978_, _09977_, _09958_);
  nor (_09979_, _09978_, _09900_);
  nand (_09980_, _09305_, \oc8051_golden_model_1.PSW [7]);
  nor (_09981_, _05528_, \oc8051_golden_model_1.ACC [7]);
  nor (_09982_, _07710_, _07626_);
  nor (_09983_, _09982_, _07625_);
  not (_09984_, _07733_);
  or (_09985_, _09984_, _07683_);
  nor (_09986_, _07682_, _07671_);
  and (_09987_, _09986_, _09985_);
  or (_09988_, _07704_, _07653_);
  or (_09989_, _09988_, _09987_);
  not (_09990_, _07652_);
  and (_09991_, _09330_, _09990_);
  and (_09992_, _09991_, _09989_);
  nor (_09993_, _09992_, _09983_);
  nor (_09994_, _09993_, _07611_);
  or (_09995_, _09994_, _07612_);
  and (_09996_, _09995_, _09331_);
  nor (_09997_, _09996_, _09981_);
  nor (_09998_, _09334_, _03377_);
  not (_09999_, _09998_);
  nor (_10000_, _09999_, _09997_);
  nor (_10001_, _03671_, \oc8051_golden_model_1.ACC [1]);
  and (_10002_, _03671_, \oc8051_golden_model_1.ACC [1]);
  and (_10003_, _02832_, \oc8051_golden_model_1.ACC [0]);
  nor (_10004_, _10003_, _10002_);
  nor (_10005_, _10004_, _10001_);
  not (_10006_, _10005_);
  nand (_10007_, _10006_, _09324_);
  nor (_10008_, _02932_, \oc8051_golden_model_1.ACC [6]);
  not (_10009_, _10008_);
  nor (_10010_, _10009_, _07820_);
  and (_10011_, _02768_, _05768_);
  nor (_10012_, _10011_, _10010_);
  and (_10013_, _03215_, \oc8051_golden_model_1.ACC [5]);
  nor (_10014_, _03215_, \oc8051_golden_model_1.ACC [5]);
  nor (_10015_, _03625_, \oc8051_golden_model_1.ACC [4]);
  nor (_10016_, _10015_, _10014_);
  nor (_10017_, _10016_, _10013_);
  and (_10018_, _10017_, _09322_);
  not (_10019_, _10018_);
  and (_10020_, _10019_, _10012_);
  and (_10021_, _02799_, \oc8051_golden_model_1.ACC [3]);
  nor (_10022_, _02799_, \oc8051_golden_model_1.ACC [3]);
  nor (_10023_, _03260_, \oc8051_golden_model_1.ACC [2]);
  nor (_10024_, _10023_, _10022_);
  nor (_10025_, _10024_, _10021_);
  nand (_10026_, _10025_, _09323_);
  and (_10027_, _10026_, _10020_);
  and (_10028_, _10027_, _10007_);
  not (_10029_, _03025_);
  or (_10030_, _09325_, _10029_);
  nor (_10031_, _10030_, _10028_);
  or (_10032_, _10031_, _09305_);
  or (_10033_, _10032_, _10000_);
  and (_10034_, _10033_, _09980_);
  nor (_10035_, _10034_, _09979_);
  nor (_10036_, _10035_, _02970_);
  nor (_10037_, _09922_, _05533_);
  or (_10038_, _09924_, _02881_);
  nor (_10039_, _10038_, _10037_);
  and (_10040_, _02942_, \oc8051_golden_model_1.PSW [7]);
  and (_10041_, _10040_, _09896_);
  nor (_10042_, _10041_, _10039_);
  not (_10043_, _10042_);
  nor (_10044_, _10043_, _10036_);
  nor (_10045_, _10044_, _06271_);
  and (_10046_, _10045_, _09346_);
  nor (_10047_, _10046_, _09899_);
  nor (_10048_, _10047_, _02986_);
  not (_10049_, _07423_);
  nor (_10050_, _07419_, _07421_);
  and (_10051_, _10050_, _10049_);
  not (_10052_, _10051_);
  or (_10053_, _10052_, _10048_);
  nor (_10054_, _10053_, _09898_);
  and (_10055_, _07529_, _07525_);
  nor (_10056_, _10055_, _07523_);
  not (_10057_, _10056_);
  and (_10058_, _07891_, _07525_);
  not (_10059_, _10058_);
  nor (_10060_, _10059_, _07585_);
  nor (_10061_, _10060_, _10057_);
  nor (_10062_, _10061_, _09792_);
  nor (_10063_, _10062_, _03444_);
  nor (_10064_, _10063_, _07426_);
  nor (_10065_, _10064_, _10054_);
  not (_10066_, _03444_);
  nor (_10067_, _10062_, _10066_);
  nor (_10068_, _10067_, _10065_);
  or (_10069_, _10068_, _03441_);
  and (_10070_, _07358_, _07351_);
  nor (_10071_, _10070_, _07349_);
  and (_10072_, _07924_, _07351_);
  not (_10073_, _10072_);
  nor (_10074_, _10073_, _07412_);
  not (_10075_, _10074_);
  and (_10076_, _10075_, _10071_);
  nor (_10077_, _10076_, _07347_);
  or (_10078_, _10077_, _07344_);
  and (_10079_, _10078_, _02997_);
  and (_10080_, _10079_, _10069_);
  and (_10081_, _07972_, _07967_);
  nor (_10082_, _10081_, _07965_);
  not (_10083_, _10082_);
  nor (_10084_, _07986_, _07981_);
  nor (_10085_, _10084_, _07980_);
  and (_10086_, _07988_, _07982_);
  and (_10087_, _08000_, _07994_);
  and (_10088_, _08008_, _02549_);
  nor (_10089_, _10088_, _08004_);
  or (_10090_, _10089_, _08005_);
  and (_10091_, _10090_, _10087_);
  and (_10092_, _07998_, _07994_);
  or (_10093_, _10092_, _07992_);
  nor (_10094_, _10093_, _10091_);
  not (_10095_, _10094_);
  and (_10096_, _10095_, _10086_);
  nor (_10097_, _10096_, _10085_);
  and (_10098_, _07973_, _07967_);
  not (_10099_, _10098_);
  nor (_10100_, _10099_, _10097_);
  nor (_10101_, _10100_, _10083_);
  not (_10102_, _05528_);
  and (_10103_, _07961_, _10102_);
  or (_10104_, _10103_, _02997_);
  or (_10105_, _10104_, _10101_);
  and (_10106_, _10105_, _07277_);
  not (_10107_, _10106_);
  nor (_10108_, _10107_, _10080_);
  and (_10109_, _07280_, _04703_);
  and (_10110_, _07293_, _07287_);
  and (_10111_, _10110_, _07334_);
  not (_10112_, _10111_);
  and (_10113_, _10110_, _07336_);
  not (_10114_, _10113_);
  and (_10115_, _07291_, _07287_);
  nor (_10116_, _10115_, _07285_);
  and (_10117_, _10116_, _10114_);
  and (_10118_, _10117_, _10112_);
  nor (_10119_, _10118_, _10109_);
  nor (_10120_, _10119_, _07277_);
  nor (_10121_, _10120_, _06793_);
  not (_10122_, _10121_);
  nor (_10123_, _10122_, _10108_);
  nor (_10124_, _10123_, _09808_);
  nor (_10125_, _10124_, _02855_);
  and (_10126_, _05490_, _04709_);
  nor (_10127_, _09797_, _02856_);
  not (_10128_, _10127_);
  nor (_10129_, _10128_, _10126_);
  nor (_10130_, _10129_, _02576_);
  not (_10131_, _10130_);
  nor (_10132_, _10131_, _10125_);
  nor (_10133_, _10132_, _09805_);
  nor (_10134_, _10133_, _06807_);
  and (_10135_, _10134_, _09801_);
  nor (_10136_, _09896_, _07319_);
  and (_10137_, _10136_, _02938_);
  or (_10138_, _10137_, _03014_);
  or (_10139_, _10138_, _10135_);
  and (_10140_, _05563_, _04709_);
  nor (_10141_, _10140_, _09797_);
  nand (_10142_, _10141_, _03014_);
  and (_10143_, _10142_, _10139_);
  nor (_10144_, _10143_, _02937_);
  and (_10145_, _09896_, _07319_);
  and (_10146_, _10145_, _02937_);
  nor (_10147_, _10146_, _10144_);
  and (_10148_, _10147_, _05279_);
  and (_10149_, _05314_, _04709_);
  nor (_10150_, _10149_, _09797_);
  nor (_10151_, _10150_, _05279_);
  or (_10152_, _10151_, _10148_);
  and (_10153_, _10152_, _03131_);
  nor (_10154_, _10153_, _09800_);
  nor (_10155_, _10154_, _03020_);
  nor (_10156_, _09797_, _04733_);
  not (_10157_, _10156_);
  nor (_10158_, _10141_, _05274_);
  and (_10159_, _10158_, _10157_);
  nor (_10160_, _10159_, _10155_);
  nor (_10161_, _10160_, _03139_);
  nor (_10162_, _09905_, _03140_);
  and (_10163_, _10162_, _10157_);
  or (_10164_, _10163_, _10161_);
  and (_10165_, _10164_, _05781_);
  nor (_10166_, _05312_, _09802_);
  nor (_10167_, _10166_, _09797_);
  nor (_10168_, _10167_, _05781_);
  or (_10169_, _10168_, _10165_);
  and (_10170_, _10169_, _05786_);
  not (_10171_, _07889_);
  nor (_10172_, _05770_, _09802_);
  nor (_10173_, _10172_, _09797_);
  nor (_10174_, _10173_, _05786_);
  nor (_10175_, _10174_, _10171_);
  not (_10176_, _10175_);
  nor (_10177_, _10176_, _10170_);
  nor (_10178_, _10177_, _09796_);
  nor (_10179_, _10178_, _07917_);
  and (_10180_, _07348_, \oc8051_golden_model_1.ACC [7]);
  nor (_10181_, _10180_, _07944_);
  nor (_10182_, _07347_, _07922_);
  and (_10183_, _10182_, _10181_);
  nor (_10184_, _10183_, _03137_);
  not (_10185_, _10184_);
  nor (_10186_, _10185_, _10179_);
  nor (_10187_, _07964_, _05768_);
  nor (_10188_, _10187_, _08023_);
  nor (_10189_, _07950_, _10103_);
  nand (_10190_, _10189_, _10188_);
  and (_10191_, _10190_, _08861_);
  nor (_10192_, _10191_, _10186_);
  nor (_10193_, _07284_, _05768_);
  nor (_10194_, _10193_, _08053_);
  and (_10195_, _07279_, _04704_);
  nor (_10196_, _10195_, _08031_);
  and (_10197_, _10196_, _10194_);
  or (_10198_, _10197_, _08029_);
  nor (_10199_, _10198_, _10192_);
  and (_10200_, _08029_, \oc8051_golden_model_1.ACC [7]);
  nor (_10201_, _10200_, _07258_);
  not (_10202_, _10201_);
  nor (_10203_, _10202_, _10199_);
  nor (_10204_, _07221_, _07219_);
  nor (_10205_, _10204_, _07218_);
  and (_10206_, _07253_, _07220_);
  or (_10207_, _10206_, _07259_);
  nor (_10208_, _10207_, _10205_);
  nor (_10209_, _10208_, _10203_);
  nor (_10210_, _10209_, _07217_);
  not (_10211_, _07266_);
  nor (_10212_, _08096_, _07807_);
  nor (_10213_, _10212_, _08064_);
  and (_10214_, _10213_, _10211_);
  or (_10215_, _10214_, _02899_);
  nor (_10216_, _10215_, _10210_);
  not (_10217_, _07598_);
  not (_10218_, _07599_);
  and (_10219_, _08128_, _10218_);
  nor (_10220_, _10219_, _02901_);
  nand (_10221_, _10220_, _10217_);
  and (_10222_, _10221_, _08106_);
  not (_10223_, _10222_);
  nor (_10224_, _10223_, _10216_);
  nor (_10225_, _10224_, _09790_);
  and (_10226_, _10225_, _03563_);
  nor (_10227_, _09902_, _03563_);
  or (_10228_, _10227_, _10226_);
  and (_10229_, _10228_, _09787_);
  and (_10230_, _08184_, \oc8051_golden_model_1.ACC [0]);
  or (_10231_, _10230_, _10229_);
  and (_10232_, _10231_, _02501_);
  nor (_10233_, _09935_, _02501_);
  or (_10234_, _10233_, _10232_);
  nor (_10235_, _10234_, _03174_);
  and (_10236_, _05257_, _04709_);
  nor (_10237_, _10236_, _09797_);
  and (_10238_, _10237_, _03174_);
  nor (_10239_, _10238_, _10235_);
  or (_10240_, _10239_, _34702_);
  or (_10241_, _34698_, \oc8051_golden_model_1.PSW [7]);
  and (_10242_, _10241_, _36029_);
  and (_32497_, _10242_, _10240_);
  and (_32498_, \oc8051_golden_model_1.PCON [7], _36029_);
  and (_32499_, \oc8051_golden_model_1.SBUF [7], _36029_);
  and (_32500_, \oc8051_golden_model_1.SCON [7], _36029_);
  and (_10243_, _04248_, \oc8051_golden_model_1.SP [4]);
  and (_10244_, _10243_, \oc8051_golden_model_1.SP [5]);
  and (_10245_, _10244_, \oc8051_golden_model_1.SP [6]);
  nor (_10246_, _10245_, \oc8051_golden_model_1.SP [7]);
  and (_10247_, _10245_, \oc8051_golden_model_1.SP [7]);
  nor (_10248_, _10247_, _10246_);
  nor (_10249_, _10248_, _03916_);
  not (_10250_, _03148_);
  not (_10251_, _08877_);
  not (_10252_, \oc8051_golden_model_1.SP [7]);
  nor (_10253_, _04650_, _10252_);
  and (_10254_, _05771_, _04650_);
  nor (_10255_, _10254_, _10253_);
  nor (_10256_, _10255_, _03131_);
  nor (_10257_, _10248_, _04126_);
  and (_10258_, _05502_, _04650_);
  nor (_10259_, _10258_, _10253_);
  and (_10260_, _10259_, _02952_);
  and (_10261_, _04650_, \oc8051_golden_model_1.ACC [7]);
  nor (_10262_, _10261_, _10253_);
  or (_10263_, _10262_, _03826_);
  nand (_10264_, _09213_, \oc8051_golden_model_1.SP [7]);
  not (_10265_, _10248_);
  nor (_10266_, _10265_, _02558_);
  nor (_10267_, _10266_, _02952_);
  and (_10268_, _10267_, _10264_);
  and (_10269_, _10268_, _10263_);
  nor (_10270_, _10269_, _05382_);
  not (_10271_, _10270_);
  nor (_10272_, _10271_, _10260_);
  nor (_10273_, _10265_, _02556_);
  or (_10274_, _10273_, _02947_);
  nor (_10275_, _10274_, _10272_);
  not (_10276_, \oc8051_golden_model_1.SP [6]);
  not (_10277_, \oc8051_golden_model_1.SP [5]);
  not (_10278_, \oc8051_golden_model_1.SP [4]);
  and (_10279_, _05407_, _10278_);
  and (_10280_, _10279_, _10277_);
  and (_10281_, _10280_, _10276_);
  and (_10282_, _10281_, _02877_);
  nor (_10283_, _10282_, _10252_);
  and (_10284_, _10282_, _10252_);
  nor (_10285_, _10284_, _10283_);
  and (_10286_, _10285_, _02947_);
  nor (_10287_, _10286_, _10275_);
  and (_10288_, _10287_, _02959_);
  nor (_10289_, _10262_, _02959_);
  or (_10290_, _10289_, _10288_);
  and (_10291_, _10290_, _03947_);
  not (_10292_, _04126_);
  and (_10293_, _10245_, \oc8051_golden_model_1.SP [0]);
  nor (_10294_, _10293_, _10252_);
  and (_10295_, _10293_, _10252_);
  nor (_10296_, _10295_, _10294_);
  nor (_10297_, _10296_, _03947_);
  nor (_10298_, _10297_, _10292_);
  not (_10299_, _10298_);
  nor (_10300_, _10299_, _10291_);
  nor (_10301_, _10300_, _10257_);
  nor (_10302_, _02865_, _02844_);
  not (_10303_, _10302_);
  nor (_10304_, _10303_, _06240_);
  not (_10305_, _10304_);
  nor (_10306_, _10305_, _10301_);
  not (_10307_, _04650_);
  nor (_10308_, _10307_, _04623_);
  nor (_10309_, _10308_, _10253_);
  and (_10310_, _10309_, _10305_);
  nor (_10311_, _10310_, _02863_);
  not (_10312_, _10311_);
  nor (_10313_, _10312_, _10306_);
  not (_10314_, _02863_);
  nor (_10315_, _10309_, _10314_);
  nor (_10316_, _10315_, _02855_);
  not (_10317_, _10316_);
  nor (_10318_, _10317_, _10313_);
  and (_10319_, _05490_, _04650_);
  nor (_10320_, _10253_, _02856_);
  not (_10321_, _10320_);
  nor (_10322_, _10321_, _10319_);
  nor (_10323_, _10322_, _02576_);
  not (_10324_, _10323_);
  nor (_10325_, _10324_, _10318_);
  nor (_10326_, _05755_, _10307_);
  nor (_10327_, _10326_, _10253_);
  nor (_10328_, _10327_, _02851_);
  or (_10329_, _10328_, _03014_);
  or (_10330_, _10329_, _10325_);
  and (_10331_, _05563_, _04650_);
  nor (_10332_, _10331_, _10253_);
  nand (_10333_, _10332_, _03014_);
  and (_10334_, _10333_, _10330_);
  nor (_10335_, _10334_, _02517_);
  and (_10336_, _10265_, _02517_);
  nor (_10337_, _10336_, _10335_);
  and (_10338_, _10337_, _05279_);
  and (_10339_, _05314_, _04650_);
  nor (_10340_, _10339_, _10253_);
  nor (_10341_, _10340_, _05279_);
  or (_10342_, _10341_, _10338_);
  and (_10343_, _10342_, _03131_);
  nor (_10344_, _10343_, _10256_);
  nor (_10345_, _10344_, _03020_);
  not (_10346_, _10253_);
  and (_10347_, _10346_, _04732_);
  or (_10348_, _10347_, _05274_);
  nor (_10349_, _10348_, _10332_);
  nor (_10350_, _10349_, _10345_);
  nor (_10351_, _10350_, _10251_);
  and (_10352_, _10248_, _02533_);
  nor (_10353_, _10352_, _03036_);
  or (_10354_, _10262_, _03140_);
  or (_10355_, _10354_, _10347_);
  nand (_10356_, _10355_, _10353_);
  nor (_10357_, _10356_, _10351_);
  nor (_10358_, _05312_, _10307_);
  or (_10359_, _10253_, _05781_);
  nor (_10360_, _10359_, _10358_);
  nor (_10361_, _10360_, _10357_);
  and (_10362_, _10361_, _05786_);
  nor (_10363_, _05770_, _10307_);
  nor (_10364_, _10363_, _10253_);
  nor (_10365_, _10364_, _05786_);
  or (_10366_, _10365_, _10362_);
  and (_10367_, _10366_, _10250_);
  nor (_10368_, _10281_, \oc8051_golden_model_1.SP [7]);
  and (_10369_, _10281_, \oc8051_golden_model_1.SP [7]);
  nor (_10370_, _10369_, _10368_);
  and (_10371_, _10370_, _03148_);
  or (_10372_, _10371_, _02531_);
  nor (_10373_, _10372_, _10367_);
  and (_10374_, _10265_, _02531_);
  nor (_10375_, _10374_, _10373_);
  and (_10376_, _10375_, _02898_);
  and (_10377_, _10370_, _02897_);
  or (_10378_, _10377_, _10376_);
  and (_10379_, _10378_, _03563_);
  nor (_10380_, _10259_, _03563_);
  nor (_10381_, _10380_, _04159_);
  not (_10382_, _10381_);
  nor (_10383_, _10382_, _10379_);
  nor (_10384_, _10383_, _10249_);
  and (_10385_, _10384_, _03178_);
  and (_10386_, _05257_, _04650_);
  nor (_10387_, _10386_, _10253_);
  nor (_10388_, _10387_, _03178_);
  or (_10389_, _10388_, _10385_);
  or (_10390_, _10389_, _34702_);
  or (_10391_, _34698_, \oc8051_golden_model_1.SP [7]);
  and (_10392_, _10391_, _36029_);
  and (_32501_, _10392_, _10390_);
  and (_32503_, \oc8051_golden_model_1.TCON [7], _36029_);
  and (_32504_, \oc8051_golden_model_1.TH0 [7], _36029_);
  and (_32505_, \oc8051_golden_model_1.TH1 [7], _36029_);
  and (_32506_, \oc8051_golden_model_1.TL0 [7], _36029_);
  and (_32507_, \oc8051_golden_model_1.TL1 [7], _36029_);
  and (_32508_, \oc8051_golden_model_1.TMOD [7], _36029_);
  and (_10393_, _34702_, \oc8051_golden_model_1.P0INREG [7]);
  or (_10394_, _10393_, _00711_);
  and (_32509_, _10394_, _36029_);
  and (_10395_, _34702_, \oc8051_golden_model_1.P1INREG [7]);
  or (_10396_, _10395_, _00455_);
  and (_32510_, _10396_, _36029_);
  and (_10397_, _34702_, \oc8051_golden_model_1.P2INREG [7]);
  or (_10398_, _10397_, _00592_);
  and (_32512_, _10398_, _36029_);
  and (_10399_, _34702_, \oc8051_golden_model_1.P3INREG [7]);
  or (_10400_, _10399_, _00671_);
  and (_32513_, _10400_, _36029_);
  nor (_10401_, _04558_, _04535_);
  nor (_10402_, _10401_, _04564_);
  and (_10403_, _10402_, _04557_);
  nor (_10404_, _04187_, _03932_);
  nor (_10405_, _10404_, _04188_);
  and (_10406_, _10405_, _10403_);
  or (_10407_, _10406_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_10408_, _04550_, _04104_);
  not (_10409_, _10408_);
  not (_10410_, _03939_);
  and (_10411_, _10408_, _04543_);
  and (_10412_, _10408_, _04546_);
  or (_10413_, _10412_, _10411_);
  or (_10414_, _10413_, _10410_);
  or (_10415_, _10414_, _10409_);
  and (_10416_, _10415_, _10407_);
  nor (_10417_, _04558_, _04103_);
  nor (_10418_, _10417_, _04559_);
  nand (_10419_, _10418_, _10403_);
  and (_10420_, _02528_, \oc8051_golden_model_1.PC [0]);
  and (_10421_, _05044_, _02549_);
  nand (_10422_, _10421_, _05787_);
  and (_10423_, _05044_, _03492_);
  nor (_10424_, _05044_, _03492_);
  nor (_10425_, _10424_, _10423_);
  and (_10426_, _10425_, _05280_);
  or (_10427_, _05551_, _03817_);
  nand (_10428_, _07700_, _02984_);
  nand (_10429_, _09857_, _09658_);
  nand (_10430_, _10429_, _02883_);
  nor (_10431_, _10430_, _09858_);
  and (_10432_, _05044_, _03822_);
  not (_10433_, _05387_);
  nand (_10434_, _10433_, _03817_);
  nor (_10435_, _02558_, _02247_);
  and (_10436_, _02558_, \oc8051_golden_model_1.ACC [0]);
  nor (_10437_, _10436_, _10435_);
  and (_10438_, _10437_, _05387_);
  nor (_10439_, _10438_, _03822_);
  and (_10440_, _10439_, _10434_);
  or (_10441_, _10440_, _10432_);
  and (_10442_, _10441_, _05383_);
  and (_10443_, _10429_, _02894_);
  or (_10444_, _10443_, _10442_);
  and (_10445_, _10444_, _02556_);
  nor (_10446_, _02556_, _02247_);
  or (_10447_, _03845_, _10446_);
  or (_10448_, _10447_, _10445_);
  or (_10449_, _04256_, _03817_);
  and (_10450_, _10449_, _05368_);
  and (_10451_, _10450_, _10448_);
  nor (_10452_, _09857_, _04667_);
  and (_10453_, _10452_, _03853_);
  or (_10454_, _10453_, _02886_);
  or (_10455_, _10454_, _10451_);
  nand (_10456_, _07700_, _02886_);
  and (_10457_, _10456_, _02884_);
  and (_10458_, _10457_, _10455_);
  or (_10459_, _10458_, _10431_);
  and (_10460_, _10459_, _02561_);
  or (_10461_, _02561_, _02247_);
  nand (_10462_, _02983_, _10461_);
  or (_10463_, _10462_, _10460_);
  and (_10464_, _10463_, _10428_);
  or (_10465_, _10464_, _03867_);
  and (_10466_, _06174_, _02858_);
  nand (_10467_, _07699_, _03867_);
  or (_10468_, _10467_, _10466_);
  and (_10469_, _10468_, _10465_);
  or (_10470_, _10469_, _03626_);
  nor (_10471_, _09680_, _04667_);
  and (_10472_, _04667_, \oc8051_golden_model_1.PSW [7]);
  nor (_10473_, _10472_, _10471_);
  nand (_10474_, _10473_, _03626_);
  and (_10475_, _10474_, _05325_);
  and (_10476_, _10475_, _10470_);
  nand (_10477_, _02578_, \oc8051_golden_model_1.PC [0]);
  nand (_10478_, _05551_, _10477_);
  or (_10479_, _10478_, _10476_);
  and (_10480_, _10479_, _10427_);
  or (_10481_, _10480_, _02857_);
  or (_10482_, _06174_, _05558_);
  and (_10483_, _10482_, _02853_);
  and (_10484_, _10483_, _10481_);
  and (_10485_, _05311_, _03817_);
  and (_10486_, _05749_, \oc8051_golden_model_1.DPL [0]);
  and (_10487_, _05677_, \oc8051_golden_model_1.TL0 [0]);
  nor (_10488_, _10487_, _10486_);
  and (_10489_, _05681_, \oc8051_golden_model_1.TH1 [0]);
  and (_10490_, _05672_, \oc8051_golden_model_1.DPH [0]);
  nor (_10491_, _10490_, _10489_);
  and (_10492_, _10491_, _10488_);
  and (_10493_, _05689_, \oc8051_golden_model_1.IP [0]);
  and (_10494_, _05694_, \oc8051_golden_model_1.B [0]);
  nor (_10495_, _10494_, _10493_);
  and (_10496_, _05699_, \oc8051_golden_model_1.PSW [0]);
  and (_10497_, _05703_, \oc8051_golden_model_1.ACC [0]);
  nor (_10498_, _10497_, _10496_);
  and (_10499_, _10498_, _10495_);
  and (_10500_, _05708_, \oc8051_golden_model_1.IE [0]);
  and (_10501_, _05712_, \oc8051_golden_model_1.SBUF [0]);
  and (_10502_, _05714_, \oc8051_golden_model_1.SCON [0]);
  or (_10503_, _10502_, _10501_);
  nor (_10504_, _10503_, _10500_);
  and (_10505_, _10504_, _10499_);
  and (_10506_, _10505_, _10492_);
  and (_10507_, _05720_, \oc8051_golden_model_1.TH0 [0]);
  and (_10508_, _05722_, \oc8051_golden_model_1.TL1 [0]);
  nor (_10509_, _10508_, _10507_);
  and (_10510_, _05725_, \oc8051_golden_model_1.TCON [0]);
  and (_10511_, _05729_, \oc8051_golden_model_1.PCON [0]);
  nor (_10512_, _10511_, _10510_);
  and (_10513_, _10512_, _10509_);
  and (_10514_, _05733_, \oc8051_golden_model_1.P1INREG [0]);
  not (_10515_, _10514_);
  and (_10516_, _05736_, \oc8051_golden_model_1.P0INREG [0]);
  not (_10517_, _10516_);
  and (_10518_, _05739_, \oc8051_golden_model_1.P2INREG [0]);
  and (_10519_, _05741_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_10520_, _10519_, _10518_);
  and (_10521_, _10520_, _10517_);
  and (_10522_, _10521_, _10515_);
  and (_10523_, _05747_, \oc8051_golden_model_1.SP [0]);
  and (_10524_, _05667_, \oc8051_golden_model_1.TMOD [0]);
  nor (_10525_, _10524_, _10523_);
  and (_10526_, _10525_, _10522_);
  and (_10527_, _10526_, _10513_);
  and (_10528_, _10527_, _10506_);
  not (_10529_, _10528_);
  nor (_10530_, _10529_, _10485_);
  nor (_10531_, _10530_, _02853_);
  or (_10532_, _10531_, _05562_);
  or (_10533_, _10532_, _10484_);
  and (_10534_, _05562_, _02832_);
  nor (_10535_, _10534_, _03885_);
  and (_10536_, _10535_, _10533_);
  and (_10537_, _03885_, _05566_);
  or (_10538_, _10537_, _02517_);
  or (_10539_, _10538_, _10536_);
  and (_10540_, _02517_, _02247_);
  nor (_10541_, _10540_, _05280_);
  and (_10542_, _10541_, _10539_);
  or (_10543_, _10542_, _10426_);
  and (_10544_, _10543_, _05278_);
  nor (_10545_, _05044_, _02549_);
  nor (_10546_, _10545_, _10421_);
  and (_10547_, _10546_, _05277_);
  or (_10548_, _10547_, _10544_);
  and (_10549_, _10548_, _05276_);
  and (_10550_, _10424_, _05275_);
  or (_10551_, _10550_, _10549_);
  and (_10552_, _10551_, _05273_);
  and (_10553_, _10545_, _03891_);
  or (_10554_, _10553_, _02533_);
  or (_10555_, _10554_, _10552_);
  and (_10556_, _02533_, _02247_);
  nor (_10557_, _10556_, _05782_);
  and (_10558_, _10557_, _10555_);
  nor (_10559_, _10423_, _05788_);
  or (_10560_, _10559_, _05787_);
  or (_10561_, _10560_, _10558_);
  and (_10562_, _10561_, _10422_);
  or (_10563_, _10562_, _02531_);
  nand (_10564_, _02531_, _02247_);
  and (_10565_, _10564_, _05271_);
  and (_10566_, _10565_, _10563_);
  nor (_10567_, _05271_, _03817_);
  or (_10568_, _10567_, _10566_);
  and (_10569_, _10568_, _03910_);
  and (_10570_, _05938_, _03909_);
  or (_10571_, _10570_, _03908_);
  or (_10572_, _10571_, _10569_);
  or (_10573_, _05044_, _05801_);
  and (_10574_, _10573_, _03916_);
  and (_10575_, _10574_, _10572_);
  and (_10576_, _03004_, _02247_);
  or (_10577_, _10576_, _10575_);
  or (_10578_, _10577_, _10420_);
  or (_10579_, _10578_, _03627_);
  or (_10580_, _10471_, _03936_);
  and (_10581_, _10580_, _06154_);
  and (_10582_, _10581_, _10579_);
  nor (_10583_, _06154_, _03817_);
  or (_10584_, _10583_, _10582_);
  and (_10585_, _10584_, _03927_);
  and (_10586_, _05938_, _03926_);
  or (_10587_, _10586_, _03925_);
  or (_10588_, _10587_, _10585_);
  or (_10589_, _05044_, _04176_);
  and (_10590_, _10589_, _04557_);
  and (_10591_, _10590_, _10588_);
  or (_10592_, _10591_, _10419_);
  and (_10593_, _10592_, _10416_);
  and (_10594_, _04551_, _04543_);
  nor (_10595_, _10594_, _04552_);
  and (_10596_, _04551_, _03939_);
  and (_10597_, _10596_, _10595_);
  nand (_10598_, _09109_, _03004_);
  or (_10599_, _08917_, _03004_);
  and (_10600_, _10599_, _10598_);
  and (_10601_, _10600_, _04551_);
  and (_10602_, _10601_, _10597_);
  or (_32540_, _10602_, _10593_);
  or (_10603_, _10406_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_10604_, _10603_, _10415_);
  or (_10605_, _06175_, _05939_);
  and (_10606_, _10605_, _03909_);
  nand (_10607_, _05269_, _02497_);
  nor (_10608_, _06161_, _05261_);
  nor (_10609_, _10608_, _10607_);
  and (_10610_, _05095_, _03705_);
  nor (_10611_, _05095_, _03705_);
  nor (_10612_, _10611_, _10610_);
  and (_10613_, _10612_, _05280_);
  or (_10614_, _04005_, _05551_);
  nand (_10615_, _07681_, _02984_);
  not (_10616_, _09831_);
  nand (_10617_, _09830_, _09603_);
  and (_10618_, _10617_, _02883_);
  and (_10619_, _10618_, _10616_);
  nor (_10620_, _09830_, _04649_);
  or (_10621_, _10620_, _05368_);
  nor (_10622_, _05495_, _05096_);
  nand (_10623_, _10622_, _03822_);
  nand (_10624_, _10608_, _10433_);
  nor (_10625_, _02558_, \oc8051_golden_model_1.PC [1]);
  and (_10626_, _02558_, \oc8051_golden_model_1.ACC [1]);
  nor (_10627_, _10626_, _10625_);
  nand (_10628_, _10627_, _05387_);
  and (_10629_, _10628_, _10624_);
  or (_10630_, _10629_, _03822_);
  and (_10631_, _10630_, _10623_);
  or (_10632_, _10631_, _02894_);
  or (_10633_, _10617_, _05383_);
  and (_10634_, _10633_, _10632_);
  or (_10635_, _10634_, _05382_);
  nor (_10636_, _02556_, _02218_);
  nor (_10637_, _10636_, _03845_);
  and (_10638_, _10637_, _10635_);
  and (_10639_, _04005_, _03845_);
  or (_10640_, _10639_, _03853_);
  or (_10641_, _10640_, _10638_);
  and (_10642_, _10641_, _10621_);
  or (_10643_, _10642_, _02886_);
  nand (_10644_, _07681_, _02886_);
  and (_10645_, _10644_, _02884_);
  and (_10646_, _10645_, _10643_);
  or (_10647_, _10646_, _10619_);
  and (_10648_, _10647_, _02561_);
  or (_10649_, _02561_, \oc8051_golden_model_1.PC [1]);
  nand (_10650_, _02983_, _10649_);
  or (_10651_, _10650_, _10648_);
  and (_10652_, _10651_, _10615_);
  or (_10653_, _10652_, _03867_);
  and (_10654_, _06173_, _02858_);
  nand (_10655_, _07680_, _03867_);
  or (_10656_, _10655_, _10654_);
  and (_10657_, _10656_, _10653_);
  or (_10658_, _10657_, _03626_);
  nor (_10659_, _09627_, _04649_);
  and (_10660_, _04649_, \oc8051_golden_model_1.PSW [7]);
  nor (_10661_, _10660_, _10659_);
  nand (_10662_, _10661_, _03626_);
  and (_10663_, _10662_, _05325_);
  and (_10664_, _10663_, _10658_);
  nand (_10665_, _02578_, _02218_);
  nand (_10666_, _05551_, _10665_);
  or (_10667_, _10666_, _10664_);
  and (_10668_, _10667_, _10614_);
  or (_10669_, _10668_, _02857_);
  or (_10670_, _06173_, _05558_);
  and (_10671_, _10670_, _02853_);
  and (_10672_, _10671_, _10669_);
  and (_10673_, _05311_, _04005_);
  and (_10674_, _05689_, \oc8051_golden_model_1.IP [1]);
  and (_10675_, _05694_, \oc8051_golden_model_1.B [1]);
  nor (_10676_, _10675_, _10674_);
  and (_10677_, _05699_, \oc8051_golden_model_1.PSW [1]);
  and (_10678_, _05703_, \oc8051_golden_model_1.ACC [1]);
  nor (_10679_, _10678_, _10677_);
  and (_10680_, _10679_, _10676_);
  and (_10681_, _05708_, \oc8051_golden_model_1.IE [1]);
  and (_10682_, _05712_, \oc8051_golden_model_1.SBUF [1]);
  and (_10683_, _05714_, \oc8051_golden_model_1.SCON [1]);
  or (_10684_, _10683_, _10682_);
  nor (_10685_, _10684_, _10681_);
  and (_10686_, _05736_, \oc8051_golden_model_1.P0INREG [1]);
  not (_10687_, _10686_);
  and (_10688_, _05733_, \oc8051_golden_model_1.P1INREG [1]);
  not (_10689_, _10688_);
  and (_10690_, _05739_, \oc8051_golden_model_1.P2INREG [1]);
  and (_10691_, _05741_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_10692_, _10691_, _10690_);
  and (_10693_, _10692_, _10689_);
  and (_10694_, _10693_, _10687_);
  and (_10695_, _10694_, _10685_);
  and (_10696_, _10695_, _10680_);
  and (_10697_, _05720_, \oc8051_golden_model_1.TH0 [1]);
  and (_10698_, _05722_, \oc8051_golden_model_1.TL1 [1]);
  nor (_10699_, _10698_, _10697_);
  and (_10700_, _05725_, \oc8051_golden_model_1.TCON [1]);
  and (_10701_, _05729_, \oc8051_golden_model_1.PCON [1]);
  nor (_10702_, _10701_, _10700_);
  and (_10703_, _10702_, _10699_);
  and (_10704_, _05677_, \oc8051_golden_model_1.TL0 [1]);
  and (_10705_, _05681_, \oc8051_golden_model_1.TH1 [1]);
  nor (_10706_, _10705_, _10704_);
  and (_10707_, _05672_, \oc8051_golden_model_1.DPH [1]);
  not (_10708_, _10707_);
  and (_10709_, _10708_, _10706_);
  and (_10710_, _05747_, \oc8051_golden_model_1.SP [1]);
  not (_10711_, _10710_);
  and (_10712_, _05749_, \oc8051_golden_model_1.DPL [1]);
  and (_10713_, _05667_, \oc8051_golden_model_1.TMOD [1]);
  nor (_10714_, _10713_, _10712_);
  and (_10715_, _10714_, _10711_);
  and (_10716_, _10715_, _10709_);
  and (_10717_, _10716_, _10703_);
  and (_10718_, _10717_, _10696_);
  not (_10719_, _10718_);
  nor (_10720_, _10719_, _10673_);
  nor (_10721_, _10720_, _02853_);
  or (_10722_, _10721_, _05562_);
  or (_10723_, _10722_, _10672_);
  and (_10724_, _05562_, _03671_);
  nor (_10726_, _10724_, _03885_);
  and (_10727_, _10726_, _10723_);
  and (_10728_, _03885_, _05675_);
  or (_10729_, _10728_, _02517_);
  or (_10730_, _10729_, _10727_);
  and (_10731_, _02517_, \oc8051_golden_model_1.PC [1]);
  nor (_10732_, _10731_, _05280_);
  and (_10733_, _10732_, _10730_);
  or (_10734_, _10733_, _10613_);
  and (_10735_, _10734_, _05278_);
  nor (_10737_, _05095_, _02618_);
  and (_10738_, _05095_, _02618_);
  nor (_10739_, _10738_, _10737_);
  and (_10740_, _10739_, _05277_);
  or (_10741_, _10740_, _10735_);
  and (_10742_, _10741_, _05276_);
  and (_10743_, _10611_, _05275_);
  or (_10744_, _10743_, _10742_);
  and (_10745_, _10744_, _05273_);
  and (_10746_, _10737_, _03891_);
  or (_10748_, _10746_, _02533_);
  or (_10749_, _10748_, _10745_);
  and (_10750_, _02533_, \oc8051_golden_model_1.PC [1]);
  nor (_10751_, _10750_, _05782_);
  and (_10752_, _10751_, _10749_);
  nor (_10753_, _10610_, _05788_);
  or (_10754_, _10753_, _05787_);
  or (_10755_, _10754_, _10752_);
  nand (_10756_, _10738_, _05787_);
  and (_10757_, _10756_, _05792_);
  and (_10759_, _10757_, _10755_);
  and (_10760_, _02531_, _02218_);
  or (_10761_, _03351_, _10760_);
  or (_10762_, _10761_, _10759_);
  nand (_10763_, _10608_, _03351_);
  and (_10764_, _10763_, _10607_);
  and (_10765_, _10764_, _10762_);
  or (_10766_, _10765_, _10609_);
  and (_10767_, _10766_, _04517_);
  nor (_10768_, _10608_, _04517_);
  or (_10770_, _10768_, _04085_);
  or (_10771_, _10770_, _10767_);
  nand (_10772_, _10608_, _04085_);
  and (_10773_, _10772_, _03910_);
  and (_10774_, _10773_, _10771_);
  or (_10775_, _10774_, _10606_);
  and (_10776_, _10775_, _05801_);
  nor (_10777_, _10622_, _05801_);
  or (_10778_, _10777_, _03004_);
  or (_10779_, _10778_, _10776_);
  nand (_10781_, _03004_, _09082_);
  and (_10782_, _10781_, _02529_);
  and (_10783_, _10782_, _10779_);
  and (_10784_, _02528_, _02218_);
  or (_10785_, _03627_, _10784_);
  or (_10786_, _10785_, _10783_);
  or (_10787_, _10659_, _03936_);
  not (_10788_, _02498_);
  and (_10789_, _03580_, _10788_);
  and (_10790_, _02834_, _02525_);
  nor (_10792_, _10790_, _10789_);
  and (_10793_, _10792_, _10787_);
  and (_10794_, _10793_, _10786_);
  not (_10795_, _10608_);
  nor (_10796_, _10792_, _10795_);
  or (_10797_, _10796_, _06147_);
  or (_10798_, _10797_, _10794_);
  nand (_10799_, _10795_, _06147_);
  and (_10800_, _10799_, _03927_);
  and (_10801_, _10800_, _10798_);
  nor (_10802_, _06175_, _05939_);
  and (_10803_, _10802_, _03926_);
  or (_10804_, _10803_, _03925_);
  or (_10805_, _10804_, _10801_);
  or (_10806_, _10622_, _04176_);
  and (_10807_, _10806_, _04557_);
  and (_10808_, _10807_, _10805_);
  or (_10809_, _10808_, _10419_);
  and (_10810_, _10809_, _10604_);
  nand (_10811_, _09048_, _03004_);
  or (_10812_, _08913_, _03004_);
  and (_10813_, _10812_, _10811_);
  and (_10814_, _10813_, _04551_);
  and (_10815_, _10814_, _10597_);
  or (_32541_, _10815_, _10810_);
  or (_10816_, _10406_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_10817_, _10816_, _10415_);
  or (_10818_, _06161_, _04441_);
  nor (_10819_, _07546_, _06154_);
  and (_10820_, _10819_, _10818_);
  and (_10821_, _05939_, _06029_);
  nor (_10822_, _05939_, _06029_);
  or (_10823_, _10822_, _10821_);
  and (_10824_, _10823_, _03909_);
  and (_10825_, _05261_, _04440_);
  nor (_10826_, _05261_, _04440_);
  or (_10827_, _10826_, _10825_);
  or (_10828_, _10827_, _05270_);
  nor (_10829_, _05142_, _06984_);
  and (_10830_, _05142_, _06984_);
  nor (_10831_, _10830_, _10829_);
  and (_10832_, _10831_, _05277_);
  and (_10833_, _05142_, _03302_);
  nor (_10834_, _05142_, _03302_);
  nor (_10835_, _10834_, _10833_);
  and (_10836_, _10835_, _05280_);
  or (_10837_, _04441_, _05551_);
  nor (_10838_, _09819_, _04653_);
  or (_10839_, _10838_, _05368_);
  or (_10840_, _10827_, _05387_);
  nor (_10841_, _02634_, _02558_);
  and (_10842_, _02558_, \oc8051_golden_model_1.ACC [2]);
  nor (_10843_, _10842_, _10841_);
  nand (_10844_, _10843_, _05387_);
  and (_10845_, _10844_, _10840_);
  and (_10846_, _10845_, _03823_);
  and (_10847_, _05495_, _05142_);
  nor (_10848_, _05495_, _05142_);
  nor (_10849_, _10848_, _10847_);
  nor (_10850_, _10849_, _03823_);
  or (_10851_, _10850_, _10846_);
  and (_10852_, _10851_, _05383_);
  nand (_10853_, _09819_, _09631_);
  and (_10854_, _10853_, _02894_);
  or (_10855_, _10854_, _05382_);
  or (_10856_, _10855_, _10852_);
  nor (_10857_, _02633_, _02556_);
  nor (_10858_, _10857_, _03845_);
  and (_10859_, _10858_, _10856_);
  nor (_10860_, _04440_, _04256_);
  or (_10861_, _10860_, _03853_);
  or (_10862_, _10861_, _10859_);
  and (_10863_, _10862_, _10839_);
  or (_10864_, _10863_, _02886_);
  nand (_10865_, _07670_, _02886_);
  and (_10866_, _10865_, _02884_);
  and (_10867_, _10866_, _10864_);
  not (_10868_, _09820_);
  and (_10869_, _10853_, _10868_);
  and (_10870_, _10869_, _02883_);
  or (_10871_, _10870_, _10867_);
  and (_10872_, _10871_, _02561_);
  or (_10873_, _02634_, _02561_);
  nand (_10874_, _02983_, _10873_);
  or (_10875_, _10874_, _10872_);
  nand (_10876_, _07670_, _02984_);
  and (_10877_, _10876_, _10875_);
  or (_10878_, _10877_, _03867_);
  and (_10879_, _06177_, _02858_);
  nand (_10880_, _07669_, _03867_);
  or (_10881_, _10880_, _10879_);
  and (_10882_, _10881_, _10878_);
  or (_10883_, _10882_, _03626_);
  nor (_10884_, _09654_, _04653_);
  and (_10885_, _04653_, \oc8051_golden_model_1.PSW [7]);
  nor (_10886_, _10885_, _10884_);
  nand (_10887_, _10886_, _03626_);
  and (_10888_, _10887_, _05325_);
  and (_10889_, _10888_, _10883_);
  nand (_10890_, _02633_, _02578_);
  nand (_10891_, _05551_, _10890_);
  or (_10892_, _10891_, _10889_);
  and (_10893_, _10892_, _10837_);
  or (_10894_, _10893_, _02857_);
  or (_10895_, _06177_, _05558_);
  and (_10896_, _10895_, _02853_);
  and (_10897_, _10896_, _10894_);
  nor (_10898_, _05563_, _04440_);
  not (_10899_, _10898_);
  and (_10900_, _05708_, \oc8051_golden_model_1.IE [2]);
  and (_10901_, _05712_, \oc8051_golden_model_1.SBUF [2]);
  and (_10902_, _05714_, \oc8051_golden_model_1.SCON [2]);
  or (_10903_, _10902_, _10901_);
  nor (_10904_, _10903_, _10900_);
  and (_10905_, _05736_, \oc8051_golden_model_1.P0INREG [2]);
  not (_10906_, _10905_);
  and (_10907_, _05733_, \oc8051_golden_model_1.P1INREG [2]);
  not (_10908_, _10907_);
  and (_10909_, _05739_, \oc8051_golden_model_1.P2INREG [2]);
  and (_10910_, _05741_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_10911_, _10910_, _10909_);
  and (_10912_, _10911_, _10908_);
  and (_10913_, _10912_, _10906_);
  and (_10914_, _10913_, _10904_);
  and (_10915_, _05689_, \oc8051_golden_model_1.IP [2]);
  and (_10916_, _05694_, \oc8051_golden_model_1.B [2]);
  nor (_10917_, _10916_, _10915_);
  and (_10918_, _05699_, \oc8051_golden_model_1.PSW [2]);
  and (_10919_, _05703_, \oc8051_golden_model_1.ACC [2]);
  nor (_10920_, _10919_, _10918_);
  and (_10921_, _10920_, _10917_);
  and (_10922_, _05681_, \oc8051_golden_model_1.TH1 [2]);
  and (_10923_, _05672_, \oc8051_golden_model_1.DPH [2]);
  nor (_10924_, _10923_, _10922_);
  and (_10925_, _10924_, _10921_);
  and (_10926_, _10925_, _10914_);
  and (_10927_, _05720_, \oc8051_golden_model_1.TH0 [2]);
  and (_10928_, _05722_, \oc8051_golden_model_1.TL1 [2]);
  nor (_10929_, _10928_, _10927_);
  and (_10930_, _05725_, \oc8051_golden_model_1.TCON [2]);
  and (_10931_, _05729_, \oc8051_golden_model_1.PCON [2]);
  nor (_10932_, _10931_, _10930_);
  and (_10933_, _10932_, _10929_);
  and (_10934_, _05677_, \oc8051_golden_model_1.TL0 [2]);
  and (_10935_, _05667_, \oc8051_golden_model_1.TMOD [2]);
  nor (_10936_, _10935_, _10934_);
  and (_10937_, _05747_, \oc8051_golden_model_1.SP [2]);
  and (_10938_, _05749_, \oc8051_golden_model_1.DPL [2]);
  nor (_10939_, _10938_, _10937_);
  and (_10940_, _10939_, _10936_);
  and (_10941_, _10940_, _10933_);
  and (_10942_, _10941_, _10926_);
  and (_10943_, _10942_, _10899_);
  nor (_10944_, _10943_, _02853_);
  or (_10945_, _10944_, _05562_);
  or (_10946_, _10945_, _10897_);
  and (_10947_, _05562_, _03260_);
  nor (_10948_, _10947_, _03885_);
  and (_10949_, _10948_, _10946_);
  and (_10950_, _03885_, _05727_);
  or (_10951_, _10950_, _02517_);
  or (_10952_, _10951_, _10949_);
  and (_10953_, _02634_, _02517_);
  nor (_10954_, _10953_, _05280_);
  and (_10955_, _10954_, _10952_);
  or (_10956_, _10955_, _10836_);
  and (_10957_, _10956_, _05278_);
  or (_10958_, _10957_, _10832_);
  and (_10959_, _10958_, _05276_);
  and (_10960_, _10834_, _05275_);
  or (_10961_, _10960_, _10959_);
  and (_10962_, _10961_, _05273_);
  and (_10963_, _10829_, _03891_);
  or (_10964_, _10963_, _02533_);
  or (_10965_, _10964_, _10962_);
  and (_10966_, _02634_, _02533_);
  nor (_10967_, _10966_, _05782_);
  and (_10968_, _10967_, _10965_);
  nor (_10969_, _10833_, _05788_);
  or (_10970_, _10969_, _05787_);
  or (_10971_, _10970_, _10968_);
  nand (_10972_, _10830_, _05787_);
  and (_10973_, _10972_, _05792_);
  and (_10974_, _10973_, _10971_);
  or (_10975_, _03711_, _03566_);
  and (_10976_, _02633_, _02531_);
  and (_10977_, _05269_, _10788_);
  or (_10978_, _10977_, _10976_);
  or (_10979_, _10978_, _10975_);
  or (_10980_, _10979_, _10974_);
  and (_10981_, _10980_, _10828_);
  or (_10982_, _10981_, _04085_);
  or (_10983_, _10827_, _04084_);
  and (_10984_, _10983_, _03910_);
  and (_10985_, _10984_, _10982_);
  or (_10986_, _10985_, _10824_);
  and (_10987_, _10986_, _05801_);
  nor (_10988_, _10849_, _05801_);
  or (_10989_, _10988_, _03004_);
  or (_10990_, _10989_, _10987_);
  nand (_10991_, _09080_, _03004_);
  and (_10992_, _10991_, _02529_);
  and (_10993_, _10992_, _10990_);
  and (_10994_, _02633_, _02528_);
  or (_10995_, _03627_, _10994_);
  or (_10996_, _10995_, _10993_);
  or (_10997_, _10884_, _03936_);
  and (_10998_, _10997_, _06154_);
  and (_10999_, _10998_, _10996_);
  or (_11000_, _10999_, _10820_);
  and (_11001_, _11000_, _03927_);
  or (_11002_, _06175_, _06177_);
  nor (_11003_, _07376_, _03927_);
  and (_11004_, _11003_, _11002_);
  or (_11005_, _11004_, _03925_);
  or (_11006_, _11005_, _11001_);
  nor (_11007_, _05143_, _05096_);
  nor (_11008_, _11007_, _05144_);
  or (_11009_, _11008_, _04176_);
  and (_11010_, _11009_, _04557_);
  and (_11011_, _11010_, _11006_);
  or (_11012_, _11011_, _10419_);
  and (_11013_, _11012_, _10817_);
  nand (_11014_, _09040_, _03004_);
  or (_11015_, _08908_, _03004_);
  and (_11016_, _11015_, _11014_);
  and (_11017_, _11016_, _04551_);
  and (_11018_, _11017_, _10597_);
  or (_32543_, _11018_, _11013_);
  or (_11019_, _10406_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_11020_, _11019_, _10415_);
  not (_11021_, _10406_);
  nor (_11022_, _10821_, _05984_);
  or (_11023_, _11022_, _06031_);
  and (_11024_, _11023_, _03909_);
  and (_11025_, _02676_, _02531_);
  nor (_11026_, _04995_, _02701_);
  and (_11027_, _04995_, _02701_);
  nor (_11028_, _11027_, _11026_);
  and (_11029_, _11028_, _05277_);
  and (_11030_, _04995_, _03120_);
  nor (_11031_, _04995_, _03120_);
  nor (_11032_, _11031_, _11030_);
  and (_11033_, _11032_, _05280_);
  nand (_11034_, _07651_, _02984_);
  nor (_11035_, _09879_, _04631_);
  or (_11036_, _11035_, _05368_);
  nand (_11037_, _09879_, _09551_);
  or (_11038_, _11037_, _05383_);
  nor (_11039_, _10847_, _04995_);
  nor (_11040_, _11039_, _05497_);
  nor (_11041_, _11040_, _03823_);
  nor (_11042_, _10825_, _04242_);
  or (_11043_, _11042_, _05263_);
  or (_11044_, _11043_, _05387_);
  nor (_11045_, _02677_, _02558_);
  and (_11046_, _02558_, \oc8051_golden_model_1.ACC [3]);
  nor (_11047_, _11046_, _11045_);
  and (_11048_, _11047_, _05387_);
  nor (_11049_, _11048_, _03822_);
  and (_11050_, _11049_, _11044_);
  or (_11051_, _11050_, _02894_);
  or (_11052_, _11051_, _11041_);
  and (_11053_, _11052_, _11038_);
  or (_11054_, _11053_, _05382_);
  nor (_11055_, _02676_, _02556_);
  nor (_11056_, _11055_, _03845_);
  and (_11057_, _11056_, _11054_);
  nor (_11058_, _04242_, _04256_);
  or (_11059_, _11058_, _03853_);
  or (_11060_, _11059_, _11057_);
  and (_11061_, _11060_, _11036_);
  or (_11062_, _11061_, _02886_);
  nand (_11063_, _07651_, _02886_);
  and (_11064_, _11063_, _02884_);
  and (_11065_, _11064_, _11062_);
  not (_11066_, _09880_);
  and (_11067_, _11037_, _11066_);
  and (_11068_, _11067_, _02883_);
  or (_11069_, _11068_, _11065_);
  and (_11070_, _11069_, _02561_);
  or (_11071_, _02677_, _02561_);
  nand (_11072_, _02983_, _11071_);
  or (_11073_, _11072_, _11070_);
  and (_11074_, _11073_, _11034_);
  or (_11075_, _11074_, _03867_);
  and (_11076_, _06176_, _02858_);
  nand (_11077_, _07650_, _03867_);
  or (_11078_, _11077_, _11076_);
  and (_11079_, _11078_, _11075_);
  or (_11080_, _11079_, _03626_);
  and (_11081_, _04631_, \oc8051_golden_model_1.PSW [7]);
  nor (_11082_, _09574_, _04631_);
  nor (_11083_, _11082_, _11081_);
  nand (_11084_, _11083_, _03626_);
  and (_11085_, _11084_, _05325_);
  and (_11086_, _11085_, _11080_);
  nand (_11087_, _02676_, _02578_);
  nand (_11088_, _05551_, _11087_);
  or (_11089_, _11088_, _11086_);
  or (_11090_, _05412_, _05551_);
  and (_11091_, _11090_, _11089_);
  or (_11092_, _11091_, _02857_);
  or (_11093_, _06176_, _05558_);
  and (_11094_, _11093_, _02853_);
  and (_11095_, _11094_, _11092_);
  nor (_11096_, _05563_, _04242_);
  not (_11097_, _11096_);
  and (_11098_, _05689_, \oc8051_golden_model_1.IP [3]);
  and (_11099_, _05694_, \oc8051_golden_model_1.B [3]);
  nor (_11100_, _11099_, _11098_);
  and (_11101_, _05699_, \oc8051_golden_model_1.PSW [3]);
  and (_11102_, _05703_, \oc8051_golden_model_1.ACC [3]);
  nor (_11103_, _11102_, _11101_);
  and (_11104_, _11103_, _11100_);
  and (_11105_, _05708_, \oc8051_golden_model_1.IE [3]);
  and (_11106_, _05712_, \oc8051_golden_model_1.SBUF [3]);
  and (_11107_, _05714_, \oc8051_golden_model_1.SCON [3]);
  or (_11108_, _11107_, _11106_);
  nor (_11109_, _11108_, _11105_);
  and (_11110_, _05736_, \oc8051_golden_model_1.P0INREG [3]);
  not (_11111_, _11110_);
  and (_11112_, _05733_, \oc8051_golden_model_1.P1INREG [3]);
  not (_11113_, _11112_);
  and (_11114_, _05739_, \oc8051_golden_model_1.P2INREG [3]);
  and (_11115_, _05741_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_11116_, _11115_, _11114_);
  and (_11117_, _11116_, _11113_);
  and (_11118_, _11117_, _11111_);
  and (_11119_, _11118_, _11109_);
  and (_11120_, _11119_, _11104_);
  and (_11121_, _05720_, \oc8051_golden_model_1.TH0 [3]);
  and (_11122_, _05722_, \oc8051_golden_model_1.TL1 [3]);
  nor (_11123_, _11122_, _11121_);
  and (_11124_, _05725_, \oc8051_golden_model_1.TCON [3]);
  and (_11125_, _05729_, \oc8051_golden_model_1.PCON [3]);
  nor (_11126_, _11125_, _11124_);
  and (_11127_, _11126_, _11123_);
  and (_11128_, _05677_, \oc8051_golden_model_1.TL0 [3]);
  and (_11129_, _05681_, \oc8051_golden_model_1.TH1 [3]);
  nor (_11130_, _11129_, _11128_);
  and (_11131_, _05672_, \oc8051_golden_model_1.DPH [3]);
  not (_11132_, _11131_);
  and (_11133_, _11132_, _11130_);
  and (_11134_, _05747_, \oc8051_golden_model_1.SP [3]);
  not (_11135_, _11134_);
  and (_11136_, _05749_, \oc8051_golden_model_1.DPL [3]);
  and (_11137_, _05667_, \oc8051_golden_model_1.TMOD [3]);
  nor (_11138_, _11137_, _11136_);
  and (_11139_, _11138_, _11135_);
  and (_11140_, _11139_, _11133_);
  and (_11141_, _11140_, _11127_);
  and (_11142_, _11141_, _11120_);
  and (_11143_, _11142_, _11097_);
  nor (_11144_, _11143_, _02853_);
  or (_11145_, _11144_, _05562_);
  or (_11146_, _11145_, _11095_);
  and (_11147_, _05562_, _02799_);
  nor (_11148_, _11147_, _03885_);
  and (_11149_, _11148_, _11146_);
  and (_11150_, _03885_, _05664_);
  or (_11151_, _11150_, _02517_);
  or (_11152_, _11151_, _11149_);
  and (_11153_, _02677_, _02517_);
  nor (_11154_, _11153_, _05280_);
  and (_11155_, _11154_, _11152_);
  or (_11156_, _11155_, _11033_);
  and (_11157_, _11156_, _05278_);
  or (_11158_, _11157_, _11029_);
  and (_11159_, _11158_, _05276_);
  and (_11160_, _11031_, _05275_);
  or (_11161_, _11160_, _11159_);
  and (_11162_, _11161_, _05273_);
  and (_11163_, _11026_, _03891_);
  or (_11164_, _11163_, _02533_);
  or (_11165_, _11164_, _11162_);
  and (_11166_, _02677_, _02533_);
  nor (_11167_, _11166_, _05782_);
  and (_11168_, _11167_, _11165_);
  nor (_11169_, _11030_, _05788_);
  or (_11170_, _11169_, _05787_);
  or (_11171_, _11170_, _11168_);
  nand (_11172_, _11027_, _05787_);
  and (_11173_, _11172_, _05792_);
  and (_11174_, _11173_, _11171_);
  or (_11175_, _11174_, _11025_);
  and (_11176_, _11175_, _05270_);
  not (_11177_, _05270_);
  and (_11178_, _11043_, _11177_);
  or (_11179_, _11178_, _04085_);
  or (_11180_, _11179_, _11176_);
  or (_11181_, _11043_, _04084_);
  and (_11182_, _11181_, _03910_);
  and (_11183_, _11182_, _11180_);
  or (_11184_, _11183_, _11024_);
  and (_11185_, _11184_, _05801_);
  nor (_11186_, _11040_, _05801_);
  or (_11187_, _11186_, _03004_);
  or (_11188_, _11187_, _11185_);
  nand (_11189_, _09075_, _03004_);
  and (_11190_, _11189_, _02529_);
  and (_11191_, _11190_, _11188_);
  and (_11192_, _02676_, _02528_);
  or (_11193_, _03627_, _11192_);
  or (_11194_, _11193_, _11191_);
  or (_11195_, _11082_, _03936_);
  and (_11196_, _11195_, _06153_);
  and (_11197_, _11196_, _11194_);
  not (_11198_, _06149_);
  nor (_11199_, _07546_, _05412_);
  nor (_11200_, _11199_, _06163_);
  or (_11201_, _11200_, _11198_);
  and (_11202_, _11201_, _06155_);
  or (_11203_, _11202_, _11197_);
  or (_11204_, _11200_, _06149_);
  and (_11205_, _11204_, _03927_);
  and (_11206_, _11205_, _11203_);
  or (_11207_, _07376_, _06176_);
  nor (_11208_, _06179_, _03927_);
  and (_11209_, _11208_, _11207_);
  or (_11210_, _11209_, _03925_);
  or (_11211_, _11210_, _11206_);
  nor (_11212_, _05144_, _04996_);
  nor (_11213_, _11212_, _05145_);
  or (_11214_, _11213_, _04176_);
  and (_11215_, _11214_, _04186_);
  and (_11216_, _11215_, _11211_);
  or (_11217_, _11216_, _11021_);
  and (_11218_, _11217_, _11020_);
  nand (_11219_, _09033_, _03004_);
  or (_11220_, _08904_, _03004_);
  and (_11221_, _11220_, _11219_);
  and (_11222_, _11221_, _04551_);
  and (_11223_, _11222_, _10597_);
  or (_32544_, _11223_, _11218_);
  or (_11224_, _10406_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_11225_, _11224_, _10415_);
  nor (_11226_, _06179_, _06181_);
  nor (_11227_, _11226_, _07353_);
  or (_11228_, _11227_, _03927_);
  and (_11229_, _06031_, _06121_);
  nor (_11230_, _06031_, _06121_);
  or (_11231_, _11230_, _11229_);
  and (_11232_, _11231_, _03909_);
  nor (_11233_, _05263_, _05202_);
  and (_11234_, _05263_, _05202_);
  or (_11235_, _11234_, _11233_);
  or (_11236_, _11235_, _05270_);
  nor (_11237_, _05630_, _05250_);
  and (_11238_, _11237_, _05275_);
  nor (_11239_, _09705_, _09682_);
  and (_11240_, _09682_, \oc8051_golden_model_1.PSW [7]);
  nor (_11241_, _11240_, _11239_);
  nor (_11242_, _11241_, _04303_);
  nor (_11243_, _09682_, _09843_);
  or (_11244_, _11243_, _05368_);
  nand (_11245_, _09683_, _09843_);
  or (_11246_, _11245_, _05383_);
  or (_11247_, _11235_, _05387_);
  and (_11248_, _02558_, \oc8051_golden_model_1.ACC [4]);
  nor (_11249_, _08937_, _02558_);
  nor (_11250_, _11249_, _11248_);
  nand (_11251_, _11250_, _05387_);
  and (_11252_, _11251_, _11247_);
  or (_11253_, _11252_, _03818_);
  or (_11254_, _06181_, _05402_);
  and (_11255_, _11254_, _11253_);
  or (_11256_, _11255_, _03822_);
  and (_11257_, _05497_, _05250_);
  nor (_11258_, _05497_, _05250_);
  nor (_11259_, _11258_, _11257_);
  nand (_11260_, _11259_, _03822_);
  and (_11261_, _11260_, _11256_);
  or (_11262_, _11261_, _02894_);
  and (_11263_, _11262_, _11246_);
  or (_11264_, _11263_, _05382_);
  nor (_11265_, _08936_, _02556_);
  nor (_11266_, _11265_, _03845_);
  and (_11267_, _11266_, _11264_);
  nor (_11268_, _05202_, _04256_);
  or (_11269_, _11268_, _03853_);
  or (_11270_, _11269_, _11267_);
  and (_11271_, _11270_, _11244_);
  or (_11272_, _11271_, _02886_);
  nand (_11273_, _07640_, _02886_);
  and (_11274_, _11273_, _02884_);
  and (_11275_, _11274_, _11272_);
  not (_11276_, _09844_);
  and (_11277_, _11245_, _11276_);
  and (_11278_, _11277_, _02883_);
  or (_11279_, _11278_, _11275_);
  and (_11280_, _11279_, _02561_);
  or (_11281_, _08937_, _02561_);
  nand (_11282_, _11281_, _02983_);
  or (_11283_, _11282_, _11280_);
  nand (_11284_, _07640_, _02984_);
  and (_11285_, _11284_, _11283_);
  or (_11286_, _11285_, _03867_);
  and (_11287_, _06181_, _02858_);
  nand (_11288_, _07639_, _03867_);
  or (_11289_, _11288_, _11287_);
  and (_11290_, _11289_, _04303_);
  and (_11291_, _11290_, _11286_);
  or (_11292_, _11291_, _11242_);
  and (_11293_, _11292_, _05325_);
  nand (_11294_, _08936_, _02578_);
  nand (_11295_, _11294_, _05551_);
  or (_11296_, _11295_, _11293_);
  or (_11297_, _06160_, _05551_);
  and (_11298_, _11297_, _11296_);
  or (_11299_, _11298_, _02857_);
  or (_11300_, _06181_, _05558_);
  and (_11301_, _11300_, _02853_);
  and (_11302_, _11301_, _11299_);
  nor (_11303_, _05563_, _05202_);
  not (_11304_, _11303_);
  and (_11305_, _05749_, \oc8051_golden_model_1.DPL [4]);
  and (_11306_, _05677_, \oc8051_golden_model_1.TL0 [4]);
  nor (_11307_, _11306_, _11305_);
  and (_11308_, _05681_, \oc8051_golden_model_1.TH1 [4]);
  and (_11309_, _05672_, \oc8051_golden_model_1.DPH [4]);
  nor (_11310_, _11309_, _11308_);
  and (_11311_, _11310_, _11307_);
  and (_11312_, _05689_, \oc8051_golden_model_1.IP [4]);
  and (_11313_, _05694_, \oc8051_golden_model_1.B [4]);
  nor (_11314_, _11313_, _11312_);
  and (_11315_, _05699_, \oc8051_golden_model_1.PSW [4]);
  and (_11316_, _05703_, \oc8051_golden_model_1.ACC [4]);
  nor (_11317_, _11316_, _11315_);
  and (_11318_, _11317_, _11314_);
  and (_11319_, _05708_, \oc8051_golden_model_1.IE [4]);
  and (_11320_, _05712_, \oc8051_golden_model_1.SBUF [4]);
  and (_11321_, _05714_, \oc8051_golden_model_1.SCON [4]);
  or (_11322_, _11321_, _11320_);
  nor (_11323_, _11322_, _11319_);
  and (_11324_, _11323_, _11318_);
  and (_11325_, _11324_, _11311_);
  and (_11326_, _05720_, \oc8051_golden_model_1.TH0 [4]);
  and (_11327_, _05722_, \oc8051_golden_model_1.TL1 [4]);
  nor (_11328_, _11327_, _11326_);
  and (_11329_, _05725_, \oc8051_golden_model_1.TCON [4]);
  and (_11330_, _05729_, \oc8051_golden_model_1.PCON [4]);
  nor (_11331_, _11330_, _11329_);
  and (_11332_, _11331_, _11328_);
  and (_11333_, _05733_, \oc8051_golden_model_1.P1INREG [4]);
  not (_11334_, _11333_);
  and (_11335_, _05736_, \oc8051_golden_model_1.P0INREG [4]);
  not (_11336_, _11335_);
  and (_11337_, _05739_, \oc8051_golden_model_1.P2INREG [4]);
  and (_11338_, _05741_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_11339_, _11338_, _11337_);
  and (_11340_, _11339_, _11336_);
  and (_11341_, _11340_, _11334_);
  and (_11342_, _05747_, \oc8051_golden_model_1.SP [4]);
  and (_11343_, _05667_, \oc8051_golden_model_1.TMOD [4]);
  nor (_11344_, _11343_, _11342_);
  and (_11345_, _11344_, _11341_);
  and (_11346_, _11345_, _11332_);
  and (_11347_, _11346_, _11325_);
  and (_11348_, _11347_, _11304_);
  nor (_11349_, _11348_, _02853_);
  or (_11350_, _11349_, _05562_);
  or (_11351_, _11350_, _11302_);
  and (_11352_, _05562_, _03625_);
  nor (_11353_, _11352_, _03885_);
  and (_11354_, _11353_, _11351_);
  and (_11355_, _05697_, _03885_);
  or (_11356_, _11355_, _02517_);
  or (_11357_, _11356_, _11354_);
  and (_11358_, _08937_, _02517_);
  nor (_11359_, _11358_, _05280_);
  and (_11360_, _11359_, _11357_);
  and (_11361_, _05630_, _05250_);
  nor (_11362_, _11361_, _11237_);
  and (_11363_, _11362_, _05280_);
  or (_11364_, _11363_, _05277_);
  or (_11365_, _11364_, _11360_);
  nor (_11366_, _05250_, _06885_);
  and (_11367_, _05250_, _06885_);
  nor (_11368_, _11367_, _11366_);
  or (_11369_, _11368_, _05278_);
  and (_11370_, _11369_, _05276_);
  and (_11371_, _11370_, _11365_);
  or (_11372_, _11371_, _11238_);
  and (_11373_, _11372_, _05273_);
  and (_11374_, _11366_, _03891_);
  or (_11375_, _11374_, _02533_);
  or (_11376_, _11375_, _11373_);
  and (_11377_, _08937_, _02533_);
  nor (_11378_, _11377_, _05782_);
  and (_11379_, _11378_, _11376_);
  nor (_11380_, _11361_, _05788_);
  or (_11381_, _11380_, _05787_);
  or (_11382_, _11381_, _11379_);
  nand (_11383_, _11367_, _05787_);
  and (_11384_, _11383_, _05792_);
  and (_11385_, _11384_, _11382_);
  and (_11386_, _08936_, _02531_);
  or (_11387_, _11386_, _10977_);
  or (_11388_, _11387_, _10975_);
  or (_11389_, _11388_, _11385_);
  and (_11390_, _11389_, _11236_);
  or (_11391_, _11390_, _04085_);
  or (_11392_, _11235_, _04084_);
  and (_11393_, _11392_, _03910_);
  and (_11394_, _11393_, _11391_);
  or (_11395_, _11394_, _11232_);
  and (_11396_, _11395_, _05801_);
  nor (_11397_, _11259_, _05801_);
  or (_11398_, _11397_, _03004_);
  or (_11399_, _11398_, _11396_);
  nand (_11400_, _09070_, _03004_);
  and (_11401_, _11400_, _02529_);
  and (_11402_, _11401_, _11399_);
  and (_11403_, _08936_, _02528_);
  or (_11404_, _11403_, _03627_);
  or (_11405_, _11404_, _11402_);
  or (_11406_, _11239_, _03936_);
  and (_11407_, _11406_, _06154_);
  and (_11408_, _11407_, _11405_);
  or (_11409_, _06163_, _06160_);
  nor (_11410_, _06164_, _06154_);
  and (_11411_, _11410_, _11409_);
  or (_11412_, _11411_, _03926_);
  or (_11413_, _11412_, _11408_);
  and (_11414_, _11413_, _11228_);
  or (_11415_, _11414_, _03925_);
  nor (_11416_, _05251_, _05145_);
  nor (_11417_, _11416_, _05252_);
  or (_11418_, _11417_, _04176_);
  and (_11419_, _11418_, _04557_);
  and (_11420_, _11419_, _11415_);
  or (_11421_, _11420_, _10419_);
  and (_11422_, _11421_, _11225_);
  not (_11423_, _08899_);
  nor (_11424_, _11423_, _03004_);
  and (_11425_, _09027_, _03004_);
  or (_11426_, _11425_, _11424_);
  and (_11427_, _11426_, _04551_);
  and (_11428_, _11427_, _10597_);
  or (_32545_, _11428_, _11422_);
  or (_11429_, _10406_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_11430_, _11429_, _10415_);
  nor (_11431_, _11234_, _04896_);
  or (_11432_, _11431_, _05264_);
  or (_11433_, _11432_, _05271_);
  nor (_11434_, _04943_, _06879_);
  and (_11435_, _04943_, _06879_);
  nor (_11436_, _11435_, _11434_);
  and (_11437_, _11436_, _05277_);
  nor (_11438_, _09601_, _09577_);
  and (_11439_, _09577_, \oc8051_golden_model_1.PSW [7]);
  nor (_11440_, _11439_, _11438_);
  nor (_11441_, _11440_, _04303_);
  nor (_11442_, _09577_, _09892_);
  or (_11443_, _11442_, _05368_);
  nor (_11444_, _11257_, _04943_);
  nor (_11445_, _11444_, _05498_);
  nor (_11446_, _11445_, _03823_);
  or (_11447_, _06180_, _05402_);
  and (_11448_, _11432_, _10433_);
  or (_11449_, _08931_, _02558_);
  nand (_11450_, _02558_, _06879_);
  and (_11451_, _11450_, _11449_);
  and (_11452_, _11451_, _05387_);
  or (_11453_, _11452_, _03818_);
  or (_11454_, _11453_, _11448_);
  and (_11455_, _11454_, _03823_);
  and (_11456_, _11455_, _11447_);
  or (_11457_, _11456_, _11446_);
  and (_11458_, _11457_, _05383_);
  nand (_11459_, _09578_, _09892_);
  and (_11460_, _11459_, _02894_);
  or (_11461_, _11460_, _05382_);
  or (_11462_, _11461_, _11458_);
  nor (_11463_, _08931_, _02556_);
  nor (_11464_, _11463_, _03845_);
  and (_11465_, _11464_, _11462_);
  nor (_11466_, _04896_, _04256_);
  or (_11467_, _11466_, _03853_);
  or (_11468_, _11467_, _11465_);
  and (_11469_, _11468_, _11443_);
  or (_11470_, _11469_, _02886_);
  nand (_11471_, _07624_, _02886_);
  and (_11472_, _11471_, _02884_);
  and (_11473_, _11472_, _11470_);
  not (_11474_, _09893_);
  and (_11475_, _11459_, _11474_);
  and (_11476_, _11475_, _02883_);
  or (_11477_, _11476_, _11473_);
  and (_11478_, _11477_, _02561_);
  or (_11479_, _08932_, _02561_);
  nand (_11480_, _11479_, _02983_);
  or (_11481_, _11480_, _11478_);
  nand (_11482_, _07624_, _02984_);
  and (_11483_, _11482_, _11481_);
  or (_11484_, _11483_, _03867_);
  and (_11485_, _06180_, _02858_);
  nand (_11486_, _07623_, _03867_);
  or (_11487_, _11486_, _11485_);
  and (_11488_, _11487_, _04303_);
  and (_11489_, _11488_, _11484_);
  or (_11490_, _11489_, _11441_);
  and (_11491_, _11490_, _05325_);
  nand (_11492_, _08931_, _02578_);
  nand (_11493_, _11492_, _05551_);
  or (_11494_, _11493_, _11491_);
  or (_11495_, _06159_, _05551_);
  and (_11496_, _11495_, _11494_);
  or (_11497_, _11496_, _02857_);
  or (_11498_, _06180_, _05558_);
  and (_11499_, _11498_, _02853_);
  and (_11500_, _11499_, _11497_);
  nor (_11501_, _05563_, _04896_);
  not (_11502_, _11501_);
  and (_11503_, _05667_, \oc8051_golden_model_1.TMOD [5]);
  and (_11504_, _05672_, \oc8051_golden_model_1.DPH [5]);
  nor (_11505_, _11504_, _11503_);
  and (_11506_, _05677_, \oc8051_golden_model_1.TL0 [5]);
  and (_11507_, _05681_, \oc8051_golden_model_1.TH1 [5]);
  nor (_11508_, _11507_, _11506_);
  and (_11509_, _11508_, _11505_);
  and (_11510_, _05689_, \oc8051_golden_model_1.IP [5]);
  and (_11511_, _05694_, \oc8051_golden_model_1.B [5]);
  nor (_11512_, _11511_, _11510_);
  and (_11513_, _05699_, \oc8051_golden_model_1.PSW [5]);
  and (_11514_, _05703_, \oc8051_golden_model_1.ACC [5]);
  nor (_11515_, _11514_, _11513_);
  and (_11516_, _11515_, _11512_);
  and (_11517_, _05708_, \oc8051_golden_model_1.IE [5]);
  and (_11518_, _05712_, \oc8051_golden_model_1.SBUF [5]);
  and (_11519_, _05714_, \oc8051_golden_model_1.SCON [5]);
  or (_11520_, _11519_, _11518_);
  nor (_11521_, _11520_, _11517_);
  and (_11522_, _11521_, _11516_);
  and (_11523_, _11522_, _11509_);
  and (_11524_, _05720_, \oc8051_golden_model_1.TH0 [5]);
  and (_11525_, _05722_, \oc8051_golden_model_1.TL1 [5]);
  nor (_11526_, _11525_, _11524_);
  and (_11527_, _05725_, \oc8051_golden_model_1.TCON [5]);
  and (_11528_, _05729_, \oc8051_golden_model_1.PCON [5]);
  nor (_11529_, _11528_, _11527_);
  and (_11530_, _11529_, _11526_);
  and (_11531_, _05733_, \oc8051_golden_model_1.P1INREG [5]);
  not (_11532_, _11531_);
  and (_11533_, _05736_, \oc8051_golden_model_1.P0INREG [5]);
  not (_11534_, _11533_);
  and (_11535_, _05739_, \oc8051_golden_model_1.P2INREG [5]);
  and (_11536_, _05741_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_11537_, _11536_, _11535_);
  and (_11538_, _11537_, _11534_);
  and (_11539_, _11538_, _11532_);
  and (_11540_, _05747_, \oc8051_golden_model_1.SP [5]);
  and (_11541_, _05749_, \oc8051_golden_model_1.DPL [5]);
  nor (_11542_, _11541_, _11540_);
  and (_11543_, _11542_, _11539_);
  and (_11544_, _11543_, _11530_);
  and (_11545_, _11544_, _11523_);
  and (_11546_, _11545_, _11502_);
  nor (_11547_, _11546_, _02853_);
  or (_11548_, _11547_, _05562_);
  or (_11549_, _11548_, _11500_);
  and (_11550_, _05562_, _03215_);
  nor (_11551_, _11550_, _03885_);
  and (_11552_, _11551_, _11549_);
  and (_11553_, _05701_, _03885_);
  or (_11554_, _11553_, _02517_);
  or (_11555_, _11554_, _11552_);
  nand (_11556_, _08932_, _02517_);
  and (_11557_, _11556_, _11555_);
  or (_11558_, _11557_, _05280_);
  not (_11559_, _05280_);
  and (_11560_, _05661_, _04943_);
  nor (_11561_, _05661_, _04943_);
  nor (_11562_, _11561_, _11560_);
  or (_11563_, _11562_, _11559_);
  and (_11564_, _11563_, _05278_);
  and (_11565_, _11564_, _11558_);
  or (_11566_, _11565_, _11437_);
  and (_11567_, _11566_, _05276_);
  and (_11568_, _11561_, _05275_);
  or (_11569_, _11568_, _11567_);
  and (_11570_, _11569_, _05273_);
  and (_11571_, _11434_, _03891_);
  or (_11572_, _11571_, _02533_);
  or (_11573_, _11572_, _11570_);
  and (_11574_, _08932_, _02533_);
  nor (_11575_, _11574_, _05782_);
  and (_11576_, _11575_, _11573_);
  nor (_11577_, _11560_, _05788_);
  or (_11578_, _11577_, _05787_);
  or (_11579_, _11578_, _11576_);
  nand (_11580_, _11435_, _05787_);
  and (_11581_, _11580_, _05792_);
  and (_11582_, _11581_, _11579_);
  nand (_11583_, _08931_, _02531_);
  nor (_11584_, _11177_, _04083_);
  nand (_11585_, _11584_, _11583_);
  or (_11586_, _11585_, _11582_);
  and (_11587_, _11586_, _11433_);
  and (_11588_, _11432_, _03570_);
  or (_11589_, _11588_, _03909_);
  or (_11590_, _11589_, _11587_);
  nor (_11591_, _11229_, _06076_);
  or (_11592_, _06123_, _03910_);
  or (_11593_, _11592_, _11591_);
  and (_11594_, _11593_, _05801_);
  and (_11595_, _11594_, _11590_);
  nor (_11596_, _11445_, _05801_);
  or (_11597_, _11596_, _03004_);
  or (_11598_, _11597_, _11595_);
  nand (_11599_, _09065_, _03004_);
  and (_11600_, _11599_, _02529_);
  and (_11601_, _11600_, _11598_);
  and (_11602_, _08931_, _02528_);
  or (_11603_, _11602_, _03627_);
  or (_11604_, _11603_, _11601_);
  or (_11605_, _11438_, _03936_);
  and (_11606_, _11605_, _06154_);
  and (_11607_, _11606_, _11604_);
  or (_11608_, _06164_, _06159_);
  nor (_11609_, _06165_, _06154_);
  and (_11610_, _11609_, _11608_);
  or (_11611_, _11610_, _11607_);
  and (_11612_, _11611_, _03927_);
  or (_11613_, _07353_, _06180_);
  nor (_11614_, _06183_, _03927_);
  and (_11615_, _11614_, _11613_);
  or (_11616_, _11615_, _03925_);
  or (_11617_, _11616_, _11612_);
  nor (_11618_, _05252_, _04944_);
  nor (_11619_, _11618_, _05253_);
  or (_11620_, _11619_, _04176_);
  and (_11621_, _11620_, _04186_);
  and (_11622_, _11621_, _11617_);
  or (_11623_, _11622_, _11021_);
  and (_11624_, _11623_, _11430_);
  nand (_11625_, _09023_, _03004_);
  or (_11626_, _08894_, _03004_);
  and (_11627_, _11626_, _11625_);
  and (_11628_, _11627_, _04551_);
  and (_11629_, _11628_, _10597_);
  or (_32546_, _11629_, _11624_);
  or (_11630_, _10406_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_11631_, _11630_, _10415_);
  nor (_11632_, _06183_, _05847_);
  nor (_11633_, _11632_, _06184_);
  or (_11634_, _11633_, _03927_);
  nor (_11635_, _05498_, _04837_);
  nor (_11636_, _11635_, _05499_);
  nor (_11637_, _11636_, _05801_);
  nor (_11638_, _06123_, _05848_);
  or (_11639_, _11638_, _06124_);
  and (_11640_, _11639_, _03909_);
  nor (_11641_, _05264_, _04787_);
  or (_11642_, _11641_, _05265_);
  or (_11643_, _11642_, _05270_);
  and (_11644_, _05598_, _04837_);
  nor (_11645_, _05598_, _04837_);
  nor (_11646_, _11645_, _11644_);
  and (_11647_, _11646_, _05280_);
  nor (_11648_, _09549_, _09525_);
  and (_11649_, _09525_, \oc8051_golden_model_1.PSW [7]);
  nor (_11650_, _11649_, _11648_);
  nor (_11651_, _11650_, _04303_);
  nor (_11652_, _04787_, _04256_);
  nand (_11653_, _09526_, _09868_);
  or (_11654_, _11653_, _05383_);
  or (_11655_, _05847_, _05402_);
  and (_11656_, _11642_, _10433_);
  and (_11657_, _02558_, \oc8051_golden_model_1.ACC [6]);
  nor (_11658_, _08924_, _02558_);
  or (_11659_, _11658_, _11657_);
  and (_11660_, _11659_, _05387_);
  or (_11661_, _11660_, _03818_);
  or (_11662_, _11661_, _11656_);
  and (_11663_, _11662_, _11655_);
  or (_11664_, _11663_, _03822_);
  nand (_11665_, _11636_, _03822_);
  and (_11666_, _11665_, _11664_);
  or (_11667_, _11666_, _02894_);
  and (_11668_, _11667_, _11654_);
  or (_11669_, _11668_, _05382_);
  nor (_11670_, _08923_, _02556_);
  nor (_11671_, _11670_, _03845_);
  and (_11672_, _11671_, _11669_);
  or (_11673_, _11672_, _11652_);
  and (_11674_, _11673_, _05368_);
  nor (_11675_, _09525_, _09868_);
  and (_11676_, _11675_, _03853_);
  or (_11677_, _11676_, _02886_);
  or (_11678_, _11677_, _11674_);
  nand (_11679_, _07610_, _02886_);
  and (_11680_, _11679_, _02884_);
  and (_11681_, _11680_, _11678_);
  not (_11682_, _09869_);
  and (_11683_, _11653_, _11682_);
  and (_11684_, _11683_, _02883_);
  or (_11685_, _11684_, _11681_);
  and (_11686_, _11685_, _02561_);
  or (_11687_, _08924_, _02561_);
  nand (_11688_, _11687_, _02983_);
  or (_11689_, _11688_, _11686_);
  nand (_11690_, _07610_, _02984_);
  and (_11691_, _11690_, _11689_);
  or (_11692_, _11691_, _03867_);
  and (_11693_, _05847_, _02858_);
  nand (_11694_, _07609_, _03867_);
  or (_11695_, _11694_, _11693_);
  and (_11696_, _11695_, _04303_);
  and (_11697_, _11696_, _11692_);
  or (_11698_, _11697_, _11651_);
  and (_11699_, _11698_, _05325_);
  nand (_11700_, _08923_, _02578_);
  nand (_11701_, _11700_, _05551_);
  or (_11702_, _11701_, _11699_);
  or (_11703_, _06158_, _05551_);
  and (_11704_, _11703_, _11702_);
  or (_11705_, _11704_, _02857_);
  or (_11706_, _05847_, _05558_);
  and (_11707_, _11706_, _02853_);
  and (_11708_, _11707_, _11705_);
  nor (_11709_, _05563_, _04787_);
  and (_11710_, _05694_, \oc8051_golden_model_1.B [6]);
  and (_11711_, _05703_, \oc8051_golden_model_1.ACC [6]);
  or (_11712_, _11711_, _11710_);
  and (_11713_, _05689_, \oc8051_golden_model_1.IP [6]);
  and (_11714_, _05699_, \oc8051_golden_model_1.PSW [6]);
  or (_11715_, _11714_, _11713_);
  or (_11716_, _11715_, _11712_);
  and (_11717_, _05681_, \oc8051_golden_model_1.TH1 [6]);
  and (_11718_, _05672_, \oc8051_golden_model_1.DPH [6]);
  or (_11719_, _11718_, _11717_);
  and (_11720_, _05749_, \oc8051_golden_model_1.DPL [6]);
  and (_11721_, _05667_, \oc8051_golden_model_1.TMOD [6]);
  or (_11722_, _11721_, _11720_);
  or (_11723_, _11722_, _11719_);
  or (_11724_, _11723_, _11716_);
  and (_11725_, _05720_, \oc8051_golden_model_1.TH0 [6]);
  and (_11726_, _05722_, \oc8051_golden_model_1.TL1 [6]);
  or (_11727_, _11726_, _11725_);
  and (_11728_, _05725_, \oc8051_golden_model_1.TCON [6]);
  and (_11729_, _05729_, \oc8051_golden_model_1.PCON [6]);
  or (_11730_, _11729_, _11728_);
  or (_11731_, _11730_, _11727_);
  and (_11732_, _05712_, \oc8051_golden_model_1.SBUF [6]);
  and (_11733_, _05714_, \oc8051_golden_model_1.SCON [6]);
  and (_11734_, _05708_, \oc8051_golden_model_1.IE [6]);
  or (_11735_, _11734_, _11733_);
  or (_11736_, _11735_, _11732_);
  and (_11737_, _05736_, \oc8051_golden_model_1.P0INREG [6]);
  and (_11738_, _05733_, \oc8051_golden_model_1.P1INREG [6]);
  and (_11739_, _05739_, \oc8051_golden_model_1.P2INREG [6]);
  and (_11740_, _05741_, \oc8051_golden_model_1.P3INREG [6]);
  or (_11741_, _11740_, _11739_);
  or (_11742_, _11741_, _11738_);
  or (_11743_, _11742_, _11737_);
  and (_11744_, _05747_, \oc8051_golden_model_1.SP [6]);
  and (_11745_, _05677_, \oc8051_golden_model_1.TL0 [6]);
  or (_11746_, _11745_, _11744_);
  or (_11747_, _11746_, _11743_);
  or (_11748_, _11747_, _11736_);
  or (_11749_, _11748_, _11731_);
  or (_11750_, _11749_, _11724_);
  nor (_11751_, _11750_, _11709_);
  nor (_11752_, _11751_, _02853_);
  or (_11753_, _11752_, _05562_);
  or (_11754_, _11753_, _11708_);
  and (_11755_, _05562_, _02932_);
  nor (_11756_, _11755_, _03885_);
  and (_11757_, _11756_, _11754_);
  not (_11758_, _05598_);
  and (_11759_, _11758_, _03885_);
  or (_11760_, _11759_, _02517_);
  or (_11761_, _11760_, _11757_);
  and (_11762_, _08924_, _02517_);
  nor (_11763_, _11762_, _05280_);
  and (_11764_, _11763_, _11761_);
  or (_11765_, _11764_, _11647_);
  and (_11766_, _11765_, _05278_);
  nor (_11767_, _04837_, _06833_);
  and (_11768_, _04837_, _06833_);
  nor (_11769_, _11768_, _11767_);
  and (_11770_, _11769_, _05277_);
  or (_11771_, _11770_, _11766_);
  and (_11772_, _11771_, _05276_);
  and (_11773_, _11645_, _05275_);
  or (_11774_, _11773_, _11772_);
  and (_11775_, _11774_, _05273_);
  and (_11776_, _11767_, _03891_);
  or (_11777_, _11776_, _02533_);
  or (_11778_, _11777_, _11775_);
  and (_11779_, _08924_, _02533_);
  nor (_11780_, _11779_, _05782_);
  and (_11781_, _11780_, _11778_);
  nor (_11782_, _11644_, _05788_);
  or (_11783_, _11782_, _05787_);
  or (_11784_, _11783_, _11781_);
  nand (_11785_, _11768_, _05787_);
  and (_11786_, _11785_, _05792_);
  and (_11787_, _11786_, _11784_);
  and (_11788_, _08923_, _02531_);
  or (_11789_, _11788_, _10977_);
  or (_11790_, _11789_, _10975_);
  or (_11791_, _11790_, _11787_);
  and (_11792_, _11791_, _11643_);
  or (_11793_, _11792_, _04085_);
  or (_11794_, _11642_, _04084_);
  and (_11795_, _11794_, _03910_);
  and (_11796_, _11795_, _11793_);
  or (_11797_, _11796_, _11640_);
  and (_11798_, _11797_, _05801_);
  or (_11799_, _11798_, _11637_);
  and (_11800_, _11799_, _06195_);
  and (_11801_, _09056_, _03004_);
  or (_11802_, _11801_, _02528_);
  or (_11803_, _11802_, _11800_);
  and (_11804_, _08924_, _02528_);
  nor (_11805_, _11804_, _03627_);
  and (_11806_, _11805_, _11803_);
  and (_11807_, _11648_, _03627_);
  nor (_11808_, _11807_, _11806_);
  nand (_11809_, _11808_, _06153_);
  nor (_11810_, _06165_, _06158_);
  nor (_11811_, _11810_, _06166_);
  and (_11812_, _11811_, _06149_);
  or (_11813_, _11812_, _06154_);
  and (_11814_, _11813_, _11809_);
  and (_11815_, _11811_, _11198_);
  or (_11816_, _11815_, _03926_);
  or (_11817_, _11816_, _11814_);
  and (_11818_, _11817_, _11634_);
  or (_11819_, _11818_, _03925_);
  nor (_11820_, _05253_, _04838_);
  nor (_11821_, _11820_, _05254_);
  or (_11822_, _11821_, _04176_);
  and (_11823_, _11822_, _04186_);
  and (_11824_, _11823_, _11819_);
  or (_11825_, _11824_, _11021_);
  and (_11826_, _11825_, _11631_);
  not (_11827_, _08882_);
  nor (_11828_, _11827_, _03004_);
  and (_11829_, _09015_, _03004_);
  or (_11830_, _11829_, _11828_);
  and (_11831_, _11830_, _04551_);
  and (_11832_, _11831_, _10597_);
  or (_32547_, _11832_, _11826_);
  or (_11833_, _10406_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_11834_, _11833_, _10415_);
  or (_11835_, _11021_, _06191_);
  and (_11836_, _11835_, _11834_);
  and (_11837_, _10597_, _06230_);
  or (_32549_, _11837_, _11836_);
  and (_11838_, _04559_, _04103_);
  and (_11839_, _11838_, _10402_);
  or (_11840_, _11839_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_11841_, _04244_);
  or (_11842_, _10413_, _11841_);
  or (_11843_, _11842_, _10409_);
  and (_11844_, _11843_, _11840_);
  not (_11845_, _11839_);
  or (_11846_, _11845_, _10591_);
  and (_11847_, _11846_, _11844_);
  and (_11848_, _04551_, _04244_);
  and (_11849_, _11848_, _10595_);
  and (_11850_, _11849_, _10601_);
  or (_32552_, _11850_, _11847_);
  or (_11851_, _11839_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_11852_, _11851_, _11843_);
  or (_11853_, _11845_, _10808_);
  and (_11854_, _11853_, _11852_);
  and (_11855_, _11849_, _10814_);
  or (_32553_, _11855_, _11854_);
  or (_11856_, _11839_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_11857_, _11856_, _11843_);
  or (_11858_, _11845_, _11011_);
  and (_11859_, _11858_, _11857_);
  and (_11860_, _11849_, _11017_);
  or (_32554_, _11860_, _11859_);
  or (_11861_, _11839_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_11862_, _11861_, _11843_);
  or (_11863_, _11845_, _11216_);
  and (_11864_, _11863_, _11862_);
  and (_11865_, _11849_, _11222_);
  or (_32556_, _11865_, _11864_);
  or (_11866_, _11839_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_11867_, _11866_, _11843_);
  or (_11868_, _11845_, _11420_);
  and (_11869_, _11868_, _11867_);
  and (_11870_, _11849_, _11427_);
  or (_32557_, _11870_, _11869_);
  or (_11871_, _11839_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_11872_, _11871_, _11843_);
  and (_11873_, _11620_, _04557_);
  and (_11874_, _11873_, _11617_);
  or (_11875_, _11845_, _11874_);
  and (_11876_, _11875_, _11872_);
  and (_11877_, _11849_, _11628_);
  or (_32558_, _11877_, _11876_);
  or (_11878_, _11839_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_11879_, _11878_, _11843_);
  or (_11880_, _11845_, _11824_);
  and (_11881_, _11880_, _11879_);
  and (_11882_, _11849_, _11831_);
  or (_32559_, _11882_, _11881_);
  or (_11883_, _11839_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_11884_, _11883_, _11843_);
  or (_11885_, _11845_, _06192_);
  and (_11886_, _11885_, _11884_);
  and (_11887_, _11849_, _06230_);
  or (_32560_, _11887_, _11886_);
  and (_11888_, _04188_, _03932_);
  and (_11889_, _11888_, _10402_);
  not (_11890_, _11889_);
  or (_11891_, _11890_, _10591_);
  or (_11892_, _11889_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_11893_, _05403_);
  or (_11894_, _10413_, _11893_);
  or (_11895_, _11894_, _10409_);
  and (_11896_, _11895_, _11892_);
  and (_11897_, _11896_, _11891_);
  and (_11898_, _05403_, _04551_);
  and (_11899_, _11898_, _10595_);
  and (_11900_, _11899_, _10601_);
  or (_32564_, _11900_, _11897_);
  or (_11901_, _11890_, _10808_);
  or (_11902_, _11889_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_11903_, _11902_, _11895_);
  and (_11904_, _11903_, _11901_);
  and (_11905_, _11899_, _10814_);
  or (_32565_, _11905_, _11904_);
  or (_11906_, _11890_, _11011_);
  or (_11907_, _11889_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_11908_, _11907_, _11895_);
  and (_11909_, _11908_, _11906_);
  and (_11910_, _11899_, _11017_);
  or (_32566_, _11910_, _11909_);
  or (_11911_, _11890_, _11216_);
  or (_11912_, _11889_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_11913_, _11912_, _11895_);
  and (_11914_, _11913_, _11911_);
  and (_11915_, _11899_, _11222_);
  or (_32567_, _11915_, _11914_);
  or (_11916_, _11890_, _11420_);
  or (_11917_, _11889_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_11918_, _11917_, _11895_);
  and (_11919_, _11918_, _11916_);
  and (_11920_, _11899_, _11427_);
  or (_32568_, _11920_, _11919_);
  or (_11921_, _11890_, _11622_);
  or (_11922_, _11889_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_11923_, _11922_, _11895_);
  and (_11924_, _11923_, _11921_);
  and (_11925_, _11899_, _11628_);
  or (_32570_, _11925_, _11924_);
  or (_11926_, _11890_, _11824_);
  or (_11927_, _11889_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_11928_, _11927_, _11895_);
  and (_11929_, _11928_, _11926_);
  and (_11930_, _11899_, _11831_);
  or (_32571_, _11930_, _11929_);
  or (_11931_, _11889_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_11932_, _11931_, _11895_);
  or (_11933_, _11890_, _06192_);
  and (_11934_, _11933_, _11932_);
  and (_11935_, _11899_, _06230_);
  or (_32572_, _11935_, _11934_);
  and (_11936_, _10402_, _04561_);
  or (_11937_, _11936_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_11938_, _03938_);
  or (_11939_, _10413_, _11938_);
  or (_11940_, _11939_, _10409_);
  and (_11941_, _11940_, _11937_);
  not (_11942_, _11936_);
  or (_11943_, _11942_, _10591_);
  and (_11944_, _11943_, _11941_);
  and (_11945_, _04551_, _03938_);
  and (_11946_, _11945_, _10595_);
  and (_11947_, _11946_, _10601_);
  or (_32575_, _11947_, _11944_);
  or (_11948_, _11936_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_11949_, _11948_, _11940_);
  or (_11950_, _11942_, _10808_);
  and (_11951_, _11950_, _11949_);
  and (_11952_, _11946_, _10814_);
  or (_32576_, _11952_, _11951_);
  or (_11953_, _11936_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_11954_, _11953_, _11940_);
  or (_11955_, _11942_, _11011_);
  and (_11956_, _11955_, _11954_);
  and (_11957_, _11946_, _11017_);
  or (_32577_, _11957_, _11956_);
  or (_11958_, _11936_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_11959_, _11958_, _11940_);
  or (_11960_, _11942_, _11216_);
  and (_11961_, _11960_, _11959_);
  and (_11962_, _11946_, _11222_);
  or (_32579_, _11962_, _11961_);
  or (_11963_, _11936_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_11964_, _11963_, _11940_);
  or (_11965_, _11942_, _11420_);
  and (_11966_, _11965_, _11964_);
  and (_11967_, _11946_, _11427_);
  or (_32580_, _11967_, _11966_);
  or (_11968_, _11942_, _11874_);
  or (_11969_, _11936_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_11970_, _11969_, _11940_);
  and (_11971_, _11970_, _11968_);
  and (_11972_, _11946_, _11628_);
  or (_32581_, _11972_, _11971_);
  or (_11973_, _11936_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_11974_, _11973_, _11940_);
  or (_11975_, _11942_, _11824_);
  and (_11976_, _11975_, _11974_);
  and (_11977_, _11946_, _11831_);
  or (_32582_, _11977_, _11976_);
  or (_11978_, _11936_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_11979_, _11978_, _11940_);
  or (_11980_, _11942_, _06192_);
  and (_11981_, _11980_, _11979_);
  and (_11982_, _11946_, _06230_);
  or (_32583_, _11982_, _11981_);
  and (_11983_, _10401_, _04359_);
  nand (_11984_, _11983_, _10418_);
  or (_11985_, _11984_, _10591_);
  not (_11986_, _04546_);
  and (_11987_, _10411_, _11986_);
  and (_11988_, _11987_, _03939_);
  not (_11989_, _11988_);
  nand (_11990_, _11984_, _03780_);
  and (_11991_, _11990_, _11989_);
  and (_11992_, _11991_, _11985_);
  and (_11993_, _11988_, _10601_);
  or (_32587_, _11993_, _11992_);
  and (_11994_, _11988_, _10814_);
  and (_11995_, _04536_, _04359_);
  and (_11996_, _11995_, _10405_);
  or (_11997_, _11996_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_11998_, _11997_, _11989_);
  or (_11999_, _11984_, _10808_);
  and (_12000_, _11999_, _11998_);
  or (_32588_, _12000_, _11994_);
  or (_12001_, _11996_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_12002_, _12001_, _11989_);
  or (_12003_, _11984_, _11011_);
  and (_12004_, _12003_, _12002_);
  and (_12005_, _11988_, _11017_);
  or (_32589_, _12005_, _12004_);
  or (_12006_, _11996_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_12007_, _12006_, _11989_);
  not (_12008_, _11996_);
  or (_12009_, _12008_, _11216_);
  and (_12010_, _12009_, _12007_);
  and (_12011_, _11988_, _11222_);
  or (_32590_, _12011_, _12010_);
  or (_12012_, _11996_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_12013_, _12012_, _11989_);
  or (_12014_, _11984_, _11420_);
  and (_12015_, _12014_, _12013_);
  and (_12016_, _11988_, _11427_);
  or (_32591_, _12016_, _12015_);
  or (_12017_, _11996_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_12018_, _12017_, _11989_);
  or (_12019_, _12008_, _11622_);
  and (_12020_, _12019_, _12018_);
  and (_12021_, _11988_, _11628_);
  or (_32592_, _12021_, _12020_);
  and (_12022_, _11988_, _11831_);
  or (_12023_, _11996_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_12024_, _12023_, _11989_);
  or (_12025_, _12008_, _11824_);
  and (_12026_, _12025_, _12024_);
  or (_32593_, _12026_, _12022_);
  and (_12027_, _11988_, _06230_);
  or (_12028_, _11996_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_12029_, _12028_, _11989_);
  or (_12030_, _11984_, _06192_);
  and (_12031_, _12030_, _12029_);
  or (_32594_, _12031_, _12027_);
  and (_12032_, _11983_, _11838_);
  not (_12033_, _12032_);
  or (_12034_, _12033_, _10591_);
  and (_12035_, _10594_, _11986_);
  and (_12036_, _12035_, _04244_);
  nor (_12037_, _12032_, \oc8051_golden_model_1.IRAM[5] [0]);
  nor (_12038_, _12037_, _12036_);
  and (_12039_, _12038_, _12034_);
  and (_12040_, _12036_, _10601_);
  or (_32598_, _12040_, _12039_);
  nand (_12041_, _11987_, _04244_);
  and (_12042_, _10404_, _04103_);
  and (_12043_, _11995_, _12042_);
  or (_12044_, _12043_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_12045_, _12044_, _12041_);
  or (_12046_, _12033_, _10808_);
  and (_12047_, _12046_, _12045_);
  and (_12048_, _12036_, _10814_);
  or (_32599_, _12048_, _12047_);
  or (_12049_, _12043_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_12050_, _12049_, _12041_);
  or (_12051_, _12033_, _11011_);
  and (_12052_, _12051_, _12050_);
  and (_12053_, _12036_, _11017_);
  or (_32600_, _12053_, _12052_);
  or (_12054_, _12043_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_12055_, _12054_, _12041_);
  not (_12056_, _12043_);
  or (_12057_, _12056_, _11216_);
  and (_12058_, _12057_, _12055_);
  and (_12059_, _12036_, _11222_);
  or (_32601_, _12059_, _12058_);
  or (_12060_, _12043_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_12061_, _12060_, _12041_);
  or (_12062_, _12033_, _11420_);
  and (_12063_, _12062_, _12061_);
  and (_12064_, _12036_, _11427_);
  or (_32602_, _12064_, _12063_);
  or (_12065_, _12043_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_12066_, _12065_, _12041_);
  or (_12067_, _12056_, _11622_);
  and (_12068_, _12067_, _12066_);
  and (_12069_, _12036_, _11628_);
  or (_32603_, _12069_, _12068_);
  or (_12070_, _12043_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_12071_, _12070_, _12041_);
  or (_12072_, _12056_, _11824_);
  and (_12073_, _12072_, _12071_);
  and (_12074_, _12036_, _11831_);
  or (_32604_, _12074_, _12073_);
  or (_12075_, _12043_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_12076_, _12075_, _12041_);
  or (_12077_, _12033_, _06192_);
  and (_12078_, _12077_, _12076_);
  and (_12079_, _12036_, _06230_);
  or (_32605_, _12079_, _12078_);
  and (_12080_, _11983_, _11888_);
  not (_12081_, _12080_);
  or (_12082_, _12081_, _10591_);
  or (_12083_, _12080_, \oc8051_golden_model_1.IRAM[6] [0]);
  nand (_12084_, _11987_, _05403_);
  and (_12085_, _12084_, _12083_);
  and (_12086_, _12085_, _12082_);
  and (_12087_, _12035_, _05403_);
  and (_12088_, _12087_, _10601_);
  or (_32608_, _12088_, _12086_);
  or (_12089_, _12080_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_12090_, _12089_, _12084_);
  or (_12091_, _12081_, _10808_);
  and (_12092_, _12091_, _12090_);
  and (_12093_, _12087_, _10814_);
  or (_32609_, _12093_, _12092_);
  or (_12094_, _12081_, _11011_);
  or (_12095_, _12080_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_12096_, _12095_, _12084_);
  and (_12097_, _12096_, _12094_);
  and (_12098_, _12087_, _11017_);
  or (_32610_, _12098_, _12097_);
  nand (_12099_, _11995_, _11888_);
  or (_12100_, _12099_, _11216_);
  or (_12101_, _12080_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_12102_, _12101_, _12084_);
  and (_12103_, _12102_, _12100_);
  and (_12104_, _12087_, _11222_);
  or (_32611_, _12104_, _12103_);
  or (_12105_, _12081_, _11420_);
  or (_12106_, _12080_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_12107_, _12106_, _12084_);
  and (_12108_, _12107_, _12105_);
  and (_12109_, _12087_, _11427_);
  or (_32613_, _12109_, _12108_);
  or (_12110_, _12099_, _11622_);
  or (_12111_, _12080_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_12112_, _12111_, _12084_);
  and (_12113_, _12112_, _12110_);
  and (_12114_, _12087_, _11628_);
  or (_32614_, _12114_, _12113_);
  or (_12115_, _12080_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_12116_, _12115_, _12084_);
  or (_12117_, _12081_, _11824_);
  and (_12118_, _12117_, _12116_);
  and (_12119_, _12087_, _11831_);
  or (_32615_, _12119_, _12118_);
  or (_12120_, _12081_, _06192_);
  or (_12121_, _12080_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_12122_, _12121_, _12084_);
  and (_12123_, _12122_, _12120_);
  and (_12124_, _12087_, _06230_);
  or (_32616_, _12124_, _12123_);
  and (_12125_, _11983_, _04561_);
  not (_12126_, _12125_);
  or (_12127_, _12126_, _10591_);
  and (_12128_, _11987_, _03938_);
  not (_12129_, _12128_);
  or (_12130_, _12125_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_12131_, _12130_, _12129_);
  and (_12132_, _12131_, _12127_);
  and (_12133_, _12128_, _10601_);
  or (_32619_, _12133_, _12132_);
  and (_12134_, _11995_, _04189_);
  or (_12135_, _12134_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_12136_, _12135_, _12129_);
  or (_12137_, _12126_, _10808_);
  and (_12138_, _12137_, _12136_);
  and (_12139_, _12128_, _10814_);
  or (_32620_, _12139_, _12138_);
  or (_12140_, _12134_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_12141_, _12140_, _12129_);
  or (_12142_, _12126_, _11011_);
  and (_12143_, _12142_, _12141_);
  and (_12144_, _12128_, _11017_);
  or (_32621_, _12144_, _12143_);
  or (_12145_, _12134_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_12146_, _12145_, _12129_);
  not (_12147_, _12134_);
  or (_12148_, _12147_, _11216_);
  and (_12149_, _12148_, _12146_);
  and (_12150_, _12128_, _11222_);
  or (_32623_, _12150_, _12149_);
  or (_12151_, _12134_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_12152_, _12151_, _12129_);
  or (_12153_, _12126_, _11420_);
  and (_12154_, _12153_, _12152_);
  and (_12155_, _12128_, _11427_);
  or (_32624_, _12155_, _12154_);
  or (_12156_, _12134_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_12157_, _12156_, _12129_);
  or (_12158_, _12147_, _11622_);
  and (_12159_, _12158_, _12157_);
  and (_12160_, _12128_, _11628_);
  or (_32625_, _12160_, _12159_);
  or (_12161_, _12134_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_12162_, _12161_, _12129_);
  or (_12163_, _12147_, _11824_);
  and (_12164_, _12163_, _12162_);
  and (_12165_, _12128_, _11831_);
  or (_32626_, _12165_, _12164_);
  or (_12166_, _12134_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_12167_, _12166_, _12129_);
  or (_12168_, _12126_, _06192_);
  and (_12169_, _12168_, _12167_);
  and (_12170_, _12128_, _06230_);
  or (_32627_, _12170_, _12169_);
  and (_12171_, _04564_, _04535_);
  and (_12172_, _12171_, _10418_);
  or (_12173_, _12172_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_12174_, _04543_);
  and (_12175_, _04552_, _12174_);
  and (_12176_, _12175_, _03939_);
  not (_12177_, _12176_);
  and (_12178_, _12177_, _12173_);
  not (_12179_, _12172_);
  or (_12180_, _12179_, _10591_);
  and (_12181_, _12180_, _12178_);
  and (_12182_, _12176_, _10601_);
  or (_32631_, _12182_, _12181_);
  or (_12183_, _12172_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_12184_, _12183_, _12177_);
  or (_12185_, _12179_, _10808_);
  and (_12186_, _12185_, _12184_);
  and (_12187_, _12176_, _10814_);
  or (_32632_, _12187_, _12186_);
  or (_12188_, _12172_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_12189_, _12188_, _12177_);
  or (_12190_, _12179_, _11011_);
  and (_12191_, _12190_, _12189_);
  and (_12192_, _12176_, _11017_);
  or (_32633_, _12192_, _12191_);
  or (_12193_, _12172_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_12194_, _12193_, _12177_);
  or (_12195_, _12179_, _11216_);
  and (_12196_, _12195_, _12194_);
  and (_12197_, _12176_, _11222_);
  or (_32634_, _12197_, _12196_);
  or (_12198_, _12172_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_12199_, _12198_, _12177_);
  or (_12200_, _12179_, _11420_);
  and (_12201_, _12200_, _12199_);
  and (_12202_, _12176_, _11427_);
  or (_32635_, _12202_, _12201_);
  or (_12203_, _12172_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_12204_, _12203_, _12177_);
  or (_12205_, _12179_, _11874_);
  and (_12206_, _12205_, _12204_);
  and (_12207_, _12176_, _11628_);
  or (_32637_, _12207_, _12206_);
  or (_12208_, _12172_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_12209_, _12208_, _12177_);
  or (_12210_, _12179_, _11824_);
  and (_12211_, _12210_, _12209_);
  and (_12212_, _12176_, _11831_);
  or (_32638_, _12212_, _12211_);
  or (_12213_, _12172_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_12214_, _12213_, _12177_);
  or (_12215_, _12179_, _06192_);
  and (_12216_, _12215_, _12214_);
  and (_12217_, _12176_, _06230_);
  or (_32639_, _12217_, _12216_);
  and (_12218_, _12171_, _11838_);
  or (_12219_, _12218_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_12220_, _10412_, _04245_);
  and (_12221_, _12220_, _12219_);
  not (_12222_, _12218_);
  or (_12223_, _12222_, _10591_);
  and (_12224_, _12223_, _12221_);
  and (_12225_, _12175_, _04244_);
  and (_12226_, _12225_, _10601_);
  or (_32642_, _12226_, _12224_);
  or (_12227_, _12218_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_12228_, _12227_, _12220_);
  or (_12229_, _12222_, _10808_);
  and (_12230_, _12229_, _12228_);
  and (_12231_, _12225_, _10814_);
  or (_32643_, _12231_, _12230_);
  or (_12232_, _12218_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_12233_, _12232_, _12220_);
  or (_12234_, _12222_, _11011_);
  and (_12235_, _12234_, _12233_);
  and (_12236_, _12225_, _11017_);
  or (_32644_, _12236_, _12235_);
  or (_12237_, _12218_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_12238_, _12237_, _12220_);
  or (_12239_, _12222_, _11216_);
  and (_12240_, _12239_, _12238_);
  and (_12241_, _12225_, _11222_);
  or (_32645_, _12241_, _12240_);
  or (_12242_, _12218_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_12243_, _12242_, _12220_);
  or (_12244_, _12222_, _11420_);
  and (_12245_, _12244_, _12243_);
  and (_12246_, _12225_, _11427_);
  or (_32647_, _12246_, _12245_);
  or (_12247_, _12218_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_12248_, _12247_, _12220_);
  or (_12249_, _12222_, _11874_);
  and (_12250_, _12249_, _12248_);
  and (_12251_, _12225_, _11628_);
  or (_32648_, _12251_, _12250_);
  or (_12252_, _12218_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_12253_, _12252_, _12220_);
  or (_12254_, _12222_, _11824_);
  and (_12255_, _12254_, _12253_);
  and (_12256_, _12225_, _11831_);
  or (_32649_, _12256_, _12255_);
  or (_12257_, _12218_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_12258_, _12257_, _12220_);
  or (_12259_, _12222_, _06192_);
  and (_12260_, _12259_, _12258_);
  and (_12261_, _12225_, _06230_);
  or (_32650_, _12261_, _12260_);
  and (_12262_, _12171_, _11888_);
  or (_12263_, _12262_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_12264_, _12175_, _05403_);
  not (_12265_, _12264_);
  and (_12266_, _12265_, _12263_);
  not (_12267_, _12262_);
  or (_12268_, _12267_, _10591_);
  and (_12269_, _12268_, _12266_);
  and (_12270_, _12264_, _10601_);
  or (_32653_, _12270_, _12269_);
  or (_12271_, _12262_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_12272_, _12271_, _12265_);
  or (_12273_, _12267_, _10808_);
  and (_12274_, _12273_, _12272_);
  and (_12275_, _12264_, _10814_);
  or (_32654_, _12275_, _12274_);
  or (_12276_, _12262_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_12277_, _12276_, _12265_);
  or (_12278_, _12267_, _11011_);
  and (_12279_, _12278_, _12277_);
  and (_12280_, _12264_, _11017_);
  or (_32655_, _12280_, _12279_);
  or (_12281_, _12262_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_12282_, _12281_, _12265_);
  or (_12283_, _12267_, _11216_);
  and (_12284_, _12283_, _12282_);
  and (_12285_, _12264_, _11222_);
  or (_32656_, _12285_, _12284_);
  or (_12286_, _12267_, _11420_);
  or (_12287_, _12262_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_12288_, _12287_, _12265_);
  and (_12289_, _12288_, _12286_);
  and (_12290_, _12264_, _11427_);
  or (_32658_, _12290_, _12289_);
  or (_12291_, _12267_, _11874_);
  or (_12292_, _12262_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_12293_, _12292_, _12265_);
  and (_12294_, _12293_, _12291_);
  and (_12295_, _12264_, _11628_);
  or (_32659_, _12295_, _12294_);
  or (_12296_, _12262_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_12297_, _12296_, _12265_);
  or (_12298_, _12267_, _11824_);
  and (_12299_, _12298_, _12297_);
  and (_12300_, _12264_, _11831_);
  or (_32660_, _12300_, _12299_);
  or (_12301_, _12267_, _06192_);
  or (_12302_, _12262_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_12303_, _12302_, _12265_);
  and (_12304_, _12303_, _12301_);
  and (_12305_, _12264_, _06230_);
  or (_32661_, _12305_, _12304_);
  and (_12306_, _12171_, _04561_);
  or (_12307_, _12306_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_12308_, _12175_, _03938_);
  not (_12309_, _12308_);
  and (_12310_, _12309_, _12307_);
  not (_12311_, _12306_);
  or (_12312_, _12311_, _10591_);
  and (_12313_, _12312_, _12310_);
  and (_12314_, _12308_, _10601_);
  or (_32664_, _12314_, _12313_);
  or (_12315_, _12306_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_12316_, _12315_, _12309_);
  or (_12317_, _12311_, _10808_);
  and (_12318_, _12317_, _12316_);
  and (_12319_, _12308_, _10814_);
  or (_32665_, _12319_, _12318_);
  or (_12320_, _12306_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_12321_, _12320_, _12309_);
  or (_12322_, _12311_, _11011_);
  and (_12323_, _12322_, _12321_);
  and (_12324_, _12308_, _11017_);
  or (_32666_, _12324_, _12323_);
  or (_12325_, _12306_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_12326_, _12325_, _12309_);
  or (_12327_, _12311_, _11216_);
  and (_12328_, _12327_, _12326_);
  and (_12329_, _12308_, _11222_);
  or (_32668_, _12329_, _12328_);
  or (_12330_, _12306_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_12331_, _12330_, _12309_);
  or (_12332_, _12311_, _11420_);
  and (_12333_, _12332_, _12331_);
  and (_12334_, _12308_, _11427_);
  or (_32669_, _12334_, _12333_);
  or (_12335_, _12306_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_12336_, _12335_, _12309_);
  or (_12337_, _12311_, _11874_);
  and (_12338_, _12337_, _12336_);
  and (_12339_, _12308_, _11628_);
  or (_32670_, _12339_, _12338_);
  or (_12340_, _12306_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_12341_, _12340_, _12309_);
  or (_12342_, _12311_, _11824_);
  and (_12343_, _12342_, _12341_);
  and (_12344_, _12308_, _11831_);
  or (_32671_, _12344_, _12343_);
  or (_12345_, _12306_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_12346_, _12345_, _12309_);
  or (_12347_, _12311_, _06192_);
  and (_12348_, _12347_, _12346_);
  and (_12349_, _12308_, _06230_);
  or (_32672_, _12349_, _12348_);
  not (_12350_, _10418_);
  or (_12351_, _12350_, _04565_);
  or (_12352_, _12351_, _10591_);
  and (_12353_, _04553_, _03939_);
  not (_12354_, _12353_);
  nand (_12355_, _12351_, _03808_);
  and (_12356_, _12355_, _12354_);
  and (_12357_, _12356_, _12352_);
  and (_12358_, _12353_, _10601_);
  or (_32675_, _12358_, _12357_);
  and (_12359_, _10405_, _04538_);
  or (_12360_, _12359_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_12361_, _12360_, _12354_);
  or (_12362_, _12351_, _10808_);
  and (_12363_, _12362_, _12361_);
  and (_12364_, _12353_, _10814_);
  or (_32676_, _12364_, _12363_);
  or (_12365_, _12359_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_12366_, _12365_, _12354_);
  or (_12367_, _12351_, _11011_);
  and (_12368_, _12367_, _12366_);
  and (_12369_, _12353_, _11017_);
  or (_32678_, _12369_, _12368_);
  or (_12370_, _12359_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_12371_, _12370_, _12354_);
  or (_12372_, _12351_, _11216_);
  and (_12373_, _12372_, _12371_);
  and (_12374_, _12353_, _11222_);
  or (_32679_, _12374_, _12373_);
  or (_12375_, _12351_, _11420_);
  or (_12376_, _12359_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_12377_, _12376_, _12354_);
  and (_12378_, _12377_, _12375_);
  and (_12379_, _12353_, _11427_);
  or (_32680_, _12379_, _12378_);
  or (_12380_, _12351_, _11874_);
  or (_12381_, _12359_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_12382_, _12381_, _12354_);
  and (_12383_, _12382_, _12380_);
  and (_12384_, _12353_, _11628_);
  or (_32681_, _12384_, _12383_);
  or (_12385_, _12359_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_12386_, _12385_, _12354_);
  or (_12387_, _12351_, _11824_);
  and (_12388_, _12387_, _12386_);
  and (_12389_, _12353_, _11831_);
  or (_32682_, _12389_, _12388_);
  or (_12390_, _12359_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_12391_, _12390_, _12354_);
  or (_12392_, _12351_, _06192_);
  and (_12393_, _12392_, _12391_);
  and (_12394_, _12353_, _06230_);
  or (_32684_, _12394_, _12393_);
  and (_12395_, _10411_, _04546_);
  and (_12396_, _12395_, _04244_);
  not (_12397_, _12396_);
  and (_12398_, _12042_, _04538_);
  or (_12399_, _12398_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_12400_, _12399_, _12397_);
  not (_12401_, _11838_);
  or (_12402_, _12401_, _04565_);
  or (_12403_, _12402_, _10591_);
  and (_12404_, _12403_, _12400_);
  and (_12405_, _04553_, _04244_);
  and (_12406_, _12405_, _10601_);
  or (_32686_, _12406_, _12404_);
  or (_12407_, _12398_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_12408_, _12407_, _12397_);
  or (_12409_, _12402_, _10808_);
  and (_12410_, _12409_, _12408_);
  and (_12411_, _12405_, _10814_);
  or (_32688_, _12411_, _12410_);
  or (_12412_, _12398_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_12413_, _12412_, _12397_);
  or (_12414_, _12402_, _11011_);
  and (_12415_, _12414_, _12413_);
  and (_12416_, _12405_, _11017_);
  or (_32689_, _12416_, _12415_);
  or (_12417_, _12398_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_12418_, _12417_, _12397_);
  or (_12419_, _12402_, _11216_);
  and (_12420_, _12419_, _12418_);
  and (_12421_, _12405_, _11222_);
  or (_32690_, _12421_, _12420_);
  or (_12422_, _12398_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_12423_, _12422_, _12397_);
  or (_12424_, _12402_, _11420_);
  and (_12425_, _12424_, _12423_);
  and (_12426_, _12405_, _11427_);
  or (_32691_, _12426_, _12425_);
  or (_12427_, _12398_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_12428_, _12427_, _12397_);
  or (_12429_, _12402_, _11874_);
  and (_12430_, _12429_, _12428_);
  and (_12431_, _12405_, _11628_);
  or (_32692_, _12431_, _12430_);
  or (_12432_, _12398_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_12433_, _12432_, _12397_);
  or (_12434_, _12402_, _11824_);
  and (_12435_, _12434_, _12433_);
  and (_12436_, _12405_, _11831_);
  or (_32694_, _12436_, _12435_);
  or (_12437_, _12398_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_12438_, _12437_, _12397_);
  or (_12439_, _12402_, _06192_);
  and (_12440_, _12439_, _12438_);
  and (_12441_, _12405_, _06230_);
  or (_32695_, _12441_, _12440_);
  and (_12442_, _11888_, _04538_);
  or (_12443_, _12442_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_12444_, _05403_, _04553_);
  not (_12445_, _12444_);
  and (_12446_, _12445_, _12443_);
  not (_12447_, _11888_);
  or (_12448_, _12447_, _04565_);
  or (_12449_, _12448_, _10591_);
  and (_12450_, _12449_, _12446_);
  and (_12451_, _12444_, _10601_);
  or (_32697_, _12451_, _12450_);
  or (_12452_, _12442_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_12453_, _12452_, _12445_);
  or (_12454_, _12448_, _10808_);
  and (_12455_, _12454_, _12453_);
  and (_12456_, _12444_, _10814_);
  or (_32699_, _12456_, _12455_);
  or (_12457_, _12442_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_12458_, _12457_, _12445_);
  or (_12459_, _12448_, _11011_);
  and (_12460_, _12459_, _12458_);
  and (_12461_, _12444_, _11017_);
  or (_32700_, _12461_, _12460_);
  or (_12462_, _12442_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_12463_, _12462_, _12445_);
  or (_12464_, _12448_, _11216_);
  and (_12465_, _12464_, _12463_);
  and (_12466_, _12444_, _11222_);
  or (_32701_, _12466_, _12465_);
  or (_12467_, _12442_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_12468_, _12467_, _12445_);
  or (_12469_, _12448_, _11420_);
  and (_12470_, _12469_, _12468_);
  and (_12471_, _12444_, _11427_);
  or (_32702_, _12471_, _12470_);
  or (_12472_, _12442_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_12473_, _12472_, _12445_);
  or (_12474_, _12448_, _11874_);
  and (_12475_, _12474_, _12473_);
  and (_12476_, _12444_, _11628_);
  or (_32703_, _12476_, _12475_);
  or (_12477_, _12442_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_12478_, _12477_, _12445_);
  or (_12479_, _12448_, _11824_);
  and (_12480_, _12479_, _12478_);
  and (_12481_, _12444_, _11831_);
  or (_32704_, _12481_, _12480_);
  or (_12482_, _12442_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_12483_, _12482_, _12445_);
  or (_12484_, _12448_, _06192_);
  and (_12485_, _12484_, _12483_);
  and (_12486_, _12444_, _06230_);
  or (_32705_, _12486_, _12485_);
  or (_12487_, _10591_, _04566_);
  or (_12488_, _04539_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_12489_, _12488_, _04555_);
  and (_12490_, _12489_, _12487_);
  and (_12491_, _10601_, _04554_);
  or (_32708_, _12491_, _12490_);
  or (_12492_, _04539_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_12493_, _12492_, _04555_);
  or (_12494_, _10808_, _04566_);
  and (_12495_, _12494_, _12493_);
  and (_12496_, _10814_, _04554_);
  or (_32709_, _12496_, _12495_);
  or (_12497_, _04539_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_12498_, _12497_, _04555_);
  or (_12499_, _11011_, _04566_);
  and (_12500_, _12499_, _12498_);
  and (_12501_, _11017_, _04554_);
  or (_32710_, _12501_, _12500_);
  or (_12502_, _04539_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_12503_, _12502_, _04555_);
  or (_12504_, _11216_, _04566_);
  and (_12505_, _12504_, _12503_);
  and (_12506_, _11222_, _04554_);
  or (_32711_, _12506_, _12505_);
  or (_12507_, _11420_, _04566_);
  or (_12508_, _04539_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_12509_, _12508_, _04555_);
  and (_12510_, _12509_, _12507_);
  and (_12511_, _11427_, _04554_);
  or (_32712_, _12511_, _12510_);
  or (_12512_, _04539_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_12513_, _12512_, _04555_);
  or (_12514_, _11874_, _04566_);
  and (_12515_, _12514_, _12513_);
  and (_12516_, _11628_, _04554_);
  or (_32713_, _12516_, _12515_);
  or (_12517_, _04539_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_12518_, _12517_, _04555_);
  or (_12519_, _11824_, _04566_);
  and (_12520_, _12519_, _12518_);
  and (_12521_, _11831_, _04554_);
  or (_32715_, _12521_, _12520_);
  nor (_12522_, _34698_, _06820_);
  nor (_12523_, _04705_, _06820_);
  and (_12524_, _10546_, _04705_);
  or (_12525_, _12524_, _12523_);
  and (_12526_, _12525_, _03130_);
  and (_12527_, _04705_, _05566_);
  or (_12528_, _12527_, _12523_);
  or (_12529_, _12528_, _03884_);
  and (_12530_, _04705_, _03817_);
  or (_12531_, _12530_, _12523_);
  or (_12532_, _12531_, _06241_);
  and (_12533_, _05044_, _04705_);
  or (_12534_, _12533_, _12523_);
  or (_12535_, _12534_, _03821_);
  and (_12536_, _04705_, \oc8051_golden_model_1.ACC [0]);
  or (_12537_, _12536_, _12523_);
  and (_12538_, _12537_, _03825_);
  nor (_12539_, _03825_, _06820_);
  or (_12540_, _12539_, _02952_);
  or (_12541_, _12540_, _12538_);
  and (_12542_, _12541_, _02892_);
  and (_12543_, _12542_, _12535_);
  and (_12544_, _10429_, _05338_);
  nor (_12545_, _05338_, _06820_);
  or (_12546_, _12545_, _12544_);
  and (_12547_, _12546_, _02891_);
  or (_12548_, _12547_, _12543_);
  and (_12549_, _12548_, _03327_);
  and (_12550_, _12531_, _02947_);
  or (_12551_, _12550_, _02950_);
  or (_12552_, _12551_, _12549_);
  or (_12553_, _12537_, _02959_);
  and (_12554_, _12553_, _02888_);
  and (_12555_, _12554_, _12552_);
  and (_12556_, _12523_, _02887_);
  or (_12557_, _12556_, _02880_);
  or (_12558_, _12557_, _12555_);
  or (_12559_, _12534_, _02881_);
  and (_12560_, _12559_, _12558_);
  or (_12561_, _12560_, _06271_);
  nor (_12562_, _06754_, _06752_);
  nor (_12563_, _12562_, _06755_);
  or (_12564_, _12563_, _06277_);
  and (_12565_, _12564_, _02875_);
  and (_12566_, _12565_, _12561_);
  nor (_12567_, _10473_, _06794_);
  or (_12568_, _12567_, _12545_);
  and (_12569_, _12568_, _02874_);
  or (_12570_, _12569_, _06793_);
  or (_12571_, _12570_, _12566_);
  and (_12572_, _12571_, _12532_);
  or (_12573_, _12572_, _02855_);
  and (_12574_, _06174_, _04705_);
  or (_12575_, _12523_, _02856_);
  or (_12576_, _12575_, _12574_);
  and (_12577_, _12576_, _12573_);
  or (_12578_, _12577_, _02576_);
  nor (_12579_, _10530_, _06235_);
  or (_12580_, _12523_, _02851_);
  or (_12581_, _12580_, _12579_);
  and (_12582_, _12581_, _06813_);
  and (_12583_, _12582_, _12578_);
  nor (_12584_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_12585_, _12584_, _06732_);
  or (_12586_, _07164_, _12585_);
  nand (_12587_, _07164_, _02549_);
  and (_12588_, _12587_, _06807_);
  and (_12589_, _12588_, _12586_);
  or (_12590_, _12589_, _03014_);
  or (_12591_, _12590_, _12583_);
  and (_12592_, _12591_, _12529_);
  or (_12593_, _12592_, _03021_);
  and (_12594_, _10425_, _04705_);
  or (_12595_, _12523_, _05279_);
  or (_12596_, _12595_, _12594_);
  and (_12597_, _12596_, _03131_);
  and (_12598_, _12597_, _12593_);
  or (_12599_, _12598_, _12526_);
  and (_12600_, _12599_, _05274_);
  nand (_12601_, _12528_, _03020_);
  nor (_12602_, _12601_, _12533_);
  or (_12603_, _12602_, _12600_);
  and (_12604_, _12603_, _03140_);
  or (_12605_, _12523_, _09183_);
  and (_12606_, _12537_, _03139_);
  and (_12607_, _12606_, _12605_);
  or (_12608_, _12607_, _03036_);
  or (_12609_, _12608_, _12604_);
  nor (_12610_, _10423_, _06235_);
  or (_12611_, _12523_, _05781_);
  or (_12612_, _12611_, _12610_);
  and (_12613_, _12612_, _05786_);
  and (_12614_, _12613_, _12609_);
  nor (_12615_, _10421_, _06235_);
  or (_12616_, _12615_, _12523_);
  and (_12617_, _12616_, _03127_);
  or (_12618_, _12617_, _03166_);
  or (_12619_, _12618_, _12614_);
  or (_12620_, _12534_, _03563_);
  and (_12621_, _12620_, _02501_);
  and (_12622_, _12621_, _12619_);
  and (_12623_, _12523_, _02500_);
  or (_12624_, _12623_, _03174_);
  or (_12625_, _12624_, _12622_);
  or (_12627_, _12534_, _03178_);
  and (_12628_, _12627_, _34698_);
  and (_12629_, _12628_, _12625_);
  or (_12630_, _12629_, _12522_);
  and (_35155_, _12630_, _36029_);
  nor (_12631_, _34698_, _06814_);
  or (_12632_, _04705_, \oc8051_golden_model_1.B [1]);
  nand (_12633_, _04705_, _03705_);
  and (_12634_, _12633_, _03014_);
  and (_12635_, _12634_, _12632_);
  nor (_12636_, _05338_, _06814_);
  and (_12637_, _10620_, _05338_);
  or (_12638_, _12637_, _12636_);
  and (_12639_, _12638_, _02887_);
  and (_12640_, _10622_, _04705_);
  not (_12641_, _12640_);
  and (_12642_, _12641_, _12632_);
  or (_12643_, _12642_, _03821_);
  nand (_12644_, _04705_, _02618_);
  and (_12645_, _12644_, _12632_);
  and (_12647_, _12645_, _03825_);
  nor (_12648_, _03825_, _06814_);
  or (_12649_, _12648_, _02952_);
  or (_12650_, _12649_, _12647_);
  and (_12651_, _12650_, _02892_);
  and (_12652_, _12651_, _12643_);
  and (_12653_, _10617_, _05338_);
  or (_12654_, _12653_, _12636_);
  and (_12655_, _12654_, _02891_);
  or (_12656_, _12655_, _02947_);
  or (_12657_, _12656_, _12652_);
  nor (_12658_, _04705_, _06814_);
  and (_12659_, _04705_, _04005_);
  or (_12660_, _12659_, _12658_);
  or (_12661_, _12660_, _03327_);
  and (_12662_, _12661_, _12657_);
  or (_12663_, _12662_, _02950_);
  or (_12664_, _12645_, _02959_);
  and (_12665_, _12664_, _02888_);
  and (_12666_, _12665_, _12663_);
  or (_12667_, _12666_, _12639_);
  and (_12668_, _12667_, _02881_);
  or (_12669_, _12636_, _10616_);
  and (_12670_, _12669_, _02880_);
  and (_12671_, _12670_, _12654_);
  or (_12672_, _12671_, _06271_);
  or (_12673_, _12672_, _12668_);
  or (_12674_, _06698_, _06697_);
  nand (_12675_, _12674_, _06756_);
  or (_12676_, _12674_, _06756_);
  and (_12677_, _12676_, _12675_);
  or (_12678_, _12677_, _06277_);
  and (_12679_, _12678_, _02875_);
  and (_12680_, _12679_, _12673_);
  nor (_12681_, _10661_, _06794_);
  or (_12682_, _12681_, _12636_);
  and (_12683_, _12682_, _02874_);
  or (_12684_, _12683_, _06793_);
  or (_12685_, _12684_, _12680_);
  or (_12686_, _12660_, _06241_);
  and (_12687_, _12686_, _12685_);
  or (_12688_, _12687_, _02855_);
  and (_12689_, _06173_, _04705_);
  or (_12690_, _12658_, _02856_);
  or (_12691_, _12690_, _12689_);
  and (_12692_, _12691_, _02851_);
  and (_12693_, _12692_, _12688_);
  nand (_12694_, _10720_, _04705_);
  and (_12695_, _12632_, _02576_);
  and (_12696_, _12695_, _12694_);
  or (_12697_, _12696_, _06807_);
  or (_12698_, _12697_, _12693_);
  and (_12699_, _07164_, _07109_);
  nor (_12700_, _07159_, _07158_);
  or (_12701_, _12700_, _07160_);
  nor (_12702_, _12701_, _07164_);
  or (_12703_, _12702_, _12699_);
  or (_12704_, _12703_, _06813_);
  and (_12705_, _12704_, _03884_);
  and (_12706_, _12705_, _12698_);
  or (_12707_, _12706_, _12635_);
  and (_12708_, _12707_, _05279_);
  or (_12709_, _10612_, _06235_);
  and (_12710_, _12632_, _03021_);
  and (_12711_, _12710_, _12709_);
  or (_12712_, _12711_, _12708_);
  and (_12713_, _12712_, _03131_);
  or (_12714_, _10739_, _06235_);
  and (_12715_, _12632_, _03130_);
  and (_12716_, _12715_, _12714_);
  or (_12717_, _12716_, _12713_);
  and (_12718_, _12717_, _05274_);
  or (_12719_, _10611_, _06235_);
  and (_12720_, _12632_, _03020_);
  and (_12721_, _12720_, _12719_);
  or (_12722_, _12721_, _12718_);
  and (_12723_, _12722_, _03140_);
  not (_12724_, _05095_);
  or (_12725_, _12658_, _12724_);
  and (_12726_, _12645_, _03139_);
  and (_12727_, _12726_, _12725_);
  or (_12728_, _12727_, _12723_);
  and (_12729_, _12728_, _03128_);
  or (_12730_, _12644_, _12724_);
  and (_12731_, _12632_, _03127_);
  and (_12732_, _12731_, _12730_);
  or (_12733_, _12732_, _03166_);
  or (_12734_, _12633_, _12724_);
  and (_12735_, _12632_, _03036_);
  and (_12736_, _12735_, _12734_);
  or (_12737_, _12736_, _12733_);
  or (_12738_, _12737_, _12729_);
  or (_12739_, _12642_, _03563_);
  and (_12740_, _12739_, _02501_);
  and (_12741_, _12740_, _12738_);
  and (_12742_, _12638_, _02500_);
  or (_12743_, _12742_, _03174_);
  or (_12744_, _12743_, _12741_);
  or (_12745_, _12658_, _03178_);
  or (_12746_, _12745_, _12640_);
  and (_12747_, _12746_, _34698_);
  and (_12748_, _12747_, _12744_);
  or (_12749_, _12748_, _12631_);
  and (_35156_, _12749_, _36029_);
  nor (_12750_, _34698_, _06826_);
  nor (_12751_, _04705_, _06826_);
  and (_12752_, _10831_, _04705_);
  or (_12753_, _12752_, _12751_);
  and (_12754_, _12753_, _03130_);
  and (_12755_, _04705_, _05727_);
  or (_12756_, _12755_, _12751_);
  or (_12757_, _12756_, _03884_);
  nor (_12758_, _06235_, _04440_);
  or (_12759_, _12758_, _12751_);
  or (_12760_, _12759_, _06241_);
  and (_12761_, _10853_, _05338_);
  and (_12762_, _12761_, _10868_);
  nor (_12763_, _05338_, _06826_);
  or (_12764_, _12763_, _02881_);
  or (_12765_, _12764_, _12762_);
  or (_12766_, _12759_, _03327_);
  nor (_12767_, _10849_, _06235_);
  or (_12768_, _12767_, _12751_);
  or (_12769_, _12768_, _03821_);
  and (_12770_, _04705_, \oc8051_golden_model_1.ACC [2]);
  or (_12771_, _12770_, _12751_);
  and (_12772_, _12771_, _03825_);
  nor (_12773_, _03825_, _06826_);
  or (_12774_, _12773_, _02952_);
  or (_12775_, _12774_, _12772_);
  and (_12776_, _12775_, _02892_);
  and (_12777_, _12776_, _12769_);
  or (_12778_, _12763_, _12761_);
  and (_12779_, _12778_, _02891_);
  or (_12780_, _12779_, _02947_);
  or (_12781_, _12780_, _12777_);
  and (_12782_, _12781_, _12766_);
  or (_12783_, _12782_, _02950_);
  or (_12784_, _12771_, _02959_);
  and (_12785_, _12784_, _02888_);
  and (_12786_, _12785_, _12783_);
  and (_12787_, _10838_, _05338_);
  or (_12788_, _12787_, _12763_);
  and (_12789_, _12788_, _02887_);
  or (_12790_, _12789_, _02880_);
  or (_12791_, _12790_, _12786_);
  and (_12792_, _12791_, _12765_);
  or (_12793_, _12792_, _06271_);
  nor (_12794_, _06758_, _06654_);
  nor (_12795_, _12794_, _06759_);
  or (_12796_, _12795_, _06277_);
  and (_12797_, _12796_, _02875_);
  and (_12798_, _12797_, _12793_);
  nor (_12799_, _10886_, _06794_);
  or (_12800_, _12799_, _12763_);
  and (_12801_, _12800_, _02874_);
  or (_12802_, _12801_, _06793_);
  or (_12803_, _12802_, _12798_);
  and (_12804_, _12803_, _12760_);
  or (_12805_, _12804_, _02855_);
  and (_12806_, _06177_, _04705_);
  or (_12807_, _12751_, _02856_);
  or (_12808_, _12807_, _12806_);
  and (_12809_, _12808_, _12805_);
  or (_12810_, _12809_, _02576_);
  nor (_12811_, _10943_, _06235_);
  or (_12812_, _12751_, _02851_);
  or (_12813_, _12812_, _12811_);
  and (_12814_, _12813_, _06813_);
  and (_12815_, _12814_, _12810_);
  nand (_12816_, _07164_, _07099_);
  nor (_12817_, _07160_, _07110_);
  not (_12818_, _12817_);
  and (_12819_, _12818_, _07102_);
  nor (_12820_, _12818_, _07102_);
  nor (_12821_, _12820_, _12819_);
  or (_12822_, _12821_, _07164_);
  and (_12823_, _12822_, _06807_);
  and (_12824_, _12823_, _12816_);
  or (_12825_, _12824_, _03014_);
  or (_12826_, _12825_, _12815_);
  and (_12827_, _12826_, _12757_);
  or (_12828_, _12827_, _03021_);
  and (_12829_, _10835_, _04705_);
  or (_12830_, _12751_, _05279_);
  or (_12831_, _12830_, _12829_);
  and (_12832_, _12831_, _03131_);
  and (_12833_, _12832_, _12828_);
  or (_12834_, _12833_, _12754_);
  and (_12835_, _12834_, _05274_);
  or (_12836_, _12751_, _05143_);
  and (_12837_, _12756_, _03020_);
  and (_12838_, _12837_, _12836_);
  or (_12839_, _12838_, _12835_);
  and (_12840_, _12839_, _03140_);
  and (_12841_, _12771_, _03139_);
  and (_12842_, _12841_, _12836_);
  or (_12843_, _12842_, _03036_);
  or (_12844_, _12843_, _12840_);
  nor (_12845_, _10833_, _06235_);
  or (_12846_, _12751_, _05781_);
  or (_12847_, _12846_, _12845_);
  and (_12848_, _12847_, _05786_);
  and (_12849_, _12848_, _12844_);
  nor (_12850_, _10830_, _06235_);
  or (_12851_, _12850_, _12751_);
  and (_12852_, _12851_, _03127_);
  or (_12853_, _12852_, _03166_);
  or (_12854_, _12853_, _12849_);
  or (_12855_, _12768_, _03563_);
  and (_12856_, _12855_, _02501_);
  and (_12857_, _12856_, _12854_);
  and (_12858_, _12788_, _02500_);
  or (_12859_, _12858_, _03174_);
  or (_12860_, _12859_, _12857_);
  and (_12861_, _11008_, _04705_);
  or (_12862_, _12751_, _03178_);
  or (_12863_, _12862_, _12861_);
  and (_12864_, _12863_, _34698_);
  and (_12865_, _12864_, _12860_);
  or (_12866_, _12865_, _12750_);
  and (_35157_, _12866_, _36029_);
  nor (_12867_, _34698_, _06827_);
  nor (_12868_, _04705_, _06827_);
  and (_12869_, _11028_, _04705_);
  or (_12870_, _12869_, _12868_);
  and (_12871_, _12870_, _03130_);
  and (_12872_, _04705_, _05664_);
  or (_12873_, _12872_, _12868_);
  or (_12874_, _12873_, _03884_);
  nor (_12875_, _11143_, _06235_);
  or (_12876_, _12875_, _12868_);
  and (_12877_, _12876_, _02576_);
  nor (_12878_, _05338_, _06827_);
  and (_12879_, _11037_, _05338_);
  or (_12880_, _12879_, _12878_);
  or (_12881_, _12878_, _11066_);
  and (_12882_, _12881_, _12880_);
  or (_12883_, _12882_, _02881_);
  nor (_12884_, _11040_, _06235_);
  or (_12885_, _12884_, _12868_);
  or (_12886_, _12885_, _03821_);
  and (_12887_, _04705_, \oc8051_golden_model_1.ACC [3]);
  or (_12888_, _12887_, _12868_);
  and (_12889_, _12888_, _03825_);
  nor (_12890_, _03825_, _06827_);
  or (_12891_, _12890_, _02952_);
  or (_12892_, _12891_, _12889_);
  and (_12893_, _12892_, _02892_);
  and (_12894_, _12893_, _12886_);
  and (_12895_, _12880_, _02891_);
  or (_12896_, _12895_, _02947_);
  or (_12897_, _12896_, _12894_);
  nor (_12898_, _06235_, _04242_);
  or (_12899_, _12898_, _12868_);
  or (_12900_, _12899_, _03327_);
  and (_12901_, _12900_, _12897_);
  or (_12902_, _12901_, _02950_);
  or (_12903_, _12888_, _02959_);
  and (_12904_, _12903_, _02888_);
  and (_12905_, _12904_, _12902_);
  and (_12906_, _11035_, _05338_);
  or (_12907_, _12906_, _12878_);
  and (_12908_, _12907_, _02887_);
  or (_12909_, _12908_, _02880_);
  or (_12910_, _12909_, _12905_);
  and (_12911_, _12910_, _12883_);
  or (_12912_, _12911_, _06271_);
  nor (_12913_, _06761_, _06596_);
  nor (_12914_, _12913_, _06762_);
  or (_12915_, _12914_, _06277_);
  and (_12916_, _12915_, _02875_);
  and (_12917_, _12916_, _12912_);
  nor (_12918_, _11083_, _06794_);
  or (_12919_, _12918_, _12878_);
  and (_12920_, _12919_, _02874_);
  or (_12921_, _12920_, _06793_);
  or (_12922_, _12921_, _12917_);
  or (_12923_, _12899_, _06241_);
  and (_12924_, _12923_, _12922_);
  or (_12925_, _12924_, _02855_);
  and (_12926_, _06176_, _04705_);
  or (_12927_, _12868_, _02856_);
  or (_12928_, _12927_, _12926_);
  and (_12929_, _12928_, _02851_);
  and (_12930_, _12929_, _12925_);
  or (_12931_, _12930_, _12877_);
  and (_12932_, _12931_, _06813_);
  nand (_12933_, _07164_, _07090_);
  nor (_12934_, _12819_, _07101_);
  nor (_12935_, _12934_, _07093_);
  and (_12936_, _12934_, _07093_);
  or (_12937_, _12936_, _12935_);
  or (_12938_, _12937_, _07164_);
  and (_12939_, _12938_, _06807_);
  and (_12940_, _12939_, _12933_);
  or (_12941_, _12940_, _03014_);
  or (_12942_, _12941_, _12932_);
  and (_12943_, _12942_, _12874_);
  or (_12944_, _12943_, _03021_);
  and (_12945_, _11032_, _04705_);
  or (_12946_, _12868_, _05279_);
  or (_12947_, _12946_, _12945_);
  and (_12948_, _12947_, _03131_);
  and (_12949_, _12948_, _12944_);
  or (_12950_, _12949_, _12871_);
  and (_12951_, _12950_, _05274_);
  or (_12952_, _12868_, _04996_);
  and (_12953_, _12873_, _03020_);
  and (_12954_, _12953_, _12952_);
  or (_12955_, _12954_, _12951_);
  and (_12956_, _12955_, _03140_);
  and (_12957_, _12888_, _03139_);
  and (_12958_, _12957_, _12952_);
  or (_12959_, _12958_, _03036_);
  or (_12960_, _12959_, _12956_);
  nor (_12961_, _11030_, _06235_);
  or (_12962_, _12868_, _05781_);
  or (_12963_, _12962_, _12961_);
  and (_12964_, _12963_, _05786_);
  and (_12965_, _12964_, _12960_);
  nor (_12966_, _11027_, _06235_);
  or (_12967_, _12966_, _12868_);
  and (_12968_, _12967_, _03127_);
  or (_12969_, _12968_, _03166_);
  or (_12970_, _12969_, _12965_);
  or (_12971_, _12885_, _03563_);
  and (_12972_, _12971_, _02501_);
  and (_12973_, _12972_, _12970_);
  and (_12974_, _12907_, _02500_);
  or (_12975_, _12974_, _03174_);
  or (_12976_, _12975_, _12973_);
  and (_12977_, _11213_, _04705_);
  or (_12978_, _12868_, _03178_);
  or (_12979_, _12978_, _12977_);
  and (_12980_, _12979_, _34698_);
  and (_12981_, _12980_, _12976_);
  or (_12982_, _12981_, _12867_);
  and (_35159_, _12982_, _36029_);
  nor (_12983_, _34698_, _06951_);
  nor (_12984_, _04705_, _06951_);
  and (_12985_, _11368_, _04705_);
  or (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _03130_);
  and (_12988_, _05697_, _04705_);
  or (_12989_, _12988_, _12984_);
  or (_12990_, _12989_, _03884_);
  nor (_12991_, _11348_, _06235_);
  or (_12992_, _12991_, _12984_);
  and (_12993_, _12992_, _02576_);
  nor (_12994_, _05202_, _06235_);
  or (_12995_, _12994_, _12984_);
  or (_12996_, _12995_, _06241_);
  nor (_12997_, _05338_, _06951_);
  and (_12998_, _11243_, _05338_);
  or (_12999_, _12998_, _12997_);
  and (_13000_, _12999_, _02887_);
  nor (_13001_, _11259_, _06235_);
  or (_13002_, _13001_, _12984_);
  or (_13003_, _13002_, _03821_);
  and (_13004_, _04705_, \oc8051_golden_model_1.ACC [4]);
  or (_13005_, _13004_, _12984_);
  and (_13006_, _13005_, _03825_);
  nor (_13007_, _03825_, _06951_);
  or (_13008_, _13007_, _02952_);
  or (_13009_, _13008_, _13006_);
  and (_13010_, _13009_, _02892_);
  and (_13011_, _13010_, _13003_);
  and (_13012_, _11245_, _05338_);
  or (_13013_, _13012_, _12997_);
  and (_13014_, _13013_, _02891_);
  or (_13015_, _13014_, _02947_);
  or (_13016_, _13015_, _13011_);
  or (_13017_, _12995_, _03327_);
  and (_13018_, _13017_, _13016_);
  or (_13019_, _13018_, _02950_);
  or (_13020_, _13005_, _02959_);
  and (_13021_, _13020_, _02888_);
  and (_13022_, _13021_, _13019_);
  or (_13023_, _13022_, _13000_);
  and (_13024_, _13023_, _02881_);
  or (_13025_, _12997_, _11276_);
  and (_13026_, _13025_, _02880_);
  and (_13027_, _13026_, _13013_);
  or (_13028_, _13027_, _06271_);
  or (_13029_, _13028_, _13024_);
  nor (_13030_, _06766_, _06764_);
  nor (_13031_, _13030_, _06767_);
  or (_13032_, _13031_, _06277_);
  and (_13033_, _13032_, _02875_);
  and (_13034_, _13033_, _13029_);
  nor (_13035_, _11241_, _06794_);
  or (_13036_, _13035_, _12997_);
  and (_13037_, _13036_, _02874_);
  or (_13038_, _13037_, _06793_);
  or (_13039_, _13038_, _13034_);
  and (_13040_, _13039_, _12996_);
  or (_13041_, _13040_, _02855_);
  and (_13042_, _06181_, _04705_);
  or (_13043_, _12984_, _02856_);
  or (_13044_, _13043_, _13042_);
  and (_13045_, _13044_, _02851_);
  and (_13046_, _13045_, _13041_);
  or (_13047_, _13046_, _12993_);
  and (_13048_, _13047_, _06813_);
  nor (_13049_, _12934_, _07091_);
  or (_13050_, _13049_, _07092_);
  nand (_13051_, _13050_, _07133_);
  or (_13052_, _13050_, _07133_);
  and (_13053_, _13052_, _13051_);
  or (_13054_, _13053_, _07164_);
  nand (_13055_, _07164_, _07130_);
  and (_13056_, _13055_, _06807_);
  and (_13057_, _13056_, _13054_);
  or (_13058_, _13057_, _03014_);
  or (_13059_, _13058_, _13048_);
  and (_13060_, _13059_, _12990_);
  or (_13061_, _13060_, _03021_);
  and (_13062_, _11362_, _04705_);
  or (_13063_, _12984_, _05279_);
  or (_13064_, _13063_, _13062_);
  and (_13065_, _13064_, _03131_);
  and (_13066_, _13065_, _13061_);
  or (_13067_, _13066_, _12987_);
  and (_13068_, _13067_, _05274_);
  or (_13069_, _12984_, _05251_);
  and (_13070_, _12989_, _03020_);
  and (_13071_, _13070_, _13069_);
  or (_13072_, _13071_, _13068_);
  and (_13073_, _13072_, _03140_);
  and (_13074_, _13005_, _03139_);
  and (_13075_, _13074_, _13069_);
  or (_13076_, _13075_, _03036_);
  or (_13077_, _13076_, _13073_);
  nor (_13078_, _11361_, _06235_);
  or (_13079_, _12984_, _05781_);
  or (_13080_, _13079_, _13078_);
  and (_13081_, _13080_, _05786_);
  and (_13082_, _13081_, _13077_);
  nor (_13083_, _11367_, _06235_);
  or (_13084_, _13083_, _12984_);
  and (_13085_, _13084_, _03127_);
  or (_13086_, _13085_, _03166_);
  or (_13087_, _13086_, _13082_);
  or (_13088_, _13002_, _03563_);
  and (_13089_, _13088_, _02501_);
  and (_13090_, _13089_, _13087_);
  and (_13091_, _12999_, _02500_);
  or (_13092_, _13091_, _03174_);
  or (_13093_, _13092_, _13090_);
  and (_13094_, _11417_, _04705_);
  or (_13095_, _12984_, _03178_);
  or (_13096_, _13095_, _13094_);
  and (_13097_, _13096_, _34698_);
  and (_13098_, _13097_, _13093_);
  or (_13099_, _13098_, _12983_);
  and (_35160_, _13099_, _36029_);
  nor (_13100_, _34698_, _06942_);
  nor (_13101_, _04705_, _06942_);
  and (_13102_, _11436_, _04705_);
  or (_13103_, _13102_, _13101_);
  and (_13104_, _13103_, _03130_);
  and (_13105_, _05701_, _04705_);
  or (_13106_, _13105_, _13101_);
  or (_13107_, _13106_, _03884_);
  nor (_13108_, _11546_, _06235_);
  or (_13109_, _13108_, _13101_);
  and (_13110_, _13109_, _02576_);
  nor (_13111_, _04896_, _06235_);
  or (_13112_, _13111_, _13101_);
  or (_13113_, _13112_, _06241_);
  nor (_13114_, _05338_, _06942_);
  and (_13115_, _11442_, _05338_);
  or (_13116_, _13115_, _13114_);
  and (_13117_, _13116_, _02887_);
  nor (_13118_, _11445_, _06235_);
  or (_13119_, _13118_, _13101_);
  or (_13120_, _13119_, _03821_);
  and (_13121_, _04705_, \oc8051_golden_model_1.ACC [5]);
  or (_13122_, _13121_, _13101_);
  and (_13123_, _13122_, _03825_);
  nor (_13124_, _03825_, _06942_);
  or (_13125_, _13124_, _02952_);
  or (_13126_, _13125_, _13123_);
  and (_13127_, _13126_, _02892_);
  and (_13128_, _13127_, _13120_);
  and (_13129_, _11459_, _05338_);
  or (_13130_, _13129_, _13114_);
  and (_13131_, _13130_, _02891_);
  or (_13132_, _13131_, _02947_);
  or (_13133_, _13132_, _13128_);
  or (_13134_, _13112_, _03327_);
  and (_13135_, _13134_, _13133_);
  or (_13136_, _13135_, _02950_);
  or (_13137_, _13122_, _02959_);
  and (_13138_, _13137_, _02888_);
  and (_13139_, _13138_, _13136_);
  or (_13140_, _13139_, _13117_);
  and (_13141_, _13140_, _02881_);
  or (_13142_, _13114_, _11474_);
  and (_13143_, _13130_, _02880_);
  and (_13144_, _13143_, _13142_);
  or (_13145_, _13144_, _06271_);
  or (_13146_, _13145_, _13141_);
  nor (_13147_, _06769_, _06470_);
  nor (_13148_, _13147_, _06770_);
  or (_13149_, _13148_, _06277_);
  and (_13150_, _13149_, _02875_);
  and (_13151_, _13150_, _13146_);
  nor (_13152_, _11440_, _06794_);
  or (_13153_, _13152_, _13114_);
  and (_13154_, _13153_, _02874_);
  or (_13155_, _13154_, _06793_);
  or (_13156_, _13155_, _13151_);
  and (_13157_, _13156_, _13113_);
  or (_13158_, _13157_, _02855_);
  and (_13159_, _06180_, _04705_);
  or (_13160_, _13101_, _02856_);
  or (_13161_, _13160_, _13159_);
  and (_13162_, _13161_, _02851_);
  and (_13163_, _13162_, _13158_);
  or (_13164_, _13163_, _13110_);
  and (_13165_, _13164_, _06813_);
  nand (_13166_, _07164_, _07141_);
  not (_13167_, _07132_);
  and (_13168_, _13051_, _13167_);
  nor (_13169_, _13168_, _07144_);
  and (_13170_, _13168_, _07144_);
  or (_13171_, _13170_, _13169_);
  or (_13172_, _13171_, _07164_);
  and (_13173_, _13172_, _06807_);
  and (_13174_, _13173_, _13166_);
  or (_13175_, _13174_, _03014_);
  or (_13176_, _13175_, _13165_);
  and (_13177_, _13176_, _13107_);
  or (_13178_, _13177_, _03021_);
  and (_13179_, _11562_, _04705_);
  or (_13180_, _13101_, _05279_);
  or (_13181_, _13180_, _13179_);
  and (_13182_, _13181_, _03131_);
  and (_13183_, _13182_, _13178_);
  or (_13184_, _13183_, _13104_);
  and (_13185_, _13184_, _05274_);
  or (_13186_, _13101_, _04944_);
  and (_13187_, _13106_, _03020_);
  and (_13188_, _13187_, _13186_);
  or (_13189_, _13188_, _13185_);
  and (_13190_, _13189_, _03140_);
  and (_13191_, _13122_, _03139_);
  and (_13192_, _13191_, _13186_);
  or (_13193_, _13192_, _03036_);
  or (_13194_, _13193_, _13190_);
  nor (_13195_, _11560_, _06235_);
  or (_13196_, _13101_, _05781_);
  or (_13197_, _13196_, _13195_);
  and (_13198_, _13197_, _05786_);
  and (_13199_, _13198_, _13194_);
  nor (_13200_, _11435_, _06235_);
  or (_13201_, _13200_, _13101_);
  and (_13202_, _13201_, _03127_);
  or (_13203_, _13202_, _03166_);
  or (_13204_, _13203_, _13199_);
  or (_13205_, _13119_, _03563_);
  and (_13206_, _13205_, _02501_);
  and (_13207_, _13206_, _13204_);
  and (_13208_, _13116_, _02500_);
  or (_13209_, _13208_, _03174_);
  or (_13210_, _13209_, _13207_);
  and (_13211_, _11619_, _04705_);
  or (_13212_, _13101_, _03178_);
  or (_13213_, _13212_, _13211_);
  and (_13214_, _13213_, _34698_);
  and (_13215_, _13214_, _13210_);
  or (_13216_, _13215_, _13100_);
  and (_35161_, _13216_, _36029_);
  nor (_13217_, _34698_, _07066_);
  nor (_13218_, _04705_, _07066_);
  and (_13219_, _11769_, _04705_);
  or (_13220_, _13219_, _13218_);
  and (_13221_, _13220_, _03130_);
  and (_13222_, _11758_, _04705_);
  or (_13223_, _13222_, _13218_);
  or (_13224_, _13223_, _03884_);
  nor (_13225_, _11751_, _06235_);
  or (_13226_, _13225_, _13218_);
  and (_13227_, _13226_, _02576_);
  nor (_13228_, _04787_, _06235_);
  or (_13229_, _13228_, _13218_);
  or (_13230_, _13229_, _06241_);
  nor (_13231_, _05338_, _07066_);
  and (_13232_, _11675_, _05338_);
  or (_13233_, _13232_, _13231_);
  and (_13234_, _13233_, _02887_);
  nor (_13235_, _11636_, _06235_);
  or (_13236_, _13235_, _13218_);
  or (_13237_, _13236_, _03821_);
  and (_13238_, _04705_, \oc8051_golden_model_1.ACC [6]);
  or (_13239_, _13238_, _13218_);
  and (_13240_, _13239_, _03825_);
  nor (_13241_, _03825_, _07066_);
  or (_13242_, _13241_, _02952_);
  or (_13243_, _13242_, _13240_);
  and (_13244_, _13243_, _02892_);
  and (_13245_, _13244_, _13237_);
  and (_13246_, _11653_, _05338_);
  or (_13247_, _13246_, _13231_);
  and (_13248_, _13247_, _02891_);
  or (_13249_, _13248_, _02947_);
  or (_13250_, _13249_, _13245_);
  or (_13251_, _13229_, _03327_);
  and (_13252_, _13251_, _13250_);
  or (_13253_, _13252_, _02950_);
  or (_13254_, _13239_, _02959_);
  and (_13255_, _13254_, _02888_);
  and (_13256_, _13255_, _13253_);
  or (_13257_, _13256_, _13234_);
  and (_13258_, _13257_, _02881_);
  or (_13259_, _13231_, _11682_);
  and (_13260_, _13247_, _02880_);
  and (_13261_, _13260_, _13259_);
  or (_13262_, _13261_, _06271_);
  or (_13263_, _13262_, _13258_);
  nor (_13264_, _06785_, _06772_);
  nor (_13265_, _13264_, _06786_);
  or (_13266_, _13265_, _06277_);
  and (_13267_, _13266_, _02875_);
  and (_13268_, _13267_, _13263_);
  nor (_13269_, _11650_, _06794_);
  or (_13270_, _13269_, _13231_);
  and (_13271_, _13270_, _02874_);
  or (_13272_, _13271_, _06793_);
  or (_13273_, _13272_, _13268_);
  and (_13274_, _13273_, _13230_);
  or (_13275_, _13274_, _02855_);
  and (_13276_, _05847_, _04705_);
  or (_13277_, _13218_, _02856_);
  or (_13278_, _13277_, _13276_);
  and (_13279_, _13278_, _02851_);
  and (_13280_, _13279_, _13275_);
  or (_13281_, _13280_, _13227_);
  and (_13282_, _13281_, _06813_);
  nor (_13283_, _13168_, _07142_);
  or (_13284_, _13283_, _07143_);
  and (_13285_, _13284_, _07123_);
  nor (_13286_, _13284_, _07123_);
  or (_13287_, _13286_, _13285_);
  or (_13288_, _13287_, _07164_);
  nand (_13289_, _07164_, _07079_);
  and (_13290_, _13289_, _06807_);
  and (_13291_, _13290_, _13288_);
  or (_13292_, _13291_, _03014_);
  or (_13293_, _13292_, _13282_);
  and (_13294_, _13293_, _13224_);
  or (_13295_, _13294_, _03021_);
  and (_13296_, _11646_, _04705_);
  or (_13297_, _13218_, _05279_);
  or (_13298_, _13297_, _13296_);
  and (_13299_, _13298_, _03131_);
  and (_13300_, _13299_, _13295_);
  or (_13301_, _13300_, _13221_);
  and (_13302_, _13301_, _05274_);
  or (_13303_, _13218_, _04838_);
  and (_13304_, _13223_, _03020_);
  and (_13305_, _13304_, _13303_);
  or (_13306_, _13305_, _13302_);
  and (_13307_, _13306_, _03140_);
  and (_13308_, _13239_, _03139_);
  and (_13309_, _13308_, _13303_);
  or (_13310_, _13309_, _03036_);
  or (_13311_, _13310_, _13307_);
  nor (_13312_, _11644_, _06235_);
  or (_13313_, _13218_, _05781_);
  or (_13314_, _13313_, _13312_);
  and (_13315_, _13314_, _05786_);
  and (_13316_, _13315_, _13311_);
  nor (_13317_, _11768_, _06235_);
  or (_13318_, _13317_, _13218_);
  and (_13319_, _13318_, _03127_);
  or (_13320_, _13319_, _03166_);
  or (_13321_, _13320_, _13316_);
  or (_13322_, _13236_, _03563_);
  and (_13323_, _13322_, _02501_);
  and (_13324_, _13323_, _13321_);
  and (_13325_, _13233_, _02500_);
  or (_13326_, _13325_, _03174_);
  or (_13327_, _13326_, _13324_);
  and (_13328_, _11821_, _04705_);
  or (_13329_, _13218_, _03178_);
  or (_13330_, _13329_, _13328_);
  and (_13331_, _13330_, _34698_);
  and (_13332_, _13331_, _13327_);
  or (_13333_, _13332_, _13217_);
  and (_35162_, _13333_, _36029_);
  nor (_13334_, _34698_, _02549_);
  and (_13335_, _08184_, \oc8051_golden_model_1.ACC [1]);
  nand (_13336_, _08135_, _05768_);
  nand (_13337_, _07734_, _02899_);
  and (_13338_, _13337_, _08106_);
  and (_13339_, _05938_, _02549_);
  nor (_13340_, _08084_, _13339_);
  and (_13341_, _07217_, _02545_);
  nand (_13342_, _13341_, _13340_);
  nor (_13343_, _08008_, _02549_);
  nor (_13344_, _13343_, _10088_);
  nand (_13345_, _13344_, _03137_);
  and (_13346_, _13345_, _08031_);
  nand (_13347_, _07865_, _09316_);
  not (_13348_, _02537_);
  nor (_13349_, _02976_, _13348_);
  nor (_13350_, _04712_, _02549_);
  and (_13351_, _04712_, _03817_);
  nor (_13352_, _13351_, _13350_);
  nand (_13353_, _13352_, _06793_);
  and (_13354_, _07327_, _02549_);
  or (_13355_, _13354_, _08039_);
  nand (_13356_, _13355_, _07276_);
  or (_13357_, _07430_, _03817_);
  nor (_13358_, _03818_, _07435_);
  or (_13359_, _13358_, _06174_);
  or (_13360_, _07440_, _03817_);
  nor (_13361_, _07442_, \oc8051_golden_model_1.ACC [0]);
  and (_13362_, _07442_, \oc8051_golden_model_1.ACC [0]);
  or (_13363_, _13362_, _13361_);
  nand (_13364_, _13363_, _09203_);
  and (_13365_, _13364_, _13360_);
  or (_13366_, _13365_, _02954_);
  nand (_13367_, _07700_, _02954_);
  and (_13368_, _13367_, _09202_);
  and (_13369_, _13368_, _13366_);
  or (_13370_, _13369_, _03818_);
  and (_13371_, _13370_, _03821_);
  and (_13372_, _13371_, _13359_);
  and (_13373_, _05044_, _04712_);
  nor (_13374_, _13373_, _13350_);
  nor (_13375_, _13374_, _03821_);
  or (_13376_, _13375_, _02891_);
  or (_13377_, _13376_, _13372_);
  nor (_13378_, _05331_, _02549_);
  and (_13379_, _10429_, _05331_);
  nor (_13380_, _13379_, _13378_);
  nand (_13381_, _13380_, _02891_);
  and (_13382_, _13381_, _03327_);
  and (_13383_, _13382_, _13377_);
  nor (_13384_, _13352_, _03327_);
  or (_13385_, _13384_, _07431_);
  or (_13386_, _13385_, _13383_);
  and (_13387_, _13386_, _13357_);
  or (_13388_, _13387_, _03413_);
  or (_13389_, _06174_, _03849_);
  and (_13390_, _13389_, _02959_);
  and (_13391_, _13390_, _13388_);
  nor (_13392_, _07700_, _02959_);
  or (_13393_, _13392_, _07497_);
  or (_13394_, _13393_, _13391_);
  nand (_13395_, _07497_, _06885_);
  and (_13396_, _13395_, _13394_);
  or (_13397_, _13396_, _02887_);
  or (_13398_, _13350_, _02888_);
  and (_13399_, _13398_, _02881_);
  and (_13400_, _13399_, _13397_);
  nor (_13401_, _13374_, _02881_);
  or (_13402_, _13401_, _06271_);
  or (_13403_, _13402_, _13400_);
  not (_13404_, _06732_);
  nand (_13405_, _13404_, _06271_);
  and (_13406_, _13405_, _07426_);
  and (_13407_, _13406_, _13403_);
  nor (_13408_, _07577_, _07426_);
  or (_13409_, _13408_, _03441_);
  or (_13410_, _13409_, _13407_);
  nand (_13411_, _07407_, _03441_);
  and (_13412_, _13411_, _02997_);
  and (_13413_, _13412_, _13410_);
  nand (_13414_, _13344_, _07277_);
  and (_13415_, _13414_, _07597_);
  or (_13416_, _13415_, _13413_);
  and (_13417_, _13416_, _13356_);
  or (_13418_, _13417_, _02585_);
  nand (_13419_, _02832_, _02585_);
  and (_13420_, _13419_, _02875_);
  and (_13421_, _13420_, _13418_);
  nor (_13422_, _10473_, _07755_);
  nor (_13423_, _13422_, _13378_);
  nor (_13424_, _13423_, _02875_);
  or (_13425_, _13424_, _06793_);
  or (_13426_, _13425_, _13421_);
  and (_13427_, _13426_, _13353_);
  or (_13428_, _13427_, _02855_);
  and (_13429_, _06174_, _04712_);
  nor (_13430_, _13429_, _13350_);
  nand (_13431_, _13430_, _02855_);
  and (_13432_, _13431_, _02851_);
  and (_13433_, _13432_, _13428_);
  nor (_13434_, _10530_, _07272_);
  nor (_13435_, _13434_, _13350_);
  nor (_13436_, _13435_, _02851_);
  or (_13437_, _13436_, _06807_);
  or (_13438_, _13437_, _13433_);
  nand (_13439_, _07164_, _06807_);
  and (_13440_, _13439_, _13438_);
  and (_13441_, _13440_, _02584_);
  nor (_13442_, _02832_, _02584_);
  or (_13443_, _13442_, _03014_);
  or (_13444_, _13443_, _13441_);
  and (_13445_, _04712_, _05566_);
  nor (_13446_, _13445_, _13350_);
  nand (_13447_, _13446_, _03014_);
  and (_13448_, _13447_, _07783_);
  and (_13449_, _13448_, _13444_);
  nor (_13450_, _07783_, _02832_);
  or (_13451_, _13450_, _07799_);
  or (_13452_, _13451_, _13449_);
  nor (_13453_, _03817_, \oc8051_golden_model_1.ACC [0]);
  nor (_13454_, _13453_, _07242_);
  or (_13455_, _07798_, _13454_);
  and (_13456_, _13455_, _07803_);
  and (_13457_, _13456_, _13452_);
  and (_13458_, _13340_, _07802_);
  or (_13459_, _13458_, _03132_);
  or (_13460_, _13459_, _13457_);
  or (_13461_, _10546_, _07814_);
  and (_13462_, _13461_, _13460_);
  or (_13463_, _13462_, _07812_);
  or (_13464_, _07813_, _09317_);
  and (_13465_, _13464_, _13463_);
  or (_13466_, _13465_, _03021_);
  and (_13467_, _10425_, _04712_);
  nor (_13468_, _13467_, _13350_);
  nand (_13469_, _13468_, _03021_);
  and (_13470_, _13469_, _03131_);
  and (_13471_, _13470_, _13466_);
  and (_13472_, _13350_, _03130_);
  or (_13473_, _13472_, _13471_);
  and (_13474_, _13473_, _07828_);
  and (_13475_, _07827_, _07242_);
  or (_13476_, _13475_, _13474_);
  and (_13477_, _13476_, _07265_);
  and (_13478_, _08084_, _03513_);
  or (_13479_, _13478_, _03141_);
  or (_13480_, _13479_, _13477_);
  or (_13481_, _10545_, _07838_);
  and (_13482_, _13481_, _07837_);
  and (_13483_, _13482_, _13480_);
  and (_13484_, _07836_, _08157_);
  or (_13485_, _13484_, _13483_);
  and (_13486_, _13485_, _05274_);
  and (_13487_, _03360_, _10788_);
  nor (_13488_, _13446_, _13373_);
  and (_13489_, _13488_, _03020_);
  or (_13490_, _13489_, _13487_);
  or (_13491_, _13490_, _13486_);
  nand (_13492_, _13487_, _13453_);
  nand (_13493_, _13492_, _13491_);
  nor (_13494_, _13493_, _13349_);
  not (_13495_, _13453_);
  and (_13496_, _13349_, _13495_);
  or (_13497_, _13496_, _07852_);
  or (_13498_, _13497_, _13494_);
  nand (_13499_, _07852_, _13453_);
  and (_13500_, _13499_, _07854_);
  and (_13501_, _13500_, _13498_);
  nor (_13502_, _13453_, _07854_);
  or (_13503_, _13502_, _07858_);
  or (_13504_, _13503_, _13501_);
  nand (_13505_, _13339_, _07858_);
  and (_13506_, _13505_, _03126_);
  and (_13507_, _13506_, _13504_);
  nand (_13508_, _10421_, _07868_);
  and (_13509_, _13508_, _07867_);
  or (_13510_, _13509_, _13507_);
  and (_13511_, _13510_, _13347_);
  or (_13512_, _13511_, _03036_);
  nor (_13513_, _10423_, _07272_);
  nor (_13514_, _13513_, _13350_);
  nand (_13515_, _13514_, _03036_);
  not (_13516_, _07887_);
  nand (_13517_, _13516_, _07882_);
  not (_13518_, _13517_);
  and (_13519_, _13518_, _13515_);
  and (_13520_, _13519_, _13512_);
  nor (_13521_, _13518_, _07577_);
  or (_13522_, _13521_, _07886_);
  or (_13523_, _13522_, _13520_);
  nand (_13524_, _07577_, _07886_);
  and (_13525_, _13524_, _07922_);
  and (_13526_, _13525_, _13523_);
  nor (_13527_, _07407_, _07922_);
  or (_13528_, _13527_, _03137_);
  or (_13529_, _13528_, _13526_);
  and (_13530_, _13529_, _13346_);
  nor (_13531_, _08031_, _13355_);
  or (_13532_, _13531_, _08029_);
  nor (_13533_, _13532_, _13530_);
  and (_13534_, _08029_, _07319_);
  or (_13535_, _13534_, _07258_);
  or (_13536_, _13535_, _13533_);
  nand (_13537_, _13454_, _07258_);
  and (_13538_, _13537_, _13536_);
  or (_13539_, _13538_, _07217_);
  nand (_13540_, _13539_, _13342_);
  and (_13541_, _03388_, _02535_);
  nand (_13542_, _13340_, _13541_);
  nand (_13543_, _13542_, _02901_);
  or (_13544_, _13543_, _13540_);
  and (_13545_, _13544_, _13338_);
  and (_13546_, _08103_, _09317_);
  or (_13547_, _13546_, _08135_);
  or (_13548_, _13547_, _13545_);
  and (_13549_, _13548_, _13336_);
  or (_13550_, _13549_, _03166_);
  nand (_13551_, _13374_, _03166_);
  and (_13552_, _13551_, _08180_);
  and (_13553_, _13552_, _13550_);
  and (_13554_, _08179_, _02549_);
  or (_13555_, _13554_, _13553_);
  and (_13556_, _13555_, _09787_);
  or (_13557_, _13556_, _13335_);
  and (_13558_, _13557_, _02501_);
  and (_13559_, _13350_, _02500_);
  or (_13560_, _13559_, _03174_);
  or (_13562_, _13560_, _13558_);
  nand (_13563_, _13374_, _03174_);
  and (_13564_, _13563_, _08202_);
  and (_13565_, _13564_, _13562_);
  and (_13566_, _08201_, _02549_);
  or (_13567_, _13566_, _08208_);
  or (_13568_, _13567_, _13565_);
  nand (_13569_, _08208_, _02618_);
  and (_13570_, _13569_, _34698_);
  and (_13571_, _13570_, _13568_);
  or (_13573_, _13571_, _13334_);
  and (_35164_, _13573_, _36029_);
  nor (_13574_, _34698_, _02618_);
  nand (_13575_, _08135_, _02549_);
  and (_13576_, _07931_, _07405_);
  nor (_13577_, _13576_, _07932_);
  or (_13578_, _13577_, _07922_);
  nand (_13579_, _07865_, _08155_);
  or (_13580_, _08081_, _07265_);
  not (_13581_, _09468_);
  nor (_13583_, _04712_, _02618_);
  and (_13584_, _13583_, _03130_);
  and (_13585_, _04712_, _04005_);
  nor (_13586_, _13585_, _13583_);
  nand (_13587_, _13586_, _06793_);
  and (_13588_, \oc8051_golden_model_1.PSW [7], _02549_);
  and (_13589_, _07319_, \oc8051_golden_model_1.ACC [0]);
  nor (_13590_, _13589_, _02832_);
  nor (_13591_, _13590_, _13588_);
  and (_13592_, _13591_, _08156_);
  nor (_13594_, _13591_, _08156_);
  nor (_13595_, _13594_, _13592_);
  nand (_13596_, _13595_, _07276_);
  or (_13597_, _07430_, _04005_);
  or (_13598_, _07440_, _04005_);
  or (_13599_, _07442_, _02618_);
  nand (_13600_, _07442_, _02618_);
  and (_13601_, _13600_, _13599_);
  nand (_13602_, _13601_, _09203_);
  and (_13603_, _13602_, _13598_);
  or (_13605_, _13603_, _02954_);
  nand (_13606_, _07681_, _02954_);
  and (_13607_, _13606_, _09202_);
  and (_13608_, _13607_, _13605_);
  or (_13609_, _13608_, _03818_);
  or (_13610_, _13358_, _06173_);
  and (_13611_, _13610_, _13609_);
  and (_13612_, _13611_, _03821_);
  nor (_13613_, _04712_, \oc8051_golden_model_1.ACC [1]);
  and (_13614_, _10622_, _04712_);
  nor (_13616_, _13614_, _13613_);
  and (_13617_, _13616_, _02952_);
  or (_13618_, _13617_, _07455_);
  or (_13619_, _13618_, _13612_);
  nor (_13620_, _07462_, \oc8051_golden_model_1.PSW [6]);
  nor (_13621_, _13620_, \oc8051_golden_model_1.ACC [1]);
  and (_13622_, _13620_, \oc8051_golden_model_1.ACC [1]);
  nor (_13623_, _13622_, _13621_);
  nand (_13624_, _13623_, _07455_);
  and (_13625_, _13624_, _02951_);
  and (_13627_, _13625_, _13619_);
  nor (_13628_, _05331_, _02618_);
  and (_13629_, _10617_, _05331_);
  nor (_13630_, _13629_, _13628_);
  nor (_13631_, _13630_, _02892_);
  nor (_13632_, _13586_, _03327_);
  or (_13633_, _13632_, _07431_);
  or (_13634_, _13633_, _13631_);
  or (_13635_, _13634_, _13627_);
  and (_13636_, _13635_, _13597_);
  or (_13638_, _13636_, _03413_);
  or (_13639_, _06173_, _03849_);
  and (_13640_, _13639_, _02959_);
  and (_13641_, _13640_, _13638_);
  nor (_13642_, _07681_, _02959_);
  or (_13643_, _13642_, _07497_);
  or (_13644_, _13643_, _13641_);
  nand (_13645_, _07497_, _06879_);
  and (_13646_, _13645_, _13644_);
  or (_13647_, _13646_, _02887_);
  and (_13649_, _10620_, _05331_);
  nor (_13650_, _13649_, _13628_);
  nand (_13651_, _13650_, _02887_);
  and (_13652_, _13651_, _02881_);
  and (_13653_, _13652_, _13647_);
  and (_13654_, _13629_, _10616_);
  nor (_13655_, _13654_, _13628_);
  nor (_13656_, _13655_, _02881_);
  or (_13657_, _13656_, _06271_);
  or (_13658_, _13657_, _13653_);
  and (_13660_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_13661_, _13660_, _07105_);
  nor (_13662_, _13661_, _06733_);
  or (_13663_, _13662_, _06277_);
  and (_13664_, _13663_, _07426_);
  and (_13665_, _13664_, _13658_);
  not (_13666_, _09005_);
  not (_13667_, _13589_);
  and (_13668_, _13667_, _03817_);
  nor (_13669_, _13668_, _13588_);
  and (_13671_, _13669_, _07241_);
  nor (_13672_, _13669_, _07241_);
  or (_13673_, _13672_, _13671_);
  or (_13674_, _13673_, _03441_);
  and (_13675_, _13674_, _13666_);
  or (_13676_, _13675_, _13665_);
  and (_13677_, _13667_, _06174_);
  nor (_13678_, _13677_, _13588_);
  and (_13679_, _13678_, _08083_);
  nor (_13680_, _13678_, _08083_);
  or (_13682_, _13680_, _13679_);
  or (_13683_, _13682_, _07344_);
  and (_13684_, _13683_, _02997_);
  and (_13685_, _13684_, _13676_);
  nor (_13686_, _07700_, _13589_);
  nor (_13687_, _13686_, _13588_);
  and (_13688_, _13687_, _07732_);
  nor (_13689_, _13687_, _07732_);
  or (_13690_, _13689_, _13688_);
  nand (_13691_, _13690_, _07277_);
  and (_13693_, _13691_, _07597_);
  or (_13694_, _13693_, _13685_);
  and (_13695_, _13694_, _13596_);
  or (_13696_, _13695_, _02585_);
  nand (_13697_, _03671_, _02585_);
  and (_13698_, _13697_, _02875_);
  and (_13699_, _13698_, _13696_);
  nor (_13700_, _10661_, _07755_);
  nor (_13701_, _13700_, _13628_);
  nor (_13702_, _13701_, _02875_);
  or (_13704_, _13702_, _06793_);
  or (_13705_, _13704_, _13699_);
  and (_13706_, _13705_, _13587_);
  or (_13707_, _13706_, _02855_);
  and (_13708_, _06173_, _04712_);
  nor (_13709_, _13708_, _13583_);
  nand (_13710_, _13709_, _02855_);
  and (_13711_, _13710_, _02851_);
  and (_13712_, _13711_, _13707_);
  nor (_13713_, _10720_, _07272_);
  nor (_13714_, _13713_, _13583_);
  nor (_13715_, _13714_, _02851_);
  or (_13716_, _13715_, _06807_);
  or (_13717_, _13716_, _13712_);
  or (_13718_, _07069_, _06813_);
  and (_13719_, _13718_, _13717_);
  and (_13720_, _13719_, _02584_);
  nor (_13721_, _03671_, _02584_);
  or (_13722_, _13721_, _03014_);
  or (_13723_, _13722_, _13720_);
  and (_13724_, _04712_, _03705_);
  nor (_13725_, _13724_, _13613_);
  or (_13726_, _13725_, _03884_);
  and (_13727_, _13726_, _07783_);
  and (_13728_, _13727_, _13723_);
  nor (_13729_, _07783_, _03671_);
  or (_13730_, _13729_, _07791_);
  or (_13731_, _13730_, _13728_);
  not (_13732_, _07793_);
  or (_13733_, _07792_, _07241_);
  and (_13734_, _13733_, _13732_);
  and (_13735_, _13734_, _13731_);
  and (_13736_, _07793_, _07241_);
  or (_13737_, _13736_, _07796_);
  or (_13738_, _13737_, _13735_);
  not (_13739_, _07796_);
  or (_13740_, _13739_, _07241_);
  and (_13741_, _13740_, _07803_);
  and (_13742_, _13741_, _13738_);
  and (_13743_, _08083_, _07802_);
  or (_13744_, _13743_, _03132_);
  or (_13745_, _13744_, _13742_);
  or (_13746_, _10739_, _07814_);
  and (_13747_, _13746_, _07813_);
  and (_13748_, _13747_, _13745_);
  and (_13749_, _07812_, _08156_);
  or (_13750_, _13749_, _03021_);
  or (_13751_, _13750_, _13748_);
  and (_13752_, _10612_, _04712_);
  nor (_13753_, _13752_, _13583_);
  nand (_13754_, _13753_, _03021_);
  and (_13755_, _13754_, _03131_);
  and (_13756_, _13755_, _13751_);
  or (_13757_, _13756_, _13584_);
  and (_13758_, _13757_, _13581_);
  and (_13759_, _09468_, _07239_);
  or (_13760_, _13759_, _09467_);
  or (_13761_, _13760_, _13758_);
  not (_13762_, _09467_);
  or (_13763_, _13762_, _07239_);
  and (_13764_, _13763_, _09471_);
  and (_13765_, _13764_, _13761_);
  not (_13766_, _07239_);
  nor (_13767_, _09471_, _13766_);
  or (_13768_, _13767_, _03513_);
  or (_13769_, _13768_, _13765_);
  and (_13770_, _13769_, _13580_);
  or (_13771_, _13770_, _03141_);
  or (_13772_, _10737_, _07838_);
  and (_13773_, _13772_, _07837_);
  and (_13774_, _13773_, _13771_);
  and (_13775_, _07836_, _08154_);
  or (_13776_, _13775_, _13774_);
  and (_13777_, _13776_, _05274_);
  and (_13778_, _10611_, _04712_);
  nor (_13779_, _13778_, _13583_);
  nor (_13780_, _13779_, _05274_);
  or (_13781_, _13780_, _09487_);
  or (_13782_, _13781_, _13777_);
  nand (_13783_, _08082_, _07858_);
  not (_13784_, _08872_);
  nand (_13785_, _13784_, _07240_);
  and (_13786_, _13785_, _03126_);
  and (_13787_, _13786_, _13783_);
  and (_13788_, _13787_, _13782_);
  nand (_13789_, _10738_, _07868_);
  and (_13790_, _13789_, _07867_);
  or (_13791_, _13790_, _13788_);
  and (_13792_, _13791_, _13579_);
  or (_13793_, _13792_, _03036_);
  nor (_13794_, _10610_, _07272_);
  or (_13795_, _13794_, _13583_);
  or (_13796_, _13795_, _05781_);
  and (_13797_, _13796_, _07889_);
  and (_13798_, _13797_, _13793_);
  and (_13799_, _07898_, _07575_);
  nor (_13800_, _13799_, _07899_);
  and (_13801_, _13800_, _10171_);
  or (_13802_, _13801_, _07917_);
  or (_13803_, _13802_, _13798_);
  and (_13804_, _13803_, _13578_);
  or (_13805_, _13804_, _03137_);
  and (_13806_, _08010_, _08006_);
  nor (_13807_, _13806_, _08011_);
  or (_13808_, _13807_, _03138_);
  and (_13809_, _13808_, _08031_);
  and (_13810_, _13809_, _13805_);
  and (_13811_, _08040_, _08038_);
  nor (_13812_, _13811_, _08041_);
  and (_13813_, _13812_, _07950_);
  or (_13814_, _13813_, _08029_);
  or (_13815_, _13814_, _13810_);
  nand (_13816_, _08029_, _02549_);
  and (_13817_, _13816_, _07259_);
  and (_13818_, _13817_, _13815_);
  or (_13819_, _07242_, _07241_);
  nor (_13820_, _07259_, _07243_);
  and (_13821_, _13820_, _13819_);
  or (_13822_, _13821_, _13818_);
  and (_13823_, _13822_, _08064_);
  nor (_13824_, _08084_, _08083_);
  or (_13825_, _08085_, _08064_);
  nor (_13826_, _13825_, _13824_);
  or (_13827_, _13826_, _02899_);
  or (_13828_, _13827_, _13823_);
  and (_13829_, _08114_, _07732_);
  nor (_13830_, _13829_, _08115_);
  or (_13831_, _13830_, _02901_);
  and (_13832_, _13831_, _08106_);
  and (_13833_, _13832_, _13828_);
  nor (_13834_, _08157_, _08156_);
  nor (_13835_, _13834_, _08158_);
  and (_13836_, _13835_, _08103_);
  or (_13837_, _13836_, _08135_);
  or (_13838_, _13837_, _13833_);
  and (_13839_, _13838_, _13575_);
  or (_13840_, _13839_, _03166_);
  or (_13841_, _13616_, _03563_);
  and (_13842_, _13841_, _08180_);
  and (_13843_, _13842_, _13840_);
  nor (_13844_, _08209_, _08185_);
  nor (_13845_, _13844_, _08180_);
  or (_13846_, _13845_, _08184_);
  or (_13847_, _13846_, _13843_);
  nand (_13848_, _08184_, _06984_);
  and (_13849_, _13848_, _02501_);
  and (_13850_, _13849_, _13847_);
  nor (_13851_, _13650_, _02501_);
  or (_13852_, _13851_, _03174_);
  or (_13853_, _13852_, _13850_);
  nor (_13854_, _13614_, _13583_);
  nand (_13855_, _13854_, _03174_);
  and (_13856_, _13855_, _08202_);
  and (_13857_, _13856_, _13853_);
  and (_13858_, _13844_, _08201_);
  or (_13859_, _13858_, _08208_);
  or (_13860_, _13859_, _13857_);
  nand (_13861_, _08208_, _06984_);
  and (_13862_, _13861_, _34698_);
  and (_13863_, _13862_, _13860_);
  or (_13864_, _13863_, _13574_);
  and (_35165_, _13864_, _36029_);
  nor (_13865_, _34698_, _06984_);
  nand (_13866_, _08029_, _02618_);
  nand (_13867_, _07865_, _08151_);
  nand (_13868_, _07263_, _07236_);
  not (_13869_, _02835_);
  nand (_13870_, _02976_, _13869_);
  and (_13871_, _13870_, _02532_);
  nor (_13872_, _13871_, _03356_);
  or (_13873_, _07813_, _08152_);
  nor (_13874_, _07783_, _03260_);
  nor (_13875_, _04712_, _06984_);
  nor (_13876_, _07272_, _04440_);
  nor (_13877_, _13876_, _13875_);
  nand (_13878_, _13877_, _06793_);
  nor (_13879_, _07705_, _07703_);
  nor (_13880_, _13879_, _07706_);
  and (_13881_, _07735_, \oc8051_golden_model_1.PSW [7]);
  not (_13882_, _13881_);
  nor (_13883_, _13882_, _13880_);
  and (_13884_, _13882_, _13880_);
  or (_13885_, _13884_, _13883_);
  or (_13886_, _13885_, _02997_);
  and (_13887_, _13886_, _07277_);
  nand (_13888_, _07431_, _04440_);
  not (_13889_, _07440_);
  nand (_13890_, _13889_, _04440_);
  or (_13891_, _07442_, _06984_);
  nand (_13892_, _07442_, _06984_);
  and (_13893_, _13892_, _13891_);
  nand (_13894_, _13893_, _09203_);
  and (_13895_, _13894_, _13890_);
  or (_13896_, _13895_, _02954_);
  nand (_13897_, _07670_, _02954_);
  and (_13898_, _13897_, _09202_);
  and (_13899_, _13898_, _13896_);
  or (_13900_, _13899_, _03818_);
  or (_13901_, _13358_, _06177_);
  and (_13902_, _13901_, _13900_);
  and (_13903_, _13902_, _03821_);
  nor (_13904_, _10849_, _07272_);
  nor (_13905_, _13904_, _13875_);
  nor (_13906_, _13905_, _03821_);
  or (_13907_, _13906_, _07455_);
  or (_13908_, _13907_, _13903_);
  nand (_13909_, _13620_, \oc8051_golden_model_1.ACC [2]);
  and (_13910_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_13911_, _13910_, _07461_);
  or (_13912_, _13911_, _13620_);
  and (_13913_, _13912_, _13909_);
  nand (_13914_, _13913_, _07455_);
  and (_13915_, _13914_, _02951_);
  and (_13916_, _13915_, _13908_);
  nor (_13917_, _05331_, _06984_);
  and (_13918_, _10853_, _05331_);
  nor (_13919_, _13918_, _13917_);
  nor (_13920_, _13919_, _02892_);
  nor (_13921_, _13877_, _03327_);
  or (_13922_, _13921_, _07431_);
  or (_13923_, _13922_, _13920_);
  or (_13924_, _13923_, _13916_);
  and (_13925_, _13924_, _13888_);
  or (_13926_, _13925_, _03413_);
  or (_13927_, _06177_, _03849_);
  and (_13928_, _13927_, _02959_);
  and (_13929_, _13928_, _13926_);
  nor (_13930_, _07670_, _02959_);
  or (_13931_, _13930_, _07497_);
  or (_13932_, _13931_, _13929_);
  nand (_13933_, _07497_, _06833_);
  and (_13934_, _13933_, _13932_);
  or (_13935_, _13934_, _02887_);
  and (_13936_, _10838_, _05331_);
  nor (_13937_, _13936_, _13917_);
  nand (_13938_, _13937_, _02887_);
  and (_13939_, _13938_, _02881_);
  and (_13940_, _13939_, _13935_);
  and (_13941_, _13918_, _10868_);
  nor (_13942_, _13941_, _13917_);
  nor (_13943_, _13942_, _02881_);
  or (_13944_, _13943_, _06271_);
  or (_13945_, _13944_, _13940_);
  nor (_13946_, _06735_, _06733_);
  nor (_13947_, _13946_, _06736_);
  or (_13948_, _13947_, _06277_);
  and (_13949_, _13948_, _13945_);
  or (_13950_, _13949_, _07427_);
  and (_13951_, _04038_, \oc8051_golden_model_1.ACC [1]);
  and (_13952_, _03817_, _02549_);
  nor (_13953_, _13952_, _07241_);
  nor (_13954_, _13953_, _13951_);
  nor (_13955_, _13954_, _07237_);
  and (_13956_, _13954_, _07237_);
  nor (_13957_, _13956_, _13955_);
  nor (_13958_, _13454_, _07241_);
  not (_13959_, _13958_);
  or (_13960_, _13959_, _13957_);
  and (_13961_, _13960_, \oc8051_golden_model_1.PSW [7]);
  nor (_13962_, _13957_, \oc8051_golden_model_1.PSW [7]);
  or (_13963_, _13962_, _13961_);
  nand (_13964_, _13959_, _13957_);
  and (_13965_, _13964_, _13963_);
  nand (_13966_, _13965_, _07427_);
  and (_13967_, _13966_, _07344_);
  and (_13968_, _13967_, _13950_);
  and (_13969_, _05893_, \oc8051_golden_model_1.ACC [1]);
  and (_13970_, _06174_, _02549_);
  nor (_13971_, _13970_, _08083_);
  nor (_13972_, _13971_, _13969_);
  nor (_13973_, _08079_, _13972_);
  and (_13974_, _08079_, _13972_);
  nor (_13975_, _13974_, _13973_);
  nor (_13976_, _13340_, _08083_);
  not (_13977_, _13976_);
  or (_13978_, _13977_, _13975_);
  and (_13979_, _13978_, \oc8051_golden_model_1.PSW [7]);
  nor (_13980_, _13975_, \oc8051_golden_model_1.PSW [7]);
  or (_13981_, _13980_, _13979_);
  nand (_13982_, _13977_, _13975_);
  and (_13983_, _13982_, _13981_);
  or (_13984_, _13983_, _07344_);
  nand (_13985_, _13984_, _02997_);
  or (_13986_, _13985_, _13968_);
  and (_13987_, _13986_, _13887_);
  nor (_13988_, _02832_, \oc8051_golden_model_1.ACC [0]);
  nor (_13989_, _13988_, _08156_);
  nor (_13990_, _13989_, _10002_);
  nor (_13991_, _08152_, _13990_);
  and (_13992_, _08152_, _13990_);
  nor (_13993_, _13992_, _13991_);
  not (_13994_, _09318_);
  or (_13995_, _13994_, _13993_);
  and (_13996_, _13995_, \oc8051_golden_model_1.PSW [7]);
  nor (_13997_, _13993_, \oc8051_golden_model_1.PSW [7]);
  or (_13998_, _13997_, _13996_);
  nand (_13999_, _13994_, _13993_);
  and (_14000_, _13999_, _13998_);
  nor (_14001_, _14000_, _07277_);
  or (_14002_, _14001_, _02585_);
  or (_14003_, _14002_, _13987_);
  nand (_14004_, _03260_, _02585_);
  and (_14005_, _14004_, _02875_);
  and (_14006_, _14005_, _14003_);
  nor (_14007_, _10886_, _07755_);
  nor (_14008_, _14007_, _13917_);
  nor (_14009_, _14008_, _02875_);
  or (_14010_, _14009_, _06793_);
  or (_14011_, _14010_, _14006_);
  and (_14012_, _14011_, _13878_);
  or (_14013_, _14012_, _02855_);
  and (_14014_, _06177_, _04712_);
  nor (_14015_, _14014_, _13875_);
  nand (_14016_, _14015_, _02855_);
  and (_14017_, _14016_, _02851_);
  and (_14018_, _14017_, _14013_);
  nor (_14019_, _10943_, _07272_);
  nor (_14020_, _14019_, _13875_);
  nor (_14021_, _14020_, _02851_);
  or (_14022_, _14021_, _06807_);
  or (_14023_, _14022_, _14018_);
  or (_14024_, _07004_, _06813_);
  and (_14025_, _14024_, _14023_);
  and (_14026_, _14025_, _02584_);
  nor (_14027_, _03260_, _02584_);
  or (_14028_, _14027_, _03014_);
  or (_14029_, _14028_, _14026_);
  and (_14030_, _04712_, _05727_);
  nor (_14031_, _14030_, _13875_);
  nand (_14032_, _14031_, _03014_);
  and (_14033_, _14032_, _07783_);
  and (_14034_, _14033_, _14029_);
  or (_14035_, _14034_, _13874_);
  and (_14036_, _14035_, _07792_);
  and (_14037_, _07791_, _07237_);
  or (_14038_, _14037_, _07793_);
  or (_14039_, _14038_, _14036_);
  or (_14040_, _13732_, _07237_);
  and (_14041_, _14040_, _13739_);
  and (_14042_, _14041_, _14039_);
  and (_14043_, _07796_, _07237_);
  or (_14044_, _14043_, _07802_);
  or (_14045_, _14044_, _14042_);
  or (_14046_, _08079_, _07803_);
  and (_14047_, _14046_, _07814_);
  and (_14048_, _14047_, _14045_);
  or (_14049_, _10831_, _07812_);
  and (_14050_, _14049_, _09451_);
  or (_14051_, _14050_, _14048_);
  and (_14052_, _14051_, _13873_);
  or (_14053_, _14052_, _03021_);
  and (_14054_, _10835_, _04712_);
  nor (_14055_, _14054_, _13875_);
  nand (_14056_, _14055_, _03021_);
  and (_14057_, _14056_, _03131_);
  and (_14058_, _14057_, _14053_);
  and (_14059_, _13875_, _03130_);
  or (_14060_, _14059_, _14058_);
  and (_14061_, _14060_, _13872_);
  and (_14062_, _04148_, _02532_);
  or (_14063_, _14062_, _07235_);
  and (_14064_, _14063_, _07827_);
  or (_14065_, _14064_, _14061_);
  not (_14066_, _14062_);
  or (_14067_, _14066_, _07235_);
  and (_14068_, _14067_, _07265_);
  and (_14069_, _14068_, _14065_);
  and (_14070_, _08077_, _03513_);
  or (_14071_, _14070_, _03141_);
  or (_14072_, _14071_, _14069_);
  or (_14073_, _10829_, _07838_);
  and (_14074_, _14073_, _07837_);
  and (_14075_, _14074_, _14072_);
  and (_14076_, _07836_, _08150_);
  or (_14077_, _14076_, _14075_);
  and (_14078_, _14077_, _05274_);
  or (_14079_, _14031_, _10830_);
  nor (_14080_, _14079_, _05274_);
  or (_14081_, _14080_, _07263_);
  or (_14082_, _14081_, _14078_);
  and (_14083_, _14082_, _13868_);
  or (_14084_, _14083_, _07852_);
  nand (_14085_, _07852_, _07236_);
  and (_14086_, _14085_, _07854_);
  and (_14087_, _14086_, _14084_);
  nor (_14088_, _07236_, _07854_);
  or (_14089_, _14088_, _07858_);
  or (_14090_, _14089_, _14087_);
  nand (_14091_, _08078_, _07858_);
  and (_14092_, _14091_, _03126_);
  and (_14093_, _14092_, _14090_);
  nand (_14094_, _10830_, _07868_);
  and (_14095_, _14094_, _07867_);
  or (_14096_, _14095_, _14093_);
  and (_14097_, _14096_, _13867_);
  or (_14098_, _14097_, _03036_);
  nor (_14099_, _10833_, _07272_);
  nor (_14100_, _14099_, _13875_);
  nand (_14101_, _14100_, _03036_);
  and (_14102_, _14101_, _07889_);
  and (_14103_, _14102_, _14098_);
  and (_14104_, _07900_, _07557_);
  nor (_14105_, _14104_, _07901_);
  and (_14106_, _14105_, _10171_);
  or (_14107_, _14106_, _14103_);
  and (_14108_, _14107_, _07922_);
  and (_14109_, _07933_, _07387_);
  nor (_14110_, _14109_, _07934_);
  and (_14111_, _14110_, _07917_);
  or (_14112_, _14111_, _03137_);
  or (_14113_, _14112_, _14108_);
  and (_14114_, _08012_, _08000_);
  nor (_14115_, _14114_, _08013_);
  or (_14116_, _14115_, _03138_);
  and (_14117_, _14116_, _08031_);
  and (_14118_, _14117_, _14113_);
  and (_14119_, _08042_, _07317_);
  nor (_14120_, _14119_, _08043_);
  and (_14121_, _14120_, _07950_);
  or (_14122_, _14121_, _08029_);
  or (_14123_, _14122_, _14118_);
  and (_14124_, _14123_, _13866_);
  or (_14125_, _14124_, _07258_);
  and (_14126_, _07244_, _07238_);
  nor (_14127_, _14126_, _07245_);
  or (_14128_, _14127_, _07259_);
  and (_14129_, _14128_, _08064_);
  and (_14130_, _14129_, _14125_);
  and (_14131_, _08086_, _08080_);
  nor (_14132_, _14131_, _08087_);
  and (_14133_, _14132_, _07217_);
  or (_14134_, _14133_, _08105_);
  or (_14135_, _14134_, _14130_);
  and (_14136_, _08116_, _07705_);
  nor (_14137_, _14136_, _08117_);
  or (_14138_, _14137_, _02901_);
  and (_14139_, _08159_, _08153_);
  nor (_14140_, _14139_, _08160_);
  or (_14141_, _14140_, _08106_);
  and (_14142_, _14141_, _08136_);
  and (_14143_, _14142_, _14138_);
  and (_14144_, _14143_, _14135_);
  and (_14145_, _08135_, \oc8051_golden_model_1.ACC [1]);
  or (_14146_, _14145_, _03166_);
  or (_14147_, _14146_, _14144_);
  nand (_14148_, _13905_, _03166_);
  and (_14149_, _14148_, _08180_);
  and (_14150_, _14149_, _14147_);
  and (_14151_, _07461_, _02549_);
  nor (_14152_, _08185_, _06984_);
  or (_14153_, _14152_, _14151_);
  and (_14154_, _14153_, _08179_);
  or (_14155_, _14154_, _08184_);
  or (_14156_, _14155_, _14150_);
  nand (_14157_, _08184_, _02701_);
  and (_14158_, _14157_, _02501_);
  and (_14159_, _14158_, _14156_);
  nor (_14160_, _13937_, _02501_);
  or (_14161_, _14160_, _03174_);
  or (_14162_, _14161_, _14159_);
  and (_14163_, _11008_, _04712_);
  nor (_14164_, _14163_, _13875_);
  nand (_14165_, _14164_, _03174_);
  and (_14166_, _14165_, _08202_);
  and (_14167_, _14166_, _14162_);
  and (_14168_, _08209_, \oc8051_golden_model_1.ACC [2]);
  nor (_14169_, _08209_, \oc8051_golden_model_1.ACC [2]);
  nor (_14170_, _14169_, _14168_);
  nor (_14171_, _14170_, _08208_);
  nor (_14172_, _14171_, _09765_);
  or (_14173_, _14172_, _14167_);
  nand (_14174_, _08208_, _02701_);
  and (_14175_, _14174_, _34698_);
  and (_14176_, _14175_, _14173_);
  or (_14177_, _14176_, _13865_);
  and (_35166_, _14177_, _36029_);
  nor (_14178_, _34698_, _02701_);
  nor (_14179_, _07231_, _07233_);
  nor (_14180_, _14179_, _07246_);
  and (_14181_, _14179_, _07246_);
  nor (_14182_, _14181_, _14180_);
  nand (_14183_, _14182_, _07258_);
  and (_14184_, _07902_, _07552_);
  nor (_14185_, _14184_, _07903_);
  and (_14186_, _14185_, _07888_);
  or (_14187_, _14186_, _07889_);
  and (_14188_, _04148_, _02537_);
  nor (_14189_, _04712_, _02701_);
  and (_14190_, _11032_, _04712_);
  nor (_14191_, _14190_, _14189_);
  nand (_14192_, _14191_, _03021_);
  nor (_14193_, _07272_, _04242_);
  nor (_14194_, _14193_, _14189_);
  nand (_14195_, _14194_, _06793_);
  and (_14196_, _06029_, \oc8051_golden_model_1.ACC [2]);
  nor (_14197_, _13973_, _14196_);
  nor (_14198_, _08075_, _08073_);
  nor (_14199_, _14198_, _14197_);
  and (_14200_, _14198_, _14197_);
  nor (_14201_, _14200_, _14199_);
  and (_14202_, _14201_, \oc8051_golden_model_1.PSW [7]);
  nor (_14203_, _14201_, \oc8051_golden_model_1.PSW [7]);
  nor (_14204_, _14203_, _14202_);
  and (_14205_, _14204_, _13979_);
  nor (_14206_, _14204_, _13979_);
  or (_14207_, _14206_, _14205_);
  nand (_14208_, _14207_, _03441_);
  nor (_14209_, _05331_, _02701_);
  and (_14210_, _11037_, _05331_);
  and (_14211_, _14210_, _11066_);
  nor (_14212_, _14211_, _14209_);
  nor (_14213_, _14212_, _02881_);
  nand (_14214_, _07431_, _04242_);
  or (_14215_, _13358_, _06176_);
  nor (_14216_, _07651_, _07433_);
  nor (_14217_, _07440_, _04242_);
  nand (_14218_, _07442_, _02701_);
  or (_14219_, _07442_, _02701_);
  and (_14220_, _14219_, _07436_);
  nand (_14221_, _14220_, _14218_);
  and (_14222_, _14221_, _07440_);
  or (_14223_, _14222_, _14217_);
  and (_14224_, _14223_, _07433_);
  or (_14225_, _14224_, _14216_);
  and (_14226_, _14225_, _09202_);
  or (_14227_, _14226_, _03818_);
  and (_14228_, _14227_, _03821_);
  and (_14229_, _14228_, _14215_);
  nor (_14230_, _11040_, _07272_);
  nor (_14231_, _14230_, _14189_);
  nor (_14232_, _14231_, _03821_);
  or (_14233_, _14232_, _07455_);
  or (_14234_, _14233_, _14229_);
  not (_14235_, \oc8051_golden_model_1.PSW [6]);
  nor (_14236_, _07461_, _14235_);
  nor (_14237_, _14236_, \oc8051_golden_model_1.ACC [3]);
  nor (_14238_, _14237_, _07462_);
  not (_14239_, _14238_);
  nand (_14240_, _14239_, _07455_);
  and (_14241_, _14240_, _14234_);
  or (_14242_, _14241_, _02891_);
  nor (_14243_, _14210_, _14209_);
  nand (_14244_, _14243_, _02891_);
  and (_14245_, _14244_, _03327_);
  and (_14246_, _14245_, _14242_);
  nor (_14247_, _14194_, _03327_);
  or (_14248_, _14247_, _07431_);
  or (_14249_, _14248_, _14246_);
  and (_14250_, _14249_, _14214_);
  or (_14251_, _14250_, _03413_);
  or (_14252_, _06176_, _03849_);
  and (_14253_, _14252_, _02959_);
  and (_14254_, _14253_, _14251_);
  nor (_14255_, _07651_, _02959_);
  or (_14256_, _14255_, _07497_);
  or (_14257_, _14256_, _14254_);
  nand (_14258_, _07497_, _05768_);
  and (_14259_, _14258_, _14257_);
  or (_14260_, _14259_, _02887_);
  and (_14261_, _11035_, _05331_);
  nor (_14262_, _14261_, _14209_);
  nand (_14263_, _14262_, _02887_);
  and (_14264_, _14263_, _02881_);
  and (_14265_, _14264_, _14260_);
  or (_14266_, _14265_, _14213_);
  and (_14267_, _14266_, _06277_);
  nor (_14268_, _06738_, _06736_);
  nor (_14269_, _14268_, _06739_);
  nand (_14270_, _14269_, _06271_);
  nand (_14271_, _14270_, _10051_);
  or (_14272_, _14271_, _14267_);
  and (_14273_, _04440_, \oc8051_golden_model_1.ACC [2]);
  nor (_14274_, _13955_, _14273_);
  and (_14275_, _14274_, _14179_);
  nor (_14276_, _14274_, _14179_);
  or (_14277_, _14276_, _14275_);
  nor (_14278_, _14277_, _07319_);
  and (_14279_, _14277_, _07319_);
  nor (_14280_, _14279_, _14278_);
  and (_14281_, _14280_, _13961_);
  nor (_14282_, _14280_, _13961_);
  nor (_14283_, _14282_, _14281_);
  and (_14284_, _14283_, _10066_);
  or (_14285_, _14284_, _07426_);
  and (_14286_, _14285_, _14272_);
  and (_14287_, _14283_, _03444_);
  or (_14288_, _14287_, _03441_);
  or (_14289_, _14288_, _14286_);
  and (_14290_, _14289_, _14208_);
  or (_14291_, _14290_, _02992_);
  not (_14292_, _07730_);
  and (_14293_, _14292_, _07707_);
  nor (_14294_, _14292_, _07707_);
  nor (_14295_, _14294_, _14293_);
  not (_14296_, _13883_);
  and (_14297_, _14296_, _14295_);
  or (_14298_, _14297_, _07737_);
  or (_14299_, _14298_, _02997_);
  and (_14300_, _14299_, _07277_);
  and (_14301_, _14300_, _14291_);
  and (_14302_, _03260_, \oc8051_golden_model_1.ACC [2]);
  nor (_14303_, _13991_, _14302_);
  nor (_14304_, _09319_, _14303_);
  and (_14305_, _09319_, _14303_);
  nor (_14306_, _14305_, _14304_);
  and (_14307_, _14306_, \oc8051_golden_model_1.PSW [7]);
  nor (_14308_, _14306_, \oc8051_golden_model_1.PSW [7]);
  nor (_14309_, _14308_, _14307_);
  and (_14310_, _14309_, _13996_);
  nor (_14311_, _14309_, _13996_);
  or (_14312_, _14311_, _14310_);
  nor (_14313_, _14312_, _07277_);
  or (_14314_, _14313_, _02585_);
  or (_14315_, _14314_, _14301_);
  nand (_14316_, _02799_, _02585_);
  and (_14317_, _14316_, _02875_);
  and (_14318_, _14317_, _14315_);
  nor (_14319_, _11083_, _07755_);
  nor (_14320_, _14319_, _14209_);
  nor (_14321_, _14320_, _02875_);
  or (_14322_, _14321_, _06793_);
  or (_14323_, _14322_, _14318_);
  and (_14324_, _14323_, _14195_);
  or (_14325_, _14324_, _02855_);
  and (_14326_, _06176_, _04712_);
  nor (_14327_, _14326_, _14189_);
  nand (_14328_, _14327_, _02855_);
  and (_14329_, _14328_, _02851_);
  and (_14330_, _14329_, _14325_);
  nor (_14331_, _11143_, _07272_);
  nor (_14332_, _14331_, _14189_);
  nor (_14333_, _14332_, _02851_);
  or (_14334_, _14333_, _06807_);
  or (_14335_, _14334_, _14330_);
  or (_14336_, _06948_, _06813_);
  and (_14337_, _14336_, _14335_);
  and (_14338_, _14337_, _02584_);
  nor (_14339_, _02799_, _02584_);
  or (_14340_, _14339_, _03014_);
  or (_14341_, _14340_, _14338_);
  and (_14342_, _04712_, _05664_);
  nor (_14343_, _14342_, _14189_);
  nand (_14344_, _14343_, _03014_);
  and (_14345_, _14344_, _07783_);
  and (_14346_, _14345_, _14341_);
  nor (_14347_, _07783_, _02799_);
  or (_14348_, _14347_, _07799_);
  or (_14349_, _14348_, _14346_);
  or (_14350_, _07798_, _14179_);
  and (_14351_, _14350_, _07803_);
  and (_14352_, _14351_, _14349_);
  and (_14353_, _14198_, _07802_);
  or (_14354_, _14353_, _03132_);
  or (_14355_, _14354_, _14352_);
  or (_14356_, _11028_, _07814_);
  and (_14357_, _14356_, _07813_);
  and (_14358_, _14357_, _14355_);
  and (_14359_, _07812_, _09319_);
  or (_14360_, _14359_, _03021_);
  or (_14361_, _14360_, _14358_);
  and (_14362_, _14361_, _14192_);
  or (_14363_, _14362_, _03130_);
  or (_14364_, _14189_, _03131_);
  and (_14365_, _14364_, _13872_);
  and (_14366_, _14365_, _14363_);
  or (_14367_, _14062_, _07233_);
  and (_14368_, _14367_, _07827_);
  or (_14369_, _14368_, _14366_);
  or (_14370_, _14066_, _07233_);
  and (_14371_, _14370_, _07265_);
  and (_14372_, _14371_, _14369_);
  and (_14373_, _08075_, _03513_);
  or (_14374_, _14373_, _03141_);
  or (_14375_, _14374_, _14372_);
  or (_14376_, _11026_, _07838_);
  and (_14377_, _14376_, _07837_);
  and (_14378_, _14377_, _14375_);
  and (_14379_, _07836_, _08148_);
  or (_14380_, _14379_, _14378_);
  and (_14381_, _14380_, _05274_);
  or (_14382_, _14343_, _11027_);
  nor (_14383_, _14382_, _05274_);
  or (_14384_, _14383_, _07263_);
  or (_14385_, _14384_, _14381_);
  nand (_14386_, _07263_, _07231_);
  nand (_14387_, _14386_, _14385_);
  nor (_14388_, _14387_, _14188_);
  and (_14389_, _14188_, _07232_);
  or (_14390_, _14389_, _07858_);
  or (_14391_, _14390_, _14388_);
  nand (_14392_, _08073_, _07858_);
  and (_14393_, _14392_, _03126_);
  and (_14394_, _14393_, _14391_);
  nand (_14395_, _11027_, _07868_);
  and (_14396_, _14395_, _07867_);
  or (_14397_, _14396_, _14394_);
  nand (_14398_, _07865_, _08149_);
  and (_14399_, _14398_, _05781_);
  and (_14400_, _14399_, _14397_);
  nor (_14401_, _11030_, _07272_);
  nor (_14402_, _14401_, _14189_);
  nor (_14403_, _14402_, _05781_);
  or (_14404_, _14403_, _07883_);
  or (_14405_, _14404_, _14400_);
  and (_14406_, _14405_, _14187_);
  and (_14407_, _14185_, _07918_);
  or (_14408_, _14407_, _07917_);
  or (_14409_, _14408_, _14406_);
  and (_14410_, _07935_, _07382_);
  nor (_14411_, _14410_, _07936_);
  or (_14412_, _14411_, _07922_);
  and (_14413_, _14412_, _03138_);
  and (_14414_, _14413_, _14409_);
  and (_14415_, _08014_, _07994_);
  nor (_14416_, _14415_, _08015_);
  and (_14417_, _14416_, _03137_);
  or (_14418_, _14417_, _07950_);
  or (_14419_, _14418_, _14414_);
  and (_14420_, _08044_, _07315_);
  nor (_14421_, _14420_, _08045_);
  or (_14422_, _14421_, _08031_);
  and (_14423_, _14422_, _08030_);
  and (_14424_, _14423_, _14419_);
  and (_14425_, _08029_, \oc8051_golden_model_1.ACC [2]);
  or (_14426_, _14425_, _07258_);
  or (_14427_, _14426_, _14424_);
  and (_14428_, _14427_, _14183_);
  or (_14429_, _14428_, _07217_);
  nor (_14430_, _08088_, _14198_);
  and (_14431_, _08088_, _14198_);
  nor (_14432_, _14431_, _14430_);
  nand (_14433_, _14432_, _07217_);
  and (_14434_, _14433_, _02901_);
  and (_14435_, _14434_, _14429_);
  nor (_14436_, _08118_, _07730_);
  and (_14437_, _08118_, _07730_);
  nor (_14438_, _14437_, _14436_);
  or (_14439_, _14438_, _08103_);
  and (_14440_, _14439_, _08105_);
  or (_14441_, _14440_, _14435_);
  nor (_14442_, _08161_, _09319_);
  and (_14443_, _08161_, _09319_);
  nor (_14444_, _14443_, _14442_);
  nand (_14445_, _14444_, _08103_);
  and (_14446_, _14445_, _08136_);
  and (_14447_, _14446_, _14441_);
  and (_14448_, _08135_, \oc8051_golden_model_1.ACC [2]);
  or (_14449_, _14448_, _03166_);
  or (_14450_, _14449_, _14447_);
  nand (_14451_, _14231_, _03166_);
  and (_14452_, _14451_, _08180_);
  and (_14453_, _14452_, _14450_);
  nor (_14454_, _14151_, _02701_);
  or (_14455_, _14454_, _08186_);
  and (_14456_, _14455_, _08179_);
  or (_14457_, _14456_, _08184_);
  or (_14458_, _14457_, _14453_);
  nand (_14459_, _08184_, _06885_);
  and (_14460_, _14459_, _02501_);
  and (_14461_, _14460_, _14458_);
  nor (_14462_, _14262_, _02501_);
  or (_14463_, _14462_, _03174_);
  or (_14464_, _14463_, _14461_);
  and (_14465_, _11213_, _04712_);
  nor (_14466_, _14465_, _14189_);
  nand (_14467_, _14466_, _03174_);
  and (_14468_, _14467_, _08202_);
  and (_14469_, _14468_, _14464_);
  or (_14470_, _14168_, \oc8051_golden_model_1.ACC [3]);
  and (_14471_, _14470_, _08210_);
  and (_14472_, _14471_, _08201_);
  or (_14473_, _14472_, _08208_);
  or (_14474_, _14473_, _14469_);
  nand (_14475_, _08208_, _06885_);
  and (_14476_, _14475_, _34698_);
  and (_14477_, _14476_, _14474_);
  or (_14478_, _14477_, _14178_);
  and (_35167_, _14478_, _36029_);
  nor (_14479_, _34698_, _06885_);
  nand (_14480_, _08029_, _02701_);
  and (_14481_, _07937_, _07373_);
  nor (_14482_, _14481_, _07938_);
  or (_14483_, _14482_, _07922_);
  nand (_14484_, _07865_, _08145_);
  nand (_14485_, _13784_, _07229_);
  or (_14486_, _08070_, _07265_);
  nor (_14487_, _04712_, _06885_);
  and (_14488_, _11362_, _04712_);
  nor (_14489_, _14488_, _14487_);
  nand (_14490_, _14489_, _03021_);
  not (_14491_, _03504_);
  nor (_14492_, _05202_, _07272_);
  nor (_14493_, _14492_, _14487_);
  nand (_14494_, _14493_, _06793_);
  and (_14495_, _07738_, _07729_);
  nor (_14496_, _14495_, _07739_);
  nand (_14497_, _14496_, _02992_);
  and (_14498_, _14497_, _07277_);
  nand (_14499_, _07431_, _05202_);
  nor (_14500_, _07640_, _07433_);
  or (_14501_, _06181_, _07436_);
  nor (_14502_, _07440_, _05202_);
  nand (_14503_, _07442_, _06885_);
  or (_14504_, _07442_, _06885_);
  and (_14505_, _14504_, _07436_);
  nand (_14506_, _14505_, _14503_);
  and (_14507_, _14506_, _07440_);
  or (_14508_, _14507_, _14502_);
  and (_14509_, _14508_, _07433_);
  and (_14510_, _14509_, _14501_);
  or (_14511_, _14510_, _14500_);
  and (_14512_, _14511_, _07453_);
  nor (_14513_, _11259_, _07272_);
  nor (_14514_, _14513_, _14487_);
  nor (_14515_, _14514_, _03821_);
  or (_14516_, _14515_, _07455_);
  or (_14517_, _14516_, _14512_);
  nor (_14518_, _07462_, \oc8051_golden_model_1.ACC [4]);
  nor (_14519_, _14518_, _07468_);
  not (_14520_, _14519_);
  nand (_14521_, _14520_, _07455_);
  and (_14522_, _14521_, _02951_);
  and (_14523_, _14522_, _14517_);
  nor (_14524_, _05331_, _06885_);
  and (_14525_, _11245_, _05331_);
  nor (_14526_, _14525_, _14524_);
  nor (_14527_, _14526_, _02892_);
  nor (_14528_, _14493_, _03327_);
  or (_14529_, _14528_, _07431_);
  or (_14530_, _14529_, _14527_);
  or (_14531_, _14530_, _14523_);
  and (_14532_, _14531_, _14499_);
  or (_14533_, _14532_, _03413_);
  or (_14534_, _06181_, _03849_);
  and (_14535_, _14534_, _02959_);
  and (_14536_, _14535_, _14533_);
  nor (_14537_, _07640_, _02959_);
  or (_14538_, _14537_, _07497_);
  or (_14539_, _14538_, _14536_);
  nand (_14540_, _07497_, _02549_);
  and (_14541_, _14540_, _14539_);
  or (_14542_, _14541_, _02887_);
  and (_14543_, _11243_, _05331_);
  nor (_14544_, _14543_, _14524_);
  nand (_14545_, _14544_, _02887_);
  and (_14546_, _14545_, _02881_);
  and (_14547_, _14546_, _14542_);
  and (_14548_, _14525_, _11276_);
  nor (_14549_, _14548_, _14524_);
  nor (_14550_, _14549_, _02881_);
  or (_14551_, _14550_, _06271_);
  or (_14552_, _14551_, _14547_);
  nor (_14553_, _06741_, _06739_);
  nor (_14554_, _14553_, _06743_);
  or (_14555_, _14554_, _06277_);
  and (_14556_, _14555_, _14552_);
  or (_14557_, _14556_, _07427_);
  or (_14558_, _14281_, _14278_);
  nor (_14559_, _04242_, \oc8051_golden_model_1.ACC [3]);
  nand (_14560_, _04242_, \oc8051_golden_model_1.ACC [3]);
  and (_14561_, _14274_, _14560_);
  or (_14562_, _14561_, _14559_);
  nor (_14563_, _14562_, _07230_);
  and (_14564_, _14562_, _07230_);
  nor (_14565_, _14564_, _14563_);
  and (_14566_, _14565_, \oc8051_golden_model_1.PSW [7]);
  nor (_14567_, _14565_, \oc8051_golden_model_1.PSW [7]);
  nor (_14568_, _14567_, _14566_);
  and (_14569_, _14568_, _14558_);
  nor (_14570_, _14568_, _14558_);
  nor (_14571_, _14570_, _14569_);
  or (_14572_, _14571_, _07426_);
  and (_14573_, _14572_, _14557_);
  or (_14574_, _14573_, _03441_);
  or (_14575_, _14205_, _14202_);
  and (_14576_, _06176_, _02701_);
  or (_14577_, _06176_, _02701_);
  and (_14578_, _14577_, _14197_);
  or (_14579_, _14578_, _14576_);
  nor (_14580_, _08072_, _14579_);
  and (_14581_, _08072_, _14579_);
  nor (_14582_, _14581_, _14580_);
  and (_14583_, _14582_, \oc8051_golden_model_1.PSW [7]);
  nor (_14584_, _14582_, \oc8051_golden_model_1.PSW [7]);
  nor (_14585_, _14584_, _14583_);
  and (_14586_, _14585_, _14575_);
  nor (_14587_, _14585_, _14575_);
  nor (_14588_, _14587_, _14586_);
  or (_14589_, _14588_, _07344_);
  and (_14590_, _14589_, _14574_);
  or (_14591_, _14590_, _02992_);
  and (_14592_, _14591_, _14498_);
  or (_14593_, _14310_, _14307_);
  nor (_14594_, _14303_, _10022_);
  nor (_14595_, _14594_, _10021_);
  nor (_14596_, _08147_, _14595_);
  and (_14597_, _08147_, _14595_);
  nor (_14598_, _14597_, _14596_);
  and (_14599_, _14598_, \oc8051_golden_model_1.PSW [7]);
  nor (_14600_, _14598_, \oc8051_golden_model_1.PSW [7]);
  nor (_14601_, _14600_, _14599_);
  and (_14602_, _14601_, _14593_);
  nor (_14603_, _14601_, _14593_);
  nor (_14604_, _14603_, _14602_);
  and (_14605_, _14604_, _07276_);
  or (_14606_, _14605_, _02585_);
  or (_14607_, _14606_, _14592_);
  nand (_14608_, _03625_, _02585_);
  and (_14609_, _14608_, _02875_);
  and (_14610_, _14609_, _14607_);
  nor (_14611_, _11241_, _07755_);
  nor (_14612_, _14611_, _14524_);
  nor (_14613_, _14612_, _02875_);
  or (_14614_, _14613_, _06793_);
  or (_14615_, _14614_, _14610_);
  and (_14616_, _14615_, _14494_);
  or (_14617_, _14616_, _02855_);
  and (_14618_, _06181_, _04712_);
  nor (_14619_, _14618_, _14487_);
  nand (_14620_, _14619_, _02855_);
  and (_14621_, _14620_, _02851_);
  and (_14622_, _14621_, _14617_);
  nor (_14623_, _11348_, _07272_);
  nor (_14624_, _14623_, _14487_);
  nor (_14625_, _14624_, _02851_);
  or (_14626_, _14625_, _06807_);
  or (_14627_, _14626_, _14622_);
  or (_14628_, _06894_, _06813_);
  and (_14629_, _14628_, _14627_);
  and (_14630_, _14629_, _02584_);
  nor (_14631_, _03625_, _02584_);
  or (_14632_, _14631_, _03014_);
  or (_14633_, _14632_, _14630_);
  and (_14634_, _05697_, _04712_);
  nor (_14635_, _14634_, _14487_);
  nand (_14636_, _14635_, _03014_);
  and (_14637_, _14636_, _07783_);
  and (_14638_, _14637_, _14633_);
  nor (_14639_, _07783_, _03625_);
  or (_14640_, _14639_, _07791_);
  or (_14641_, _14640_, _14638_);
  or (_14642_, _07792_, _07230_);
  and (_14643_, _14642_, _13732_);
  and (_14644_, _14643_, _14641_);
  and (_14645_, _07793_, _07230_);
  or (_14646_, _14645_, _07796_);
  or (_14647_, _14646_, _14644_);
  and (_14648_, _02574_, _02546_);
  and (_14649_, _14648_, _02511_);
  not (_14650_, _14649_);
  or (_14651_, _13739_, _07230_);
  and (_14652_, _14651_, _14650_);
  and (_14653_, _14652_, _14647_);
  and (_14654_, _14649_, _08072_);
  or (_14655_, _14654_, _14653_);
  and (_14656_, _14655_, _14491_);
  and (_14657_, _08072_, _03504_);
  or (_14658_, _14657_, _03132_);
  or (_14659_, _14658_, _14656_);
  or (_14660_, _11368_, _07814_);
  and (_14661_, _14660_, _07813_);
  and (_14662_, _14661_, _14659_);
  nor (_14663_, _07813_, _08146_);
  or (_14664_, _14663_, _03021_);
  or (_14665_, _14664_, _14662_);
  and (_14666_, _14665_, _14490_);
  or (_14667_, _14666_, _03130_);
  or (_14668_, _14487_, _03131_);
  and (_14669_, _14668_, _07828_);
  and (_14670_, _14669_, _14667_);
  and (_14671_, _07827_, _07228_);
  or (_14672_, _14671_, _03513_);
  or (_14673_, _14672_, _14670_);
  and (_14674_, _14673_, _14486_);
  or (_14675_, _14674_, _03141_);
  or (_14676_, _11366_, _07838_);
  and (_14677_, _14676_, _07837_);
  and (_14678_, _14677_, _14675_);
  and (_14679_, _07836_, _08144_);
  or (_14680_, _14679_, _14678_);
  and (_14682_, _14680_, _05274_);
  or (_14683_, _14635_, _11367_);
  nor (_14684_, _14683_, _05274_);
  or (_14685_, _14684_, _13784_);
  or (_14686_, _14685_, _14682_);
  and (_14687_, _14686_, _14485_);
  or (_14688_, _14687_, _07858_);
  nand (_14689_, _08071_, _07858_);
  and (_14690_, _14689_, _03126_);
  and (_14691_, _14690_, _14688_);
  nand (_14693_, _11367_, _07868_);
  and (_14694_, _14693_, _07867_);
  or (_14695_, _14694_, _14691_);
  and (_14696_, _14695_, _14484_);
  or (_14697_, _14696_, _03036_);
  nor (_14698_, _11361_, _07272_);
  nor (_14699_, _14698_, _14487_);
  nand (_14700_, _14699_, _03036_);
  and (_14701_, _14700_, _07889_);
  and (_14702_, _14701_, _14697_);
  and (_14704_, _07904_, _07543_);
  nor (_14705_, _14704_, _07905_);
  and (_14706_, _14705_, _10171_);
  or (_14707_, _14706_, _07917_);
  or (_14708_, _14707_, _14702_);
  and (_14709_, _14708_, _14483_);
  or (_14710_, _14709_, _03137_);
  and (_14711_, _08016_, _07988_);
  nor (_14712_, _14711_, _08017_);
  or (_14713_, _14712_, _03138_);
  and (_14715_, _14713_, _08031_);
  and (_14716_, _14715_, _14710_);
  and (_14717_, _08046_, _07304_);
  nor (_14718_, _14717_, _08047_);
  and (_14719_, _14718_, _07950_);
  or (_14720_, _14719_, _08029_);
  or (_14721_, _14720_, _14716_);
  and (_14722_, _14721_, _14480_);
  or (_14723_, _14722_, _07258_);
  nor (_14724_, _07248_, _07230_);
  nor (_14726_, _14724_, _07249_);
  or (_14727_, _14726_, _07259_);
  and (_14728_, _14727_, _08064_);
  and (_14729_, _14728_, _14723_);
  nor (_14730_, _08090_, _08072_);
  nor (_14731_, _14730_, _08091_);
  and (_14732_, _14731_, _07217_);
  or (_14733_, _14732_, _08105_);
  or (_14734_, _14733_, _14729_);
  nor (_14735_, _08122_, _08110_);
  nor (_14737_, _14735_, _08123_);
  or (_14738_, _14737_, _02901_);
  nor (_14739_, _08163_, _08147_);
  nor (_14740_, _14739_, _08164_);
  or (_14741_, _14740_, _08106_);
  and (_14742_, _14741_, _08136_);
  and (_14743_, _14742_, _14738_);
  and (_14744_, _14743_, _14734_);
  and (_14745_, _08135_, \oc8051_golden_model_1.ACC [3]);
  or (_14746_, _14745_, _03166_);
  or (_14748_, _14746_, _14744_);
  nand (_14749_, _14514_, _03166_);
  and (_14750_, _14749_, _08180_);
  and (_14751_, _14750_, _14748_);
  and (_14752_, _08186_, _06885_);
  nor (_14753_, _08186_, _06885_);
  nor (_14754_, _14753_, _14752_);
  not (_14755_, _14754_);
  and (_14756_, _14755_, _08179_);
  or (_14757_, _14756_, _08184_);
  or (_14759_, _14757_, _14751_);
  nand (_14760_, _08184_, _06879_);
  and (_14761_, _14760_, _02501_);
  and (_14762_, _14761_, _14759_);
  nor (_14763_, _14544_, _02501_);
  or (_14764_, _14763_, _03174_);
  or (_14765_, _14764_, _14762_);
  and (_14766_, _11417_, _04712_);
  nor (_14767_, _14766_, _14487_);
  nand (_14768_, _14767_, _03174_);
  and (_14770_, _14768_, _08202_);
  and (_14771_, _14770_, _14765_);
  and (_14772_, _08210_, _06885_);
  nor (_14773_, _14772_, _08211_);
  and (_14774_, _14773_, _08201_);
  or (_14775_, _14774_, _08208_);
  or (_14776_, _14775_, _14771_);
  nand (_14777_, _08208_, _06879_);
  and (_14778_, _14777_, _34698_);
  and (_14779_, _14778_, _14776_);
  or (_14781_, _14779_, _14479_);
  and (_35168_, _14781_, _36029_);
  nor (_14782_, _34698_, _06879_);
  and (_14783_, _07250_, _07227_);
  nor (_14784_, _14783_, _07251_);
  or (_14785_, _14784_, _07259_);
  and (_14786_, _07906_, _07536_);
  nor (_14787_, _14786_, _07907_);
  or (_14788_, _14787_, _07889_);
  nand (_14789_, _07263_, _07225_);
  or (_14791_, _11434_, _07838_);
  and (_14792_, _14791_, _07837_);
  nor (_14793_, _04712_, _06879_);
  and (_14794_, _11562_, _04712_);
  nor (_14795_, _14794_, _14793_);
  nand (_14796_, _14795_, _03021_);
  nor (_14797_, _08069_, _08068_);
  or (_14798_, _14797_, _14491_);
  nor (_14799_, _04896_, _07272_);
  nor (_14800_, _14799_, _14793_);
  nand (_14802_, _14800_, _06793_);
  and (_14803_, _03625_, \oc8051_golden_model_1.ACC [4]);
  nor (_14804_, _14596_, _14803_);
  nor (_14805_, _08142_, _14804_);
  and (_14806_, _08142_, _14804_);
  nor (_14807_, _14806_, _14805_);
  and (_14808_, _14807_, \oc8051_golden_model_1.PSW [7]);
  nor (_14809_, _14807_, \oc8051_golden_model_1.PSW [7]);
  nor (_14810_, _14809_, _14808_);
  nor (_14811_, _14602_, _14599_);
  not (_14813_, _14811_);
  and (_14814_, _14813_, _14810_);
  nor (_14815_, _14813_, _14810_);
  nor (_14816_, _14815_, _14814_);
  or (_14817_, _14816_, _07277_);
  nor (_14818_, _05331_, _06879_);
  and (_14819_, _11459_, _05331_);
  and (_14820_, _14819_, _11474_);
  nor (_14821_, _14820_, _14818_);
  nor (_14822_, _14821_, _02881_);
  nand (_14824_, _07431_, _04896_);
  nor (_14825_, _07624_, _07433_);
  or (_14826_, _06180_, _07436_);
  nor (_14827_, _07440_, _04896_);
  nand (_14828_, _07442_, _06879_);
  or (_14829_, _07442_, _06879_);
  and (_14830_, _14829_, _07436_);
  nand (_14831_, _14830_, _14828_);
  and (_14832_, _14831_, _07440_);
  or (_14833_, _14832_, _14827_);
  and (_14835_, _14833_, _07433_);
  and (_14836_, _14835_, _14826_);
  or (_14837_, _14836_, _14825_);
  and (_14838_, _14837_, _07453_);
  nor (_14839_, _11445_, _07272_);
  nor (_14840_, _14839_, _14793_);
  nor (_14841_, _14840_, _03821_);
  or (_14842_, _14841_, _07455_);
  or (_14843_, _14842_, _14838_);
  and (_14844_, _09915_, _07470_);
  nor (_14846_, _09915_, _07470_);
  nor (_14847_, _14846_, _14844_);
  nand (_14848_, _14847_, _07455_);
  and (_14849_, _14848_, _02951_);
  and (_14850_, _14849_, _14843_);
  nor (_14851_, _14819_, _14818_);
  nor (_14852_, _14851_, _02892_);
  nor (_14853_, _14800_, _03327_);
  or (_14854_, _14853_, _07431_);
  or (_14855_, _14854_, _14852_);
  or (_14856_, _14855_, _14850_);
  and (_14857_, _14856_, _14824_);
  or (_14858_, _14857_, _03413_);
  or (_14859_, _06180_, _03849_);
  and (_14860_, _14859_, _02959_);
  and (_14861_, _14860_, _14858_);
  nor (_14862_, _07624_, _02959_);
  or (_14863_, _14862_, _07497_);
  or (_14864_, _14863_, _14861_);
  nand (_14865_, _07497_, _02618_);
  and (_14867_, _14865_, _14864_);
  or (_14868_, _14867_, _02887_);
  and (_14869_, _11442_, _05331_);
  nor (_14870_, _14869_, _14818_);
  nand (_14871_, _14870_, _02887_);
  and (_14872_, _14871_, _02881_);
  and (_14873_, _14872_, _14868_);
  or (_14874_, _14873_, _14822_);
  and (_14875_, _14874_, _06277_);
  nor (_14876_, _06745_, _06743_);
  nor (_14878_, _14876_, _06746_);
  and (_14879_, _14878_, _06271_);
  or (_14880_, _14879_, _07427_);
  or (_14881_, _14880_, _14875_);
  and (_14882_, _05202_, \oc8051_golden_model_1.ACC [4]);
  nor (_14883_, _14563_, _14882_);
  nor (_14884_, _14883_, _07226_);
  and (_14885_, _14883_, _07226_);
  nor (_14886_, _14885_, _14884_);
  and (_14887_, _14886_, \oc8051_golden_model_1.PSW [7]);
  nor (_14889_, _14886_, \oc8051_golden_model_1.PSW [7]);
  nor (_14890_, _14889_, _14887_);
  nor (_14891_, _14569_, _14566_);
  not (_14892_, _14891_);
  and (_14893_, _14892_, _14890_);
  nor (_14894_, _14892_, _14890_);
  nor (_14895_, _14894_, _14893_);
  or (_14896_, _14895_, _07426_);
  and (_14897_, _14896_, _14881_);
  or (_14898_, _14897_, _03441_);
  and (_14900_, _06121_, \oc8051_golden_model_1.ACC [4]);
  nor (_14901_, _14580_, _14900_);
  nor (_14902_, _14797_, _14901_);
  and (_14903_, _14797_, _14901_);
  nor (_14904_, _14903_, _14902_);
  and (_14905_, _14904_, \oc8051_golden_model_1.PSW [7]);
  nor (_14906_, _14904_, \oc8051_golden_model_1.PSW [7]);
  nor (_14907_, _14906_, _14905_);
  nor (_14908_, _14586_, _14583_);
  not (_14909_, _14908_);
  and (_14911_, _14909_, _14907_);
  nor (_14912_, _14909_, _14907_);
  nor (_14913_, _14912_, _14911_);
  or (_14914_, _14913_, _07344_);
  and (_14915_, _14914_, _02997_);
  and (_14916_, _14915_, _14898_);
  and (_14917_, _07740_, _07727_);
  nor (_14918_, _14917_, _07741_);
  nand (_14919_, _14918_, _07277_);
  and (_14920_, _14919_, _07597_);
  or (_14922_, _14920_, _14916_);
  and (_14923_, _14922_, _14817_);
  or (_14924_, _14923_, _02585_);
  nand (_14925_, _03215_, _02585_);
  and (_14926_, _14925_, _02875_);
  and (_14927_, _14926_, _14924_);
  nor (_14928_, _11440_, _07755_);
  nor (_14929_, _14928_, _14818_);
  nor (_14930_, _14929_, _02875_);
  or (_14931_, _14930_, _06793_);
  or (_14933_, _14931_, _14927_);
  and (_14934_, _14933_, _14802_);
  or (_14935_, _14934_, _02855_);
  and (_14936_, _06180_, _04712_);
  nor (_14937_, _14936_, _14793_);
  nand (_14938_, _14937_, _02855_);
  and (_14939_, _14938_, _02851_);
  and (_14940_, _14939_, _14935_);
  nor (_14941_, _11546_, _07272_);
  nor (_14942_, _14941_, _14793_);
  nor (_14943_, _14942_, _02851_);
  or (_14944_, _14943_, _06807_);
  or (_14945_, _14944_, _14940_);
  or (_14946_, _06864_, _06813_);
  and (_14947_, _14946_, _14945_);
  and (_14948_, _14947_, _02584_);
  nor (_14949_, _03215_, _02584_);
  or (_14950_, _14949_, _03014_);
  or (_14951_, _14950_, _14948_);
  and (_14952_, _05701_, _04712_);
  nor (_14955_, _14952_, _14793_);
  nand (_14956_, _14955_, _03014_);
  and (_14957_, _14956_, _07783_);
  and (_14958_, _14957_, _14951_);
  nor (_14959_, _07783_, _03215_);
  or (_14960_, _14959_, _07799_);
  or (_14961_, _14960_, _14958_);
  or (_14962_, _07798_, _07226_);
  and (_14963_, _14962_, _14650_);
  and (_14964_, _14963_, _14961_);
  or (_14966_, _14797_, _02465_);
  and (_14967_, _14966_, _07802_);
  or (_14968_, _14967_, _14964_);
  and (_14969_, _14968_, _14798_);
  or (_14970_, _14969_, _03132_);
  or (_14971_, _11436_, _07814_);
  and (_14972_, _14971_, _07813_);
  and (_14973_, _14972_, _14970_);
  and (_14974_, _07812_, _08142_);
  or (_14975_, _14974_, _03021_);
  or (_14977_, _14975_, _14973_);
  and (_14978_, _14977_, _14796_);
  or (_14979_, _14978_, _03130_);
  or (_14980_, _14793_, _03131_);
  and (_14981_, _14980_, _13872_);
  and (_14982_, _14981_, _14979_);
  or (_14983_, _14062_, _07224_);
  and (_14984_, _14983_, _07827_);
  or (_14985_, _14984_, _14982_);
  or (_14986_, _14066_, _07224_);
  and (_14988_, _14986_, _07265_);
  and (_14989_, _14988_, _14985_);
  and (_14990_, _08068_, _03513_);
  or (_14991_, _14990_, _03141_);
  or (_14992_, _14991_, _14989_);
  and (_14993_, _14992_, _14792_);
  and (_14994_, _07836_, _08140_);
  or (_14995_, _14994_, _14993_);
  and (_14996_, _14995_, _05274_);
  or (_14997_, _14955_, _11435_);
  nor (_14999_, _14997_, _05274_);
  or (_15000_, _14999_, _07263_);
  or (_15001_, _15000_, _14996_);
  and (_15002_, _15001_, _14789_);
  or (_15003_, _15002_, _07852_);
  nand (_15004_, _07852_, _07225_);
  and (_15005_, _15004_, _07854_);
  and (_15006_, _15005_, _15003_);
  nor (_15007_, _07225_, _07854_);
  or (_15008_, _15007_, _07858_);
  or (_15010_, _15008_, _15006_);
  nand (_15011_, _08069_, _07858_);
  and (_15012_, _15011_, _03126_);
  and (_15013_, _15012_, _15010_);
  nand (_15014_, _11435_, _07868_);
  and (_15015_, _15014_, _07867_);
  or (_15016_, _15015_, _15013_);
  nand (_15017_, _07865_, _08141_);
  and (_15018_, _15017_, _05781_);
  and (_15019_, _15018_, _15016_);
  nor (_15021_, _11560_, _07272_);
  nor (_15022_, _15021_, _14793_);
  nor (_15023_, _15022_, _05781_);
  or (_15024_, _15023_, _10171_);
  or (_15025_, _15024_, _15019_);
  and (_15026_, _15025_, _14788_);
  or (_15027_, _15026_, _07917_);
  and (_15028_, _07939_, _07371_);
  nor (_15029_, _15028_, _07940_);
  or (_15030_, _15029_, _07922_);
  and (_15032_, _15030_, _03138_);
  and (_15033_, _15032_, _15027_);
  and (_15034_, _08018_, _07982_);
  nor (_15035_, _15034_, _08019_);
  or (_15036_, _15035_, _07950_);
  and (_15037_, _15036_, _08861_);
  or (_15038_, _15037_, _15033_);
  and (_15039_, _08048_, _07299_);
  nor (_15040_, _15039_, _08049_);
  or (_15041_, _15040_, _08031_);
  and (_15043_, _15041_, _08030_);
  and (_15044_, _15043_, _15038_);
  and (_15045_, _08029_, \oc8051_golden_model_1.ACC [4]);
  or (_15046_, _15045_, _07258_);
  or (_15047_, _15046_, _15044_);
  and (_15048_, _15047_, _14785_);
  or (_15049_, _15048_, _07217_);
  nor (_15050_, _08092_, _14797_);
  and (_15051_, _08092_, _14797_);
  or (_15052_, _15051_, _15050_);
  or (_15054_, _15052_, _08064_);
  and (_15055_, _15054_, _02901_);
  and (_15056_, _15055_, _15049_);
  and (_15057_, _08124_, _07724_);
  nor (_15058_, _15057_, _08125_);
  or (_15059_, _15058_, _08103_);
  and (_15060_, _15059_, _08105_);
  or (_15061_, _15060_, _15056_);
  and (_15062_, _08165_, _08143_);
  nor (_15063_, _15062_, _08166_);
  or (_15065_, _15063_, _08106_);
  and (_15066_, _15065_, _08136_);
  and (_15067_, _15066_, _15061_);
  and (_15068_, _08135_, \oc8051_golden_model_1.ACC [4]);
  or (_15069_, _15068_, _03166_);
  or (_15070_, _15069_, _15067_);
  nand (_15071_, _14840_, _03166_);
  and (_15072_, _15071_, _08180_);
  and (_15073_, _15072_, _15070_);
  nor (_15074_, _14752_, _06879_);
  or (_15076_, _15074_, _08187_);
  and (_15077_, _15076_, _08179_);
  or (_15078_, _15077_, _08184_);
  or (_15079_, _15078_, _15073_);
  nand (_15080_, _08184_, _06833_);
  and (_15081_, _15080_, _02501_);
  and (_15082_, _15081_, _15079_);
  nor (_15083_, _14870_, _02501_);
  or (_15084_, _15083_, _03174_);
  or (_15085_, _15084_, _15082_);
  and (_15087_, _11619_, _04712_);
  nor (_15088_, _15087_, _14793_);
  nand (_15089_, _15088_, _03174_);
  and (_15090_, _15089_, _08202_);
  and (_15091_, _15090_, _15085_);
  nor (_15092_, _08211_, \oc8051_golden_model_1.ACC [5]);
  nor (_15093_, _15092_, _08212_);
  and (_15094_, _15093_, _08201_);
  or (_15095_, _15094_, _08208_);
  or (_15096_, _15095_, _15091_);
  nand (_15098_, _08208_, _06833_);
  and (_15099_, _15098_, _34698_);
  and (_15100_, _15099_, _15096_);
  or (_15101_, _15100_, _14782_);
  and (_35169_, _15101_, _36029_);
  nor (_15102_, _34698_, _06833_);
  and (_15103_, _08020_, _07973_);
  nor (_15104_, _15103_, _08021_);
  and (_15105_, _15104_, _03137_);
  nand (_15106_, _07865_, _08138_);
  or (_15108_, _11767_, _07838_);
  and (_15109_, _15108_, _07837_);
  and (_15110_, _07827_, _07221_);
  nor (_15111_, _04712_, _06833_);
  and (_15112_, _11646_, _04712_);
  nor (_15113_, _15112_, _15111_);
  nand (_15114_, _15113_, _03021_);
  and (_15115_, _02842_, _02511_);
  and (_15116_, _15115_, _10788_);
  and (_15117_, _03029_, _02511_);
  not (_15119_, _07223_);
  nand (_15120_, _15119_, _15117_);
  nor (_15121_, _04787_, _07272_);
  nor (_15122_, _15121_, _15111_);
  nand (_15123_, _15122_, _06793_);
  and (_15124_, _07742_, _07723_);
  or (_15125_, _15124_, _07743_);
  or (_15126_, _15125_, _02997_);
  and (_15127_, _15126_, _07277_);
  or (_15128_, _06180_, _06879_);
  and (_15130_, _06180_, _06879_);
  or (_15131_, _14901_, _15130_);
  and (_15132_, _15131_, _15128_);
  nor (_15133_, _15132_, _08067_);
  and (_15134_, _15132_, _08067_);
  nor (_15135_, _15134_, _15133_);
  nor (_15136_, _14911_, _14905_);
  and (_15137_, _15136_, \oc8051_golden_model_1.PSW [7]);
  nor (_15138_, _15137_, _15135_);
  and (_15139_, _15137_, _15135_);
  nor (_15141_, _15139_, _15138_);
  and (_15142_, _15141_, _03441_);
  nand (_15143_, _07431_, _04787_);
  nor (_15144_, _07610_, _07433_);
  or (_15145_, _05847_, _07436_);
  nor (_15146_, _07440_, _04787_);
  and (_15147_, _07442_, _06833_);
  nor (_15148_, _07442_, _06833_);
  or (_15149_, _15148_, _07435_);
  or (_15150_, _15149_, _15147_);
  and (_15152_, _15150_, _07440_);
  or (_15153_, _15152_, _15146_);
  and (_15154_, _15153_, _07433_);
  and (_15155_, _15154_, _15145_);
  or (_15156_, _15155_, _15144_);
  and (_15157_, _15156_, _07453_);
  nor (_15158_, _11636_, _07272_);
  nor (_15159_, _15158_, _15111_);
  nor (_15160_, _15159_, _03821_);
  or (_15161_, _15160_, _07455_);
  or (_15163_, _15161_, _15157_);
  not (_15164_, _07472_);
  nor (_15165_, _14846_, _15164_);
  and (_15166_, _09914_, _07473_);
  nor (_15167_, _15166_, _15165_);
  nand (_15168_, _15167_, _07455_);
  and (_15169_, _15168_, _02951_);
  and (_15170_, _15169_, _15163_);
  nor (_15171_, _05331_, _06833_);
  and (_15172_, _11653_, _05331_);
  nor (_15174_, _15172_, _15171_);
  nor (_15175_, _15174_, _02892_);
  nor (_15176_, _15122_, _03327_);
  or (_15177_, _15176_, _07431_);
  or (_15178_, _15177_, _15175_);
  or (_15179_, _15178_, _15170_);
  and (_15180_, _15179_, _15143_);
  or (_15181_, _15180_, _03413_);
  or (_15182_, _05847_, _03849_);
  and (_15183_, _15182_, _02959_);
  and (_15185_, _15183_, _15181_);
  nor (_15186_, _07610_, _02959_);
  or (_15187_, _15186_, _07497_);
  or (_15188_, _15187_, _15185_);
  nand (_15189_, _07497_, _06984_);
  and (_15190_, _15189_, _15188_);
  or (_15191_, _15190_, _02887_);
  and (_15192_, _11675_, _05331_);
  nor (_15193_, _15192_, _15171_);
  nand (_15194_, _15193_, _02887_);
  and (_15196_, _15194_, _02881_);
  and (_15197_, _15196_, _15191_);
  and (_15198_, _15172_, _11682_);
  nor (_15199_, _15198_, _15171_);
  nor (_15200_, _15199_, _02881_);
  or (_15201_, _15200_, _06271_);
  or (_15202_, _15201_, _15197_);
  nor (_15203_, _06748_, _06746_);
  nor (_15204_, _15203_, _06749_);
  or (_15205_, _15204_, _06277_);
  and (_15207_, _15205_, _15202_);
  or (_15208_, _15207_, _07427_);
  nand (_15209_, _04896_, \oc8051_golden_model_1.ACC [5]);
  nor (_15210_, _04896_, \oc8051_golden_model_1.ACC [5]);
  or (_15211_, _14883_, _15210_);
  and (_15212_, _15211_, _15209_);
  nor (_15213_, _15212_, _07223_);
  and (_15214_, _15212_, _07223_);
  nor (_15215_, _15214_, _15213_);
  nor (_15216_, _14893_, _14887_);
  and (_15218_, _15216_, \oc8051_golden_model_1.PSW [7]);
  or (_15219_, _15218_, _15215_);
  nand (_15220_, _15218_, _15215_);
  and (_15221_, _15220_, _15219_);
  or (_15222_, _15221_, _07426_);
  and (_15223_, _15222_, _07344_);
  and (_15224_, _15223_, _15208_);
  or (_15225_, _15224_, _02992_);
  or (_15226_, _15225_, _15142_);
  and (_15227_, _15226_, _15127_);
  nor (_15229_, _14804_, _10014_);
  nor (_15230_, _15229_, _10013_);
  nor (_15231_, _15230_, _08139_);
  and (_15232_, _15230_, _08139_);
  nor (_15233_, _15232_, _15231_);
  nor (_15234_, _14814_, _14808_);
  and (_15235_, _15234_, \oc8051_golden_model_1.PSW [7]);
  nor (_15236_, _15235_, _15233_);
  and (_15237_, _15235_, _15233_);
  nor (_15238_, _15237_, _15236_);
  and (_15240_, _15238_, _07276_);
  or (_15241_, _15240_, _02585_);
  or (_15242_, _15241_, _15227_);
  nand (_15243_, _02932_, _02585_);
  and (_15244_, _15243_, _02875_);
  and (_15245_, _15244_, _15242_);
  nor (_15246_, _11650_, _07755_);
  nor (_15247_, _15246_, _15171_);
  nor (_15248_, _15247_, _02875_);
  or (_15249_, _15248_, _06793_);
  or (_15251_, _15249_, _15245_);
  and (_15252_, _15251_, _15123_);
  or (_15253_, _15252_, _02855_);
  and (_15254_, _05847_, _04712_);
  nor (_15255_, _15254_, _15111_);
  nand (_15256_, _15255_, _02855_);
  and (_15257_, _15256_, _02851_);
  and (_15258_, _15257_, _15253_);
  nor (_15259_, _11751_, _07272_);
  nor (_15260_, _15259_, _15111_);
  nor (_15262_, _15260_, _02851_);
  or (_15263_, _15262_, _06807_);
  or (_15264_, _15263_, _15258_);
  not (_15265_, _06834_);
  and (_15266_, _06837_, _15265_);
  or (_15267_, _15266_, _06813_);
  and (_15268_, _15267_, _15264_);
  and (_15269_, _15268_, _02584_);
  nor (_15270_, _02932_, _02584_);
  or (_15271_, _15270_, _03014_);
  or (_15273_, _15271_, _15269_);
  and (_15274_, _11758_, _04712_);
  nor (_15275_, _15274_, _15111_);
  nand (_15276_, _15275_, _03014_);
  and (_15277_, _15276_, _07783_);
  and (_15278_, _15277_, _15273_);
  nor (_15279_, _07783_, _02932_);
  or (_15280_, _15279_, _15117_);
  or (_15281_, _15280_, _15278_);
  nand (_15282_, _15281_, _15120_);
  and (_15284_, _05318_, _02511_);
  nor (_15285_, _15284_, _15282_);
  and (_15286_, _15284_, _07223_);
  nor (_15287_, _15286_, _15285_);
  nor (_15288_, _15287_, _15116_);
  or (_15289_, _07223_, _02498_);
  and (_15290_, _15289_, _15115_);
  or (_15291_, _15290_, _15288_);
  nand (_15292_, _15119_, _07794_);
  and (_15293_, _15292_, _14650_);
  and (_15295_, _15293_, _15291_);
  and (_15296_, _14649_, _08067_);
  or (_15297_, _15296_, _15295_);
  and (_15298_, _15297_, _14491_);
  and (_15299_, _08067_, _03504_);
  or (_15300_, _15299_, _03132_);
  or (_15301_, _15300_, _15298_);
  or (_15302_, _11769_, _07814_);
  and (_15303_, _15302_, _07813_);
  and (_15304_, _15303_, _15301_);
  and (_15306_, _07812_, _08139_);
  or (_15307_, _15306_, _03021_);
  or (_15308_, _15307_, _15304_);
  and (_15309_, _15308_, _15114_);
  or (_15310_, _15309_, _03130_);
  or (_15311_, _15111_, _03131_);
  and (_15312_, _15311_, _07828_);
  and (_15313_, _15312_, _15310_);
  or (_15314_, _15313_, _15110_);
  and (_15315_, _15314_, _07265_);
  and (_15317_, _08065_, _03513_);
  or (_15318_, _15317_, _03141_);
  or (_15319_, _15318_, _15315_);
  and (_15320_, _15319_, _15109_);
  and (_15321_, _07836_, _08137_);
  or (_15322_, _15321_, _15320_);
  and (_15323_, _15322_, _05274_);
  or (_15324_, _15275_, _11768_);
  or (_15325_, _15324_, _05274_);
  nand (_15326_, _15325_, _08871_);
  or (_15328_, _15326_, _15323_);
  not (_15329_, _08870_);
  nor (_15330_, _15329_, _07222_);
  or (_15331_, _15330_, _08872_);
  and (_15332_, _15331_, _15328_);
  nor (_15333_, _08870_, _07222_);
  or (_15334_, _15333_, _07858_);
  or (_15335_, _15334_, _15332_);
  nand (_15336_, _08066_, _07858_);
  and (_15337_, _15336_, _03126_);
  and (_15339_, _15337_, _15335_);
  nand (_15340_, _11768_, _07868_);
  and (_15341_, _15340_, _07867_);
  or (_15342_, _15341_, _15339_);
  and (_15343_, _15342_, _15106_);
  or (_15344_, _15343_, _03036_);
  nor (_15345_, _11644_, _07272_);
  nor (_15346_, _15345_, _15111_);
  nand (_15347_, _15346_, _03036_);
  and (_15348_, _15347_, _07889_);
  and (_15350_, _15348_, _15344_);
  and (_15351_, _07908_, _07891_);
  nor (_15352_, _15351_, _07909_);
  and (_15353_, _15352_, _10171_);
  or (_15354_, _15353_, _15350_);
  and (_15355_, _15354_, _07922_);
  and (_15356_, _07941_, _07924_);
  nor (_15357_, _15356_, _07942_);
  and (_15358_, _15357_, _07917_);
  or (_15359_, _15358_, _15355_);
  and (_15361_, _15359_, _03138_);
  or (_15362_, _15361_, _15105_);
  and (_15363_, _15362_, _08031_);
  and (_15364_, _08050_, _07293_);
  nor (_15365_, _15364_, _08051_);
  and (_15366_, _15365_, _07950_);
  or (_15367_, _15366_, _08029_);
  or (_15368_, _15367_, _15363_);
  nand (_15369_, _08029_, _06879_);
  and (_15370_, _15369_, _07259_);
  and (_15372_, _15370_, _15368_);
  nor (_15373_, _07252_, _07223_);
  nor (_15374_, _15373_, _07253_);
  or (_15375_, _15374_, _07217_);
  and (_15376_, _15375_, _09524_);
  or (_15377_, _15376_, _15372_);
  nor (_15378_, _08094_, _08067_);
  nor (_15379_, _15378_, _08095_);
  or (_15380_, _15379_, _08064_);
  and (_15381_, _15380_, _02901_);
  and (_15383_, _15381_, _15377_);
  and (_15384_, _08126_, _07613_);
  nor (_15385_, _15384_, _08127_);
  or (_15386_, _15385_, _08103_);
  and (_15387_, _15386_, _08105_);
  or (_15388_, _15387_, _15383_);
  nor (_15389_, _08167_, _08139_);
  nor (_15390_, _15389_, _08168_);
  or (_15391_, _15390_, _08106_);
  and (_15392_, _15391_, _08136_);
  and (_15394_, _15392_, _15388_);
  and (_15395_, _08135_, \oc8051_golden_model_1.ACC [5]);
  or (_15396_, _15395_, _03166_);
  or (_15397_, _15396_, _15394_);
  nand (_15398_, _15159_, _03166_);
  and (_15399_, _15398_, _08180_);
  and (_15400_, _15399_, _15397_);
  nor (_15401_, _08187_, _06833_);
  or (_15402_, _15401_, _08188_);
  and (_15403_, _15402_, _08179_);
  or (_15405_, _15403_, _08184_);
  or (_15406_, _15405_, _15400_);
  nand (_15407_, _08184_, _05768_);
  and (_15408_, _15407_, _02501_);
  and (_15409_, _15408_, _15406_);
  nor (_15410_, _15193_, _02501_);
  or (_15411_, _15410_, _03174_);
  or (_15412_, _15411_, _15409_);
  and (_15413_, _11821_, _04712_);
  nor (_15414_, _15413_, _15111_);
  nand (_15416_, _15414_, _03174_);
  and (_15417_, _15416_, _08202_);
  and (_15418_, _15417_, _15412_);
  nor (_15419_, _08212_, \oc8051_golden_model_1.ACC [6]);
  nor (_15420_, _15419_, _08213_);
  and (_15421_, _15420_, _08201_);
  or (_15422_, _15421_, _08208_);
  or (_15423_, _15422_, _15418_);
  nand (_15424_, _08208_, _05768_);
  and (_15425_, _15424_, _34698_);
  and (_15427_, _15425_, _15423_);
  or (_15428_, _15427_, _15102_);
  and (_35170_, _15428_, _36029_);
  not (_15429_, \oc8051_golden_model_1.DPL [0]);
  nor (_15430_, _34698_, _15429_);
  and (_15431_, _05044_, _04654_);
  nor (_15432_, _04654_, _15429_);
  and (_15433_, _04654_, _05566_);
  or (_15434_, _15433_, _15432_);
  nand (_15435_, _15434_, _03020_);
  nor (_15437_, _15435_, _15431_);
  and (_15438_, _04654_, _03817_);
  or (_15439_, _15438_, _15432_);
  or (_15440_, _15439_, _06241_);
  and (_15441_, _04654_, \oc8051_golden_model_1.ACC [0]);
  or (_15442_, _15441_, _15432_);
  or (_15443_, _15442_, _02959_);
  or (_15444_, _15432_, _15431_);
  or (_15445_, _15444_, _03821_);
  and (_15446_, _15442_, _03825_);
  nor (_15448_, _03825_, _15429_);
  or (_15449_, _15448_, _02952_);
  or (_15450_, _15449_, _15446_);
  and (_15451_, _15450_, _03327_);
  and (_15452_, _15451_, _15445_);
  and (_15453_, _15439_, _02947_);
  or (_15454_, _15453_, _02950_);
  or (_15455_, _15454_, _15452_);
  and (_15456_, _15455_, _15443_);
  or (_15457_, _15456_, _08250_);
  nand (_15459_, _08250_, \oc8051_golden_model_1.DPL [0]);
  and (_15460_, _15459_, _08235_);
  and (_15461_, _15460_, _15457_);
  nor (_15462_, _03492_, _08235_);
  or (_15463_, _15462_, _06793_);
  or (_15464_, _15463_, _15461_);
  and (_15465_, _15464_, _15440_);
  or (_15466_, _15465_, _02855_);
  and (_15467_, _06174_, _04654_);
  or (_15468_, _15432_, _02856_);
  or (_15470_, _15468_, _15467_);
  and (_15471_, _15470_, _15466_);
  or (_15472_, _15471_, _02576_);
  nor (_15473_, _10530_, _08231_);
  or (_15474_, _15432_, _02851_);
  or (_15475_, _15474_, _15473_);
  and (_15476_, _15475_, _03884_);
  and (_15477_, _15476_, _15472_);
  and (_15478_, _15434_, _03014_);
  or (_15479_, _15478_, _03021_);
  or (_15481_, _15479_, _15477_);
  and (_15482_, _10425_, _04654_);
  or (_15483_, _15482_, _15432_);
  or (_15484_, _15483_, _05279_);
  and (_15485_, _15484_, _15481_);
  or (_15486_, _15485_, _03130_);
  and (_15487_, _10546_, _04654_);
  or (_15488_, _15432_, _03131_);
  or (_15489_, _15488_, _15487_);
  and (_15490_, _15489_, _05274_);
  and (_15492_, _15490_, _15486_);
  or (_15493_, _15492_, _15437_);
  and (_15494_, _15493_, _03140_);
  or (_15495_, _15432_, _09183_);
  and (_15496_, _15442_, _03139_);
  and (_15497_, _15496_, _15495_);
  or (_15498_, _15497_, _03036_);
  or (_15499_, _15498_, _15494_);
  nor (_15500_, _10423_, _08231_);
  or (_15501_, _15432_, _05781_);
  or (_15503_, _15501_, _15500_);
  and (_15504_, _15503_, _05786_);
  and (_15505_, _15504_, _15499_);
  not (_15506_, _03265_);
  nor (_15507_, _10421_, _08231_);
  or (_15508_, _15507_, _15432_);
  and (_15509_, _15508_, _03127_);
  or (_15510_, _15509_, _15506_);
  or (_15511_, _15510_, _15505_);
  or (_15512_, _15444_, _03265_);
  and (_15514_, _15512_, _34698_);
  and (_15515_, _15514_, _15511_);
  or (_15516_, _15515_, _15430_);
  and (_35172_, _15516_, _36029_);
  not (_15517_, \oc8051_golden_model_1.DPL [1]);
  nor (_15518_, _34698_, _15517_);
  or (_15519_, _10739_, _08231_);
  or (_15520_, _04654_, \oc8051_golden_model_1.DPL [1]);
  and (_15521_, _15520_, _03130_);
  and (_15522_, _15521_, _15519_);
  nand (_15524_, _10720_, _04654_);
  and (_15525_, _15520_, _02576_);
  and (_15526_, _15525_, _15524_);
  nor (_15527_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_15528_, _15527_, _08255_);
  and (_15529_, _15528_, _08250_);
  and (_15530_, _10622_, _04654_);
  not (_15531_, _15530_);
  and (_15532_, _15531_, _15520_);
  or (_15533_, _15532_, _03821_);
  nand (_15535_, _04654_, _02618_);
  and (_15536_, _15535_, _15520_);
  and (_15537_, _15536_, _03825_);
  nor (_15538_, _03825_, _15517_);
  or (_15539_, _15538_, _02952_);
  or (_15540_, _15539_, _15537_);
  and (_15541_, _15540_, _03327_);
  and (_15542_, _15541_, _15533_);
  nor (_15543_, _04654_, _15517_);
  and (_15544_, _04654_, _04005_);
  or (_15546_, _15544_, _15543_);
  and (_15547_, _15546_, _02947_);
  or (_15548_, _15547_, _02950_);
  or (_15549_, _15548_, _15542_);
  or (_15550_, _15536_, _02959_);
  and (_15551_, _15550_, _08251_);
  and (_15552_, _15551_, _15549_);
  or (_15553_, _15552_, _15529_);
  and (_15554_, _15553_, _08235_);
  nor (_15555_, _03705_, _08235_);
  or (_15557_, _15555_, _06793_);
  or (_15558_, _15557_, _15554_);
  or (_15559_, _15546_, _06241_);
  and (_15560_, _15559_, _15558_);
  or (_15561_, _15560_, _02855_);
  and (_15562_, _06173_, _04654_);
  or (_15563_, _15543_, _02856_);
  or (_15564_, _15563_, _15562_);
  and (_15565_, _15564_, _02851_);
  and (_15566_, _15565_, _15561_);
  or (_15568_, _15566_, _15526_);
  and (_15569_, _15568_, _03884_);
  nand (_15570_, _04654_, _03705_);
  and (_15571_, _15520_, _03014_);
  and (_15572_, _15571_, _15570_);
  or (_15573_, _15572_, _15569_);
  and (_15574_, _15573_, _05279_);
  or (_15575_, _10612_, _08231_);
  and (_15576_, _15520_, _03021_);
  and (_15577_, _15576_, _15575_);
  or (_15579_, _15577_, _15574_);
  and (_15580_, _15579_, _03131_);
  or (_15581_, _15580_, _15522_);
  and (_15582_, _15581_, _05274_);
  or (_15583_, _10611_, _08231_);
  and (_15584_, _15520_, _03020_);
  and (_15585_, _15584_, _15583_);
  or (_15586_, _15585_, _15582_);
  and (_15587_, _15586_, _03140_);
  or (_15588_, _15543_, _12724_);
  and (_15590_, _15536_, _03139_);
  and (_15591_, _15590_, _15588_);
  or (_15592_, _15591_, _15587_);
  and (_15593_, _15592_, _03128_);
  or (_15594_, _15535_, _12724_);
  and (_15595_, _15520_, _03127_);
  and (_15596_, _15595_, _15594_);
  or (_15597_, _15596_, _03166_);
  or (_15598_, _15570_, _12724_);
  and (_15599_, _15520_, _03036_);
  and (_15601_, _15599_, _15598_);
  or (_15602_, _15601_, _15597_);
  or (_15603_, _15602_, _15593_);
  or (_15604_, _15532_, _03563_);
  and (_15605_, _15604_, _15603_);
  or (_15606_, _15605_, _03174_);
  or (_15607_, _15543_, _03178_);
  or (_15608_, _15607_, _15530_);
  and (_15609_, _15608_, _34698_);
  and (_15610_, _15609_, _15606_);
  or (_15612_, _15610_, _15518_);
  and (_35173_, _15612_, _36029_);
  not (_15613_, \oc8051_golden_model_1.DPL [2]);
  nor (_15614_, _34698_, _15613_);
  nor (_15615_, _04654_, _15613_);
  nor (_15616_, _10830_, _08231_);
  or (_15617_, _15616_, _15615_);
  and (_15618_, _15617_, _03127_);
  or (_15619_, _15615_, _05143_);
  and (_15620_, _04654_, _05727_);
  or (_15622_, _15620_, _15615_);
  and (_15623_, _15622_, _03020_);
  and (_15624_, _15623_, _15619_);
  and (_15625_, _10831_, _04654_);
  or (_15626_, _15625_, _15615_);
  and (_15627_, _15626_, _03130_);
  nor (_15628_, _08231_, _04440_);
  or (_15629_, _15628_, _15615_);
  or (_15630_, _15629_, _06241_);
  nor (_15631_, _10849_, _08231_);
  or (_15633_, _15631_, _15615_);
  or (_15634_, _15633_, _03821_);
  and (_15635_, _04654_, \oc8051_golden_model_1.ACC [2]);
  or (_15636_, _15635_, _15615_);
  and (_15637_, _15636_, _03825_);
  nor (_15638_, _03825_, _15613_);
  or (_15639_, _15638_, _02952_);
  or (_15640_, _15639_, _15637_);
  and (_15641_, _15640_, _03327_);
  and (_15642_, _15641_, _15634_);
  and (_15644_, _15629_, _02947_);
  or (_15645_, _15644_, _02950_);
  or (_15646_, _15645_, _15642_);
  or (_15647_, _15636_, _02959_);
  and (_15648_, _15647_, _08251_);
  and (_15649_, _15648_, _15646_);
  nor (_15650_, _08255_, \oc8051_golden_model_1.DPL [2]);
  nor (_15651_, _15650_, _08256_);
  and (_15652_, _15651_, _08250_);
  or (_15653_, _15652_, _15649_);
  and (_15655_, _15653_, _08235_);
  nor (_15656_, _03302_, _08235_);
  or (_15657_, _15656_, _06793_);
  or (_15658_, _15657_, _15655_);
  and (_15659_, _15658_, _15630_);
  or (_15660_, _15659_, _02855_);
  and (_15661_, _06177_, _04654_);
  or (_15662_, _15615_, _02856_);
  or (_15663_, _15662_, _15661_);
  and (_15664_, _15663_, _02851_);
  and (_15666_, _15664_, _15660_);
  nor (_15667_, _10943_, _08231_);
  or (_15668_, _15667_, _15615_);
  and (_15669_, _15668_, _02576_);
  or (_15670_, _15669_, _03014_);
  or (_15671_, _15670_, _15666_);
  or (_15672_, _15622_, _03884_);
  and (_15673_, _15672_, _15671_);
  or (_15674_, _15673_, _03021_);
  and (_15675_, _10835_, _04654_);
  or (_15677_, _15615_, _05279_);
  or (_15678_, _15677_, _15675_);
  and (_15679_, _15678_, _03131_);
  and (_15680_, _15679_, _15674_);
  or (_15681_, _15680_, _15627_);
  and (_15682_, _15681_, _05274_);
  or (_15683_, _15682_, _15624_);
  and (_15684_, _15683_, _03140_);
  and (_15685_, _15636_, _03139_);
  and (_15686_, _15685_, _15619_);
  or (_15688_, _15686_, _03036_);
  or (_15689_, _15688_, _15684_);
  nor (_15690_, _10833_, _08231_);
  or (_15691_, _15615_, _05781_);
  or (_15692_, _15691_, _15690_);
  and (_15693_, _15692_, _05786_);
  and (_15694_, _15693_, _15689_);
  or (_15695_, _15694_, _15618_);
  and (_15696_, _15695_, _03563_);
  and (_15697_, _15633_, _03166_);
  or (_15699_, _15697_, _03174_);
  or (_15700_, _15699_, _15696_);
  and (_15701_, _11008_, _04654_);
  or (_15702_, _15615_, _03178_);
  or (_15703_, _15702_, _15701_);
  and (_15704_, _15703_, _34698_);
  and (_15705_, _15704_, _15700_);
  or (_15706_, _15705_, _15614_);
  and (_35174_, _15706_, _36029_);
  or (_15707_, _34698_, \oc8051_golden_model_1.DPL [3]);
  and (_15709_, _15707_, _36029_);
  and (_15710_, _08231_, \oc8051_golden_model_1.DPL [3]);
  and (_15711_, _11028_, _04654_);
  or (_15712_, _15711_, _15710_);
  and (_15713_, _15712_, _03130_);
  nor (_15714_, _08231_, _04242_);
  or (_15715_, _15714_, _15710_);
  or (_15716_, _15715_, _06241_);
  nor (_15717_, _08256_, \oc8051_golden_model_1.DPL [3]);
  nor (_15718_, _15717_, _08257_);
  and (_15720_, _15718_, _08250_);
  nor (_15721_, _11040_, _08231_);
  or (_15722_, _15721_, _15710_);
  or (_15723_, _15722_, _03821_);
  and (_15724_, _04654_, \oc8051_golden_model_1.ACC [3]);
  or (_15725_, _15724_, _15710_);
  and (_15726_, _15725_, _03825_);
  and (_15727_, _03826_, \oc8051_golden_model_1.DPL [3]);
  or (_15728_, _15727_, _02952_);
  or (_15729_, _15728_, _15726_);
  and (_15731_, _15729_, _03327_);
  and (_15732_, _15731_, _15723_);
  and (_15733_, _15715_, _02947_);
  or (_15734_, _15733_, _02950_);
  or (_15735_, _15734_, _15732_);
  or (_15736_, _15725_, _02959_);
  and (_15737_, _15736_, _08251_);
  and (_15738_, _15737_, _15735_);
  or (_15739_, _15738_, _15720_);
  and (_15740_, _15739_, _08235_);
  nor (_15742_, _03120_, _08235_);
  or (_15743_, _15742_, _06793_);
  or (_15744_, _15743_, _15740_);
  and (_15745_, _15744_, _15716_);
  or (_15746_, _15745_, _02855_);
  and (_15747_, _06176_, _04654_);
  or (_15748_, _15710_, _02856_);
  or (_15749_, _15748_, _15747_);
  and (_15750_, _15749_, _02851_);
  and (_15751_, _15750_, _15746_);
  nor (_15753_, _11143_, _08231_);
  or (_15754_, _15753_, _15710_);
  and (_15755_, _15754_, _02576_);
  or (_15756_, _15755_, _03014_);
  or (_15757_, _15756_, _15751_);
  and (_15758_, _04654_, _05664_);
  or (_15759_, _15758_, _15710_);
  or (_15760_, _15759_, _03884_);
  and (_15761_, _15760_, _15757_);
  or (_15762_, _15761_, _03021_);
  and (_15764_, _11032_, _04654_);
  or (_15765_, _15710_, _05279_);
  or (_15766_, _15765_, _15764_);
  and (_15767_, _15766_, _03131_);
  and (_15768_, _15767_, _15762_);
  or (_15769_, _15768_, _15713_);
  and (_15770_, _15769_, _05274_);
  or (_15771_, _15710_, _04996_);
  and (_15772_, _15759_, _03020_);
  and (_15773_, _15772_, _15771_);
  or (_15775_, _15773_, _15770_);
  and (_15776_, _15775_, _03140_);
  and (_15777_, _15725_, _03139_);
  and (_15778_, _15777_, _15771_);
  or (_15779_, _15778_, _03036_);
  or (_15780_, _15779_, _15776_);
  nor (_15781_, _11030_, _08231_);
  or (_15782_, _15710_, _05781_);
  or (_15783_, _15782_, _15781_);
  and (_15784_, _15783_, _05786_);
  and (_15786_, _15784_, _15780_);
  nor (_15787_, _11027_, _08231_);
  or (_15788_, _15787_, _15710_);
  and (_15789_, _15788_, _03127_);
  or (_15790_, _15789_, _03166_);
  or (_15791_, _15790_, _15786_);
  or (_15792_, _15722_, _03563_);
  and (_15793_, _15792_, _03178_);
  and (_15794_, _15793_, _15791_);
  and (_15795_, _11213_, _04654_);
  or (_15797_, _15795_, _15710_);
  and (_15798_, _15797_, _03174_);
  or (_15799_, _15798_, _34702_);
  or (_15800_, _15799_, _15794_);
  and (_35175_, _15800_, _15709_);
  or (_15801_, _34698_, \oc8051_golden_model_1.DPL [4]);
  and (_15802_, _15801_, _36029_);
  and (_15803_, _08231_, \oc8051_golden_model_1.DPL [4]);
  and (_15804_, _11368_, _04654_);
  or (_15805_, _15804_, _15803_);
  and (_15807_, _15805_, _03130_);
  nor (_15808_, _05202_, _08231_);
  or (_15809_, _15808_, _15803_);
  or (_15810_, _15809_, _06241_);
  nor (_15811_, _11259_, _08231_);
  or (_15812_, _15811_, _15803_);
  or (_15813_, _15812_, _03821_);
  and (_15814_, _04654_, \oc8051_golden_model_1.ACC [4]);
  or (_15815_, _15814_, _15803_);
  and (_15816_, _15815_, _03825_);
  and (_15818_, _03826_, \oc8051_golden_model_1.DPL [4]);
  or (_15819_, _15818_, _02952_);
  or (_15820_, _15819_, _15816_);
  and (_15821_, _15820_, _03327_);
  and (_15822_, _15821_, _15813_);
  and (_15823_, _15809_, _02947_);
  or (_15824_, _15823_, _02950_);
  or (_15825_, _15824_, _15822_);
  or (_15826_, _15815_, _02959_);
  and (_15827_, _15826_, _08251_);
  and (_15829_, _15827_, _15825_);
  nor (_15830_, _08257_, \oc8051_golden_model_1.DPL [4]);
  nor (_15831_, _15830_, _08258_);
  and (_15832_, _15831_, _08250_);
  or (_15833_, _15832_, _15829_);
  and (_15834_, _15833_, _08235_);
  nor (_15835_, _05630_, _08235_);
  or (_15836_, _15835_, _06793_);
  or (_15837_, _15836_, _15834_);
  and (_15838_, _15837_, _15810_);
  or (_15840_, _15838_, _02855_);
  and (_15841_, _06181_, _04654_);
  or (_15842_, _15803_, _02856_);
  or (_15843_, _15842_, _15841_);
  and (_15844_, _15843_, _02851_);
  and (_15845_, _15844_, _15840_);
  nor (_15846_, _11348_, _08231_);
  or (_15847_, _15846_, _15803_);
  and (_15848_, _15847_, _02576_);
  or (_15849_, _15848_, _03014_);
  or (_15851_, _15849_, _15845_);
  and (_15852_, _05697_, _04654_);
  or (_15853_, _15852_, _15803_);
  or (_15854_, _15853_, _03884_);
  and (_15855_, _15854_, _15851_);
  or (_15856_, _15855_, _03021_);
  and (_15857_, _11362_, _04654_);
  or (_15858_, _15803_, _05279_);
  or (_15859_, _15858_, _15857_);
  and (_15860_, _15859_, _03131_);
  and (_15862_, _15860_, _15856_);
  or (_15863_, _15862_, _15807_);
  and (_15864_, _15863_, _05274_);
  or (_15865_, _15803_, _05251_);
  and (_15866_, _15853_, _03020_);
  and (_15867_, _15866_, _15865_);
  or (_15868_, _15867_, _15864_);
  and (_15869_, _15868_, _03140_);
  and (_15870_, _15815_, _03139_);
  and (_15871_, _15870_, _15865_);
  or (_15873_, _15871_, _03036_);
  or (_15874_, _15873_, _15869_);
  nor (_15875_, _11361_, _08231_);
  or (_15876_, _15803_, _05781_);
  or (_15877_, _15876_, _15875_);
  and (_15878_, _15877_, _05786_);
  and (_15879_, _15878_, _15874_);
  nor (_15880_, _11367_, _08231_);
  or (_15881_, _15880_, _15803_);
  and (_15882_, _15881_, _03127_);
  or (_15884_, _15882_, _03166_);
  or (_15885_, _15884_, _15879_);
  or (_15886_, _15812_, _03563_);
  and (_15887_, _15886_, _03178_);
  and (_15888_, _15887_, _15885_);
  and (_15889_, _11417_, _04654_);
  or (_15890_, _15889_, _15803_);
  and (_15891_, _15890_, _03174_);
  or (_15892_, _15891_, _34702_);
  or (_15893_, _15892_, _15888_);
  and (_35176_, _15893_, _15802_);
  or (_15895_, _34698_, \oc8051_golden_model_1.DPL [5]);
  and (_15896_, _15895_, _36029_);
  and (_15897_, _08231_, \oc8051_golden_model_1.DPL [5]);
  and (_15898_, _11436_, _04654_);
  or (_15899_, _15898_, _15897_);
  and (_15900_, _15899_, _03130_);
  nor (_15901_, _04896_, _08231_);
  or (_15902_, _15901_, _15897_);
  or (_15903_, _15902_, _06241_);
  nor (_15905_, _11445_, _08231_);
  or (_15906_, _15905_, _15897_);
  or (_15907_, _15906_, _03821_);
  and (_15908_, _04654_, \oc8051_golden_model_1.ACC [5]);
  or (_15909_, _15908_, _15897_);
  and (_15910_, _15909_, _03825_);
  and (_15911_, _03826_, \oc8051_golden_model_1.DPL [5]);
  or (_15912_, _15911_, _02952_);
  or (_15913_, _15912_, _15910_);
  and (_15914_, _15913_, _03327_);
  and (_15916_, _15914_, _15907_);
  and (_15917_, _15902_, _02947_);
  or (_15918_, _15917_, _02950_);
  or (_15919_, _15918_, _15916_);
  or (_15920_, _15909_, _02959_);
  and (_15921_, _15920_, _08251_);
  and (_15922_, _15921_, _15919_);
  nor (_15923_, _08258_, \oc8051_golden_model_1.DPL [5]);
  nor (_15924_, _15923_, _08259_);
  and (_15925_, _15924_, _08250_);
  or (_15927_, _15925_, _15922_);
  and (_15928_, _15927_, _08235_);
  nor (_15929_, _05661_, _08235_);
  or (_15930_, _15929_, _06793_);
  or (_15931_, _15930_, _15928_);
  and (_15932_, _15931_, _15903_);
  or (_15933_, _15932_, _02855_);
  and (_15934_, _06180_, _04654_);
  or (_15935_, _15897_, _02856_);
  or (_15936_, _15935_, _15934_);
  and (_15938_, _15936_, _02851_);
  and (_15939_, _15938_, _15933_);
  nor (_15940_, _11546_, _08231_);
  or (_15941_, _15940_, _15897_);
  and (_15942_, _15941_, _02576_);
  or (_15943_, _15942_, _03014_);
  or (_15944_, _15943_, _15939_);
  and (_15945_, _05701_, _04654_);
  or (_15946_, _15945_, _15897_);
  or (_15947_, _15946_, _03884_);
  and (_15949_, _15947_, _15944_);
  or (_15950_, _15949_, _03021_);
  and (_15951_, _11562_, _04654_);
  or (_15952_, _15897_, _05279_);
  or (_15953_, _15952_, _15951_);
  and (_15954_, _15953_, _03131_);
  and (_15955_, _15954_, _15950_);
  or (_15956_, _15955_, _15900_);
  and (_15957_, _15956_, _05274_);
  or (_15958_, _15897_, _04944_);
  and (_15960_, _15946_, _03020_);
  and (_15961_, _15960_, _15958_);
  or (_15962_, _15961_, _15957_);
  and (_15963_, _15962_, _03140_);
  and (_15964_, _15909_, _03139_);
  and (_15965_, _15964_, _15958_);
  or (_15966_, _15965_, _03036_);
  or (_15967_, _15966_, _15963_);
  nor (_15968_, _11560_, _08231_);
  or (_15969_, _15897_, _05781_);
  or (_15971_, _15969_, _15968_);
  and (_15972_, _15971_, _05786_);
  and (_15973_, _15972_, _15967_);
  nor (_15974_, _11435_, _08231_);
  or (_15975_, _15974_, _15897_);
  and (_15976_, _15975_, _03127_);
  or (_15977_, _15976_, _03166_);
  or (_15978_, _15977_, _15973_);
  or (_15979_, _15906_, _03563_);
  and (_15980_, _15979_, _03178_);
  and (_15982_, _15980_, _15978_);
  and (_15983_, _11619_, _04654_);
  or (_15984_, _15983_, _15897_);
  and (_15985_, _15984_, _03174_);
  or (_15986_, _15985_, _34702_);
  or (_15987_, _15986_, _15982_);
  and (_35178_, _15987_, _15896_);
  or (_15988_, _34698_, \oc8051_golden_model_1.DPL [6]);
  and (_15989_, _15988_, _36029_);
  not (_15990_, \oc8051_golden_model_1.DPL [6]);
  nor (_15992_, _04654_, _15990_);
  and (_15993_, _11769_, _04654_);
  or (_15994_, _15993_, _15992_);
  and (_15995_, _15994_, _03130_);
  nor (_15996_, _04787_, _08231_);
  or (_15997_, _15996_, _15992_);
  or (_15998_, _15997_, _06241_);
  nor (_15999_, _11636_, _08231_);
  or (_16000_, _15999_, _15992_);
  or (_16001_, _16000_, _03821_);
  and (_16003_, _04654_, \oc8051_golden_model_1.ACC [6]);
  or (_16004_, _16003_, _15992_);
  and (_16005_, _16004_, _03825_);
  nor (_16006_, _03825_, _15990_);
  or (_16007_, _16006_, _02952_);
  or (_16008_, _16007_, _16005_);
  and (_16009_, _16008_, _03327_);
  and (_16010_, _16009_, _16001_);
  and (_16011_, _15997_, _02947_);
  or (_16012_, _16011_, _02950_);
  or (_16014_, _16012_, _16010_);
  or (_16015_, _16004_, _02959_);
  and (_16016_, _16015_, _08251_);
  and (_16017_, _16016_, _16014_);
  nor (_16018_, _08259_, \oc8051_golden_model_1.DPL [6]);
  nor (_16019_, _16018_, _08260_);
  and (_16020_, _16019_, _08250_);
  or (_16021_, _16020_, _16017_);
  and (_16022_, _16021_, _08235_);
  nor (_16023_, _05598_, _08235_);
  or (_16025_, _16023_, _06793_);
  or (_16026_, _16025_, _16022_);
  and (_16027_, _16026_, _15998_);
  or (_16028_, _16027_, _02855_);
  and (_16029_, _05847_, _04654_);
  or (_16030_, _15992_, _02856_);
  or (_16031_, _16030_, _16029_);
  and (_16032_, _16031_, _02851_);
  and (_16033_, _16032_, _16028_);
  nor (_16034_, _11751_, _08231_);
  or (_16036_, _16034_, _15992_);
  and (_16037_, _16036_, _02576_);
  or (_16038_, _16037_, _03014_);
  or (_16039_, _16038_, _16033_);
  and (_16040_, _11758_, _04654_);
  or (_16041_, _16040_, _15992_);
  or (_16042_, _16041_, _03884_);
  and (_16043_, _16042_, _16039_);
  or (_16044_, _16043_, _03021_);
  and (_16045_, _11646_, _04654_);
  or (_16047_, _15992_, _05279_);
  or (_16048_, _16047_, _16045_);
  and (_16049_, _16048_, _03131_);
  and (_16050_, _16049_, _16044_);
  or (_16051_, _16050_, _15995_);
  and (_16052_, _16051_, _05274_);
  or (_16053_, _15992_, _04838_);
  and (_16054_, _16041_, _03020_);
  and (_16055_, _16054_, _16053_);
  or (_16056_, _16055_, _16052_);
  and (_16058_, _16056_, _03140_);
  and (_16059_, _16004_, _03139_);
  and (_16060_, _16059_, _16053_);
  or (_16061_, _16060_, _03036_);
  or (_16062_, _16061_, _16058_);
  nor (_16063_, _11644_, _08231_);
  or (_16064_, _15992_, _05781_);
  or (_16065_, _16064_, _16063_);
  and (_16066_, _16065_, _05786_);
  and (_16067_, _16066_, _16062_);
  nor (_16069_, _11768_, _08231_);
  or (_16070_, _16069_, _15992_);
  and (_16071_, _16070_, _03127_);
  or (_16072_, _16071_, _03166_);
  or (_16073_, _16072_, _16067_);
  or (_16074_, _16000_, _03563_);
  and (_16075_, _16074_, _03178_);
  and (_16076_, _16075_, _16073_);
  and (_16077_, _11821_, _04654_);
  or (_16078_, _16077_, _15992_);
  and (_16080_, _16078_, _03174_);
  or (_16081_, _16080_, _34702_);
  or (_16082_, _16081_, _16076_);
  and (_35179_, _16082_, _15989_);
  nor (_16083_, _34698_, _09403_);
  nor (_16084_, _08262_, \oc8051_golden_model_1.DPH [0]);
  nor (_16085_, _16084_, _08349_);
  and (_16086_, _16085_, _08250_);
  nor (_16087_, _05038_, _09403_);
  and (_16088_, _05044_, _04632_);
  or (_16090_, _16088_, _16087_);
  or (_16091_, _16090_, _03821_);
  and (_16092_, _05038_, \oc8051_golden_model_1.ACC [0]);
  or (_16093_, _16092_, _16087_);
  and (_16094_, _16093_, _03825_);
  nor (_16095_, _03825_, _09403_);
  or (_16096_, _16095_, _02952_);
  or (_16097_, _16096_, _16094_);
  and (_16098_, _16097_, _03327_);
  and (_16099_, _16098_, _16091_);
  and (_16101_, _04632_, _03817_);
  or (_16102_, _16101_, _16087_);
  and (_16103_, _16102_, _02947_);
  or (_16104_, _16103_, _02950_);
  or (_16105_, _16104_, _16099_);
  or (_16106_, _16093_, _02959_);
  and (_16107_, _16106_, _08251_);
  and (_16108_, _16107_, _16105_);
  or (_16109_, _16108_, _16086_);
  and (_16110_, _16109_, _08235_);
  nor (_16112_, _02832_, _08235_);
  or (_16113_, _16112_, _06793_);
  or (_16114_, _16113_, _16110_);
  or (_16115_, _16102_, _06241_);
  and (_16116_, _16115_, _16114_);
  or (_16117_, _16116_, _02855_);
  and (_16118_, _06174_, _05038_);
  or (_16119_, _16087_, _02856_);
  or (_16120_, _16119_, _16118_);
  and (_16121_, _16120_, _16117_);
  or (_16123_, _16121_, _02576_);
  nor (_16124_, _10530_, _08328_);
  or (_16125_, _16087_, _02851_);
  or (_16126_, _16125_, _16124_);
  and (_16127_, _16126_, _03884_);
  and (_16128_, _16127_, _16123_);
  and (_16129_, _05038_, _05566_);
  or (_16130_, _16129_, _16087_);
  and (_16131_, _16130_, _03014_);
  or (_16132_, _16131_, _03021_);
  or (_16134_, _16132_, _16128_);
  and (_16135_, _10425_, _05038_);
  or (_16136_, _16135_, _16087_);
  or (_16137_, _16136_, _05279_);
  and (_16138_, _16137_, _16134_);
  or (_16139_, _16138_, _03130_);
  and (_16140_, _10546_, _04632_);
  or (_16141_, _16087_, _03131_);
  or (_16142_, _16141_, _16140_);
  and (_16143_, _16142_, _05274_);
  and (_16145_, _16143_, _16139_);
  nand (_16146_, _16130_, _03020_);
  nor (_16147_, _16146_, _16088_);
  or (_16148_, _16147_, _16145_);
  and (_16149_, _16148_, _03140_);
  or (_16150_, _16087_, _09183_);
  and (_16151_, _16093_, _03139_);
  and (_16152_, _16151_, _16150_);
  or (_16153_, _16152_, _03036_);
  or (_16154_, _16153_, _16149_);
  nor (_16156_, _10423_, _08372_);
  or (_16157_, _16156_, _16087_);
  or (_16158_, _16157_, _05781_);
  and (_16159_, _16158_, _05786_);
  and (_16160_, _16159_, _16154_);
  nor (_16161_, _10421_, _08328_);
  or (_16162_, _16161_, _16087_);
  and (_16163_, _16162_, _03127_);
  or (_16164_, _16163_, _15506_);
  or (_16165_, _16164_, _16160_);
  or (_16167_, _16090_, _03265_);
  and (_16168_, _16167_, _34698_);
  and (_16169_, _16168_, _16165_);
  or (_16170_, _16169_, _16083_);
  and (_35180_, _16170_, _36029_);
  not (_16171_, \oc8051_golden_model_1.DPH [1]);
  nor (_16172_, _34698_, _16171_);
  or (_16173_, _10739_, _08328_);
  or (_16174_, _05038_, \oc8051_golden_model_1.DPH [1]);
  and (_16175_, _16174_, _03130_);
  and (_16177_, _16175_, _16173_);
  and (_16178_, _16174_, _03014_);
  nand (_16179_, _04632_, _03705_);
  and (_16180_, _16179_, _16178_);
  nor (_16181_, _08349_, \oc8051_golden_model_1.DPH [1]);
  nor (_16182_, _16181_, _08350_);
  and (_16183_, _16182_, _08250_);
  nand (_16184_, _10622_, _04632_);
  and (_16185_, _16184_, _16174_);
  or (_16186_, _16185_, _03821_);
  nand (_16188_, _04632_, _02618_);
  and (_16189_, _16188_, _16174_);
  and (_16190_, _16189_, _03825_);
  nor (_16191_, _03825_, _16171_);
  or (_16192_, _16191_, _02952_);
  or (_16193_, _16192_, _16190_);
  and (_16194_, _16193_, _03327_);
  and (_16195_, _16194_, _16186_);
  nor (_16196_, _05038_, _16171_);
  and (_16197_, _04632_, _04005_);
  or (_16199_, _16197_, _16196_);
  and (_16200_, _16199_, _02947_);
  or (_16201_, _16200_, _02950_);
  or (_16202_, _16201_, _16195_);
  or (_16203_, _16189_, _02959_);
  and (_16204_, _16203_, _08251_);
  and (_16205_, _16204_, _16202_);
  or (_16206_, _16205_, _16183_);
  and (_16207_, _16206_, _08235_);
  nor (_16208_, _03671_, _08235_);
  or (_16210_, _16208_, _06793_);
  or (_16211_, _16210_, _16207_);
  or (_16212_, _16199_, _06241_);
  and (_16213_, _16212_, _16211_);
  or (_16214_, _16213_, _02855_);
  and (_16215_, _06173_, _05038_);
  or (_16216_, _16196_, _02856_);
  or (_16217_, _16216_, _16215_);
  and (_16218_, _16217_, _02851_);
  and (_16219_, _16218_, _16214_);
  and (_16221_, _16174_, _02576_);
  nand (_16222_, _10720_, _04632_);
  and (_16223_, _16222_, _16221_);
  or (_16224_, _16223_, _16219_);
  and (_16225_, _16224_, _03884_);
  or (_16226_, _16225_, _16180_);
  and (_16227_, _16226_, _05279_);
  or (_16228_, _10612_, _08328_);
  and (_16229_, _16174_, _03021_);
  and (_16230_, _16229_, _16228_);
  or (_16232_, _16230_, _16227_);
  and (_16233_, _16232_, _03131_);
  or (_16234_, _16233_, _16177_);
  and (_16235_, _16234_, _05274_);
  or (_16236_, _10611_, _08328_);
  and (_16237_, _16174_, _03020_);
  and (_16238_, _16237_, _16236_);
  or (_16239_, _16238_, _16235_);
  and (_16240_, _16239_, _03140_);
  or (_16241_, _16196_, _12724_);
  and (_16243_, _16189_, _03139_);
  and (_16244_, _16243_, _16241_);
  or (_16245_, _16244_, _16240_);
  and (_16246_, _16245_, _03128_);
  or (_16247_, _16188_, _12724_);
  and (_16248_, _16174_, _03127_);
  and (_16249_, _16248_, _16247_);
  or (_16250_, _16249_, _03166_);
  or (_16251_, _16179_, _12724_);
  and (_16252_, _16174_, _03036_);
  and (_16254_, _16252_, _16251_);
  or (_16255_, _16254_, _16250_);
  or (_16256_, _16255_, _16246_);
  or (_16257_, _16185_, _03563_);
  and (_16258_, _16257_, _16256_);
  or (_16259_, _16258_, _03174_);
  nor (_16260_, _16196_, _03178_);
  nand (_16261_, _16260_, _16184_);
  and (_16262_, _16261_, _34698_);
  and (_16263_, _16262_, _16259_);
  or (_16265_, _16263_, _16172_);
  and (_35182_, _16265_, _36029_);
  not (_16266_, \oc8051_golden_model_1.DPH [2]);
  nor (_16267_, _34698_, _16266_);
  nor (_16268_, _05038_, _16266_);
  nor (_16269_, _10830_, _08328_);
  or (_16270_, _16269_, _16268_);
  and (_16271_, _16270_, _03127_);
  and (_16272_, _10831_, _04632_);
  or (_16273_, _16272_, _16268_);
  and (_16275_, _16273_, _03130_);
  nor (_16276_, _08328_, _04440_);
  or (_16277_, _16276_, _16268_);
  or (_16278_, _16277_, _06241_);
  or (_16279_, _08350_, \oc8051_golden_model_1.DPH [2]);
  nor (_16280_, _08351_, _08251_);
  and (_16281_, _16280_, _16279_);
  nor (_16282_, _10849_, _08328_);
  or (_16283_, _16282_, _16268_);
  or (_16284_, _16283_, _03821_);
  and (_16286_, _05038_, \oc8051_golden_model_1.ACC [2]);
  or (_16287_, _16286_, _16268_);
  and (_16288_, _16287_, _03825_);
  nor (_16289_, _03825_, _16266_);
  or (_16290_, _16289_, _02952_);
  or (_16291_, _16290_, _16288_);
  and (_16292_, _16291_, _03327_);
  and (_16293_, _16292_, _16284_);
  and (_16294_, _16277_, _02947_);
  or (_16295_, _16294_, _02950_);
  or (_16297_, _16295_, _16293_);
  or (_16298_, _16287_, _02959_);
  and (_16299_, _16298_, _08251_);
  and (_16300_, _16299_, _16297_);
  or (_16301_, _16300_, _16281_);
  and (_16302_, _16301_, _08235_);
  nor (_16303_, _03260_, _08235_);
  or (_16304_, _16303_, _06793_);
  or (_16305_, _16304_, _16302_);
  and (_16306_, _16305_, _16278_);
  or (_16308_, _16306_, _02855_);
  or (_16309_, _16268_, _02856_);
  and (_16310_, _06177_, _05038_);
  or (_16311_, _16310_, _16309_);
  and (_16312_, _16311_, _02851_);
  and (_16313_, _16312_, _16308_);
  nor (_16314_, _10943_, _08372_);
  or (_16315_, _16314_, _16268_);
  and (_16316_, _16315_, _02576_);
  or (_16317_, _16316_, _03014_);
  or (_16319_, _16317_, _16313_);
  and (_16320_, _05038_, _05727_);
  or (_16321_, _16320_, _16268_);
  or (_16322_, _16321_, _03884_);
  and (_16323_, _16322_, _16319_);
  or (_16324_, _16323_, _03021_);
  and (_16325_, _10835_, _04632_);
  or (_16326_, _16268_, _05279_);
  or (_16327_, _16326_, _16325_);
  and (_16328_, _16327_, _03131_);
  and (_16330_, _16328_, _16324_);
  or (_16331_, _16330_, _16275_);
  and (_16332_, _16331_, _05274_);
  or (_16333_, _16268_, _05143_);
  and (_16334_, _16321_, _03020_);
  and (_16335_, _16334_, _16333_);
  or (_16336_, _16335_, _16332_);
  and (_16337_, _16336_, _03140_);
  and (_16338_, _16287_, _03139_);
  and (_16339_, _16338_, _16333_);
  or (_16341_, _16339_, _03036_);
  or (_16342_, _16341_, _16337_);
  nor (_16343_, _10833_, _08328_);
  or (_16344_, _16268_, _05781_);
  or (_16345_, _16344_, _16343_);
  and (_16346_, _16345_, _05786_);
  and (_16347_, _16346_, _16342_);
  or (_16348_, _16347_, _16271_);
  and (_16349_, _16348_, _03563_);
  and (_16350_, _16283_, _03166_);
  or (_16352_, _16350_, _03174_);
  or (_16353_, _16352_, _16349_);
  and (_16354_, _11008_, _04632_);
  or (_16355_, _16268_, _03178_);
  or (_16356_, _16355_, _16354_);
  and (_16357_, _16356_, _34698_);
  and (_16358_, _16357_, _16353_);
  or (_16359_, _16358_, _16267_);
  and (_35183_, _16359_, _36029_);
  or (_16360_, _34698_, \oc8051_golden_model_1.DPH [3]);
  and (_16362_, _16360_, _36029_);
  not (_16363_, \oc8051_golden_model_1.DPH [3]);
  nor (_16364_, _05038_, _16363_);
  and (_16365_, _11028_, _04632_);
  or (_16366_, _16365_, _16364_);
  and (_16367_, _16366_, _03130_);
  nor (_16368_, _08328_, _04242_);
  or (_16369_, _16368_, _16364_);
  or (_16370_, _16369_, _06241_);
  or (_16371_, _08351_, \oc8051_golden_model_1.DPH [3]);
  nor (_16373_, _08352_, _08251_);
  and (_16374_, _16373_, _16371_);
  nor (_16375_, _11040_, _08328_);
  or (_16376_, _16375_, _16364_);
  or (_16377_, _16376_, _03821_);
  and (_16378_, _05038_, \oc8051_golden_model_1.ACC [3]);
  or (_16379_, _16378_, _16364_);
  and (_16380_, _16379_, _03825_);
  nor (_16381_, _03825_, _16363_);
  or (_16382_, _16381_, _02952_);
  or (_16384_, _16382_, _16380_);
  and (_16385_, _16384_, _03327_);
  and (_16386_, _16385_, _16377_);
  and (_16387_, _16369_, _02947_);
  or (_16388_, _16387_, _02950_);
  or (_16389_, _16388_, _16386_);
  or (_16390_, _16379_, _02959_);
  and (_16391_, _16390_, _08251_);
  and (_16392_, _16391_, _16389_);
  or (_16393_, _16392_, _16374_);
  and (_16395_, _16393_, _08235_);
  nor (_16396_, _08235_, _02799_);
  or (_16397_, _16396_, _06793_);
  or (_16398_, _16397_, _16395_);
  and (_16399_, _16398_, _16370_);
  or (_16400_, _16399_, _02855_);
  or (_16401_, _16364_, _02856_);
  and (_16402_, _06176_, _05038_);
  or (_16403_, _16402_, _16401_);
  and (_16404_, _16403_, _02851_);
  and (_16406_, _16404_, _16400_);
  nor (_16407_, _11143_, _08372_);
  or (_16408_, _16407_, _16364_);
  and (_16409_, _16408_, _02576_);
  or (_16410_, _16409_, _03014_);
  or (_16411_, _16410_, _16406_);
  and (_16412_, _05038_, _05664_);
  or (_16413_, _16412_, _16364_);
  or (_16414_, _16413_, _03884_);
  and (_16415_, _16414_, _16411_);
  or (_16417_, _16415_, _03021_);
  and (_16418_, _11032_, _04632_);
  or (_16419_, _16364_, _05279_);
  or (_16420_, _16419_, _16418_);
  and (_16421_, _16420_, _03131_);
  and (_16422_, _16421_, _16417_);
  or (_16423_, _16422_, _16367_);
  and (_16424_, _16423_, _05274_);
  or (_16425_, _16364_, _04996_);
  and (_16426_, _16413_, _03020_);
  and (_16428_, _16426_, _16425_);
  or (_16429_, _16428_, _16424_);
  and (_16430_, _16429_, _03140_);
  and (_16431_, _16379_, _03139_);
  and (_16432_, _16431_, _16425_);
  or (_16433_, _16432_, _03036_);
  or (_16434_, _16433_, _16430_);
  nor (_16435_, _11030_, _08328_);
  or (_16436_, _16364_, _05781_);
  or (_16437_, _16436_, _16435_);
  and (_16439_, _16437_, _05786_);
  and (_16440_, _16439_, _16434_);
  nor (_16441_, _11027_, _08328_);
  or (_16442_, _16441_, _16364_);
  and (_16443_, _16442_, _03127_);
  or (_16444_, _16443_, _03166_);
  or (_16445_, _16444_, _16440_);
  or (_16446_, _16376_, _03563_);
  and (_16447_, _16446_, _03178_);
  and (_16448_, _16447_, _16445_);
  and (_16450_, _11213_, _04632_);
  or (_16451_, _16450_, _16364_);
  and (_16452_, _16451_, _03174_);
  or (_16453_, _16452_, _34702_);
  or (_16454_, _16453_, _16448_);
  and (_35184_, _16454_, _16362_);
  or (_16455_, _34698_, \oc8051_golden_model_1.DPH [4]);
  and (_16456_, _16455_, _36029_);
  not (_16457_, \oc8051_golden_model_1.DPH [4]);
  nor (_16458_, _05038_, _16457_);
  and (_16460_, _11368_, _04632_);
  or (_16461_, _16460_, _16458_);
  and (_16462_, _16461_, _03130_);
  nor (_16463_, _05202_, _08328_);
  or (_16464_, _16463_, _16458_);
  or (_16465_, _16464_, _06241_);
  nor (_16466_, _11259_, _08328_);
  or (_16467_, _16466_, _16458_);
  or (_16468_, _16467_, _03821_);
  and (_16469_, _05038_, \oc8051_golden_model_1.ACC [4]);
  or (_16471_, _16469_, _16458_);
  and (_16472_, _16471_, _03825_);
  nor (_16473_, _03825_, _16457_);
  or (_16474_, _16473_, _02952_);
  or (_16475_, _16474_, _16472_);
  and (_16476_, _16475_, _03327_);
  and (_16477_, _16476_, _16468_);
  and (_16478_, _16464_, _02947_);
  or (_16479_, _16478_, _02950_);
  or (_16480_, _16479_, _16477_);
  or (_16482_, _16471_, _02959_);
  and (_16483_, _16482_, _08251_);
  and (_16484_, _16483_, _16480_);
  or (_16485_, _08352_, \oc8051_golden_model_1.DPH [4]);
  nor (_16486_, _08353_, _08251_);
  and (_16487_, _16486_, _16485_);
  or (_16488_, _16487_, _16484_);
  and (_16489_, _16488_, _08235_);
  nor (_16490_, _03625_, _08235_);
  or (_16491_, _16490_, _06793_);
  or (_16493_, _16491_, _16489_);
  and (_16494_, _16493_, _16465_);
  or (_16495_, _16494_, _02855_);
  or (_16496_, _16458_, _02856_);
  and (_16497_, _06181_, _05038_);
  or (_16498_, _16497_, _16496_);
  and (_16499_, _16498_, _02851_);
  and (_16500_, _16499_, _16495_);
  nor (_16501_, _11348_, _08372_);
  or (_16502_, _16501_, _16458_);
  and (_16504_, _16502_, _02576_);
  or (_16505_, _16504_, _03014_);
  or (_16506_, _16505_, _16500_);
  and (_16507_, _05697_, _05038_);
  or (_16508_, _16507_, _16458_);
  or (_16509_, _16508_, _03884_);
  and (_16510_, _16509_, _16506_);
  or (_16511_, _16510_, _03021_);
  and (_16512_, _11362_, _04632_);
  or (_16513_, _16458_, _05279_);
  or (_16515_, _16513_, _16512_);
  and (_16516_, _16515_, _03131_);
  and (_16517_, _16516_, _16511_);
  or (_16518_, _16517_, _16462_);
  and (_16519_, _16518_, _05274_);
  or (_16520_, _16458_, _05251_);
  and (_16521_, _16508_, _03020_);
  and (_16522_, _16521_, _16520_);
  or (_16523_, _16522_, _16519_);
  and (_16524_, _16523_, _03140_);
  and (_16526_, _16471_, _03139_);
  and (_16527_, _16526_, _16520_);
  or (_16528_, _16527_, _03036_);
  or (_16529_, _16528_, _16524_);
  nor (_16530_, _11361_, _08328_);
  or (_16531_, _16458_, _05781_);
  or (_16532_, _16531_, _16530_);
  and (_16533_, _16532_, _05786_);
  and (_16534_, _16533_, _16529_);
  nor (_16535_, _11367_, _08328_);
  or (_16537_, _16535_, _16458_);
  and (_16538_, _16537_, _03127_);
  or (_16539_, _16538_, _03166_);
  or (_16540_, _16539_, _16534_);
  or (_16541_, _16467_, _03563_);
  and (_16542_, _16541_, _03178_);
  and (_16543_, _16542_, _16540_);
  and (_16544_, _11417_, _04632_);
  or (_16545_, _16544_, _16458_);
  and (_16546_, _16545_, _03174_);
  or (_16548_, _16546_, _34702_);
  or (_16549_, _16548_, _16543_);
  and (_35185_, _16549_, _16456_);
  or (_16550_, _34698_, \oc8051_golden_model_1.DPH [5]);
  and (_16551_, _16550_, _36029_);
  not (_16552_, \oc8051_golden_model_1.DPH [5]);
  nor (_16553_, _05038_, _16552_);
  and (_16554_, _11436_, _04632_);
  or (_16555_, _16554_, _16553_);
  and (_16556_, _16555_, _03130_);
  nor (_16558_, _04896_, _08328_);
  or (_16559_, _16558_, _16553_);
  or (_16560_, _16559_, _06241_);
  nor (_16561_, _11445_, _08328_);
  or (_16562_, _16561_, _16553_);
  or (_16563_, _16562_, _03821_);
  and (_16564_, _05038_, \oc8051_golden_model_1.ACC [5]);
  or (_16565_, _16564_, _16553_);
  and (_16566_, _16565_, _03825_);
  nor (_16567_, _03825_, _16552_);
  or (_16569_, _16567_, _02952_);
  or (_16570_, _16569_, _16566_);
  and (_16571_, _16570_, _03327_);
  and (_16572_, _16571_, _16563_);
  and (_16573_, _16559_, _02947_);
  or (_16574_, _16573_, _02950_);
  or (_16575_, _16574_, _16572_);
  or (_16576_, _16565_, _02959_);
  and (_16577_, _16576_, _08251_);
  and (_16578_, _16577_, _16575_);
  or (_16580_, _08353_, \oc8051_golden_model_1.DPH [5]);
  nor (_16581_, _08354_, _08251_);
  and (_16582_, _16581_, _16580_);
  or (_16583_, _16582_, _16578_);
  and (_16584_, _16583_, _08235_);
  nor (_16585_, _03215_, _08235_);
  or (_16586_, _16585_, _06793_);
  or (_16587_, _16586_, _16584_);
  and (_16588_, _16587_, _16560_);
  or (_16589_, _16588_, _02855_);
  or (_16591_, _16553_, _02856_);
  and (_16592_, _06180_, _05038_);
  or (_16593_, _16592_, _16591_);
  and (_16594_, _16593_, _02851_);
  and (_16595_, _16594_, _16589_);
  nor (_16596_, _11546_, _08372_);
  or (_16597_, _16596_, _16553_);
  and (_16598_, _16597_, _02576_);
  or (_16599_, _16598_, _03014_);
  or (_16600_, _16599_, _16595_);
  and (_16602_, _05701_, _05038_);
  or (_16603_, _16602_, _16553_);
  or (_16604_, _16603_, _03884_);
  and (_16605_, _16604_, _16600_);
  or (_16606_, _16605_, _03021_);
  and (_16607_, _11562_, _04632_);
  or (_16608_, _16553_, _05279_);
  or (_16609_, _16608_, _16607_);
  and (_16610_, _16609_, _03131_);
  and (_16611_, _16610_, _16606_);
  or (_16613_, _16611_, _16556_);
  and (_16614_, _16613_, _05274_);
  or (_16615_, _16553_, _04944_);
  and (_16616_, _16603_, _03020_);
  and (_16617_, _16616_, _16615_);
  or (_16618_, _16617_, _16614_);
  and (_16619_, _16618_, _03140_);
  and (_16620_, _16565_, _03139_);
  and (_16621_, _16620_, _16615_);
  or (_16622_, _16621_, _03036_);
  or (_16624_, _16622_, _16619_);
  nor (_16625_, _11560_, _08328_);
  or (_16626_, _16553_, _05781_);
  or (_16627_, _16626_, _16625_);
  and (_16628_, _16627_, _05786_);
  and (_16629_, _16628_, _16624_);
  nor (_16630_, _11435_, _08328_);
  or (_16631_, _16630_, _16553_);
  and (_16632_, _16631_, _03127_);
  or (_16633_, _16632_, _03166_);
  or (_16635_, _16633_, _16629_);
  or (_16636_, _16562_, _03563_);
  and (_16637_, _16636_, _03178_);
  and (_16638_, _16637_, _16635_);
  and (_16639_, _11619_, _04632_);
  or (_16640_, _16639_, _16553_);
  and (_16641_, _16640_, _03174_);
  or (_16642_, _16641_, _34702_);
  or (_16643_, _16642_, _16638_);
  and (_35186_, _16643_, _16551_);
  or (_16645_, _34698_, \oc8051_golden_model_1.DPH [6]);
  and (_16646_, _16645_, _36029_);
  not (_16647_, \oc8051_golden_model_1.DPH [6]);
  nor (_16648_, _05038_, _16647_);
  and (_16649_, _11769_, _04632_);
  or (_16650_, _16649_, _16648_);
  and (_16651_, _16650_, _03130_);
  nor (_16652_, _04787_, _08328_);
  or (_16653_, _16652_, _16648_);
  or (_16654_, _16653_, _06241_);
  nor (_16656_, _11636_, _08328_);
  or (_16657_, _16656_, _16648_);
  or (_16658_, _16657_, _03821_);
  and (_16659_, _05038_, \oc8051_golden_model_1.ACC [6]);
  or (_16660_, _16659_, _16648_);
  and (_16661_, _16660_, _03825_);
  nor (_16662_, _03825_, _16647_);
  or (_16663_, _16662_, _02952_);
  or (_16664_, _16663_, _16661_);
  and (_16665_, _16664_, _03327_);
  and (_16667_, _16665_, _16658_);
  and (_16668_, _16653_, _02947_);
  or (_16669_, _16668_, _02950_);
  or (_16670_, _16669_, _16667_);
  or (_16671_, _16660_, _02959_);
  and (_16672_, _16671_, _08251_);
  and (_16673_, _16672_, _16670_);
  or (_16674_, _08354_, \oc8051_golden_model_1.DPH [6]);
  nor (_16675_, _08355_, _08251_);
  and (_16676_, _16675_, _16674_);
  or (_16678_, _16676_, _16673_);
  and (_16679_, _16678_, _08235_);
  nor (_16680_, _08235_, _02932_);
  or (_16681_, _16680_, _06793_);
  or (_16682_, _16681_, _16679_);
  and (_16683_, _16682_, _16654_);
  or (_16684_, _16683_, _02855_);
  or (_16685_, _16648_, _02856_);
  and (_16686_, _05847_, _05038_);
  or (_16687_, _16686_, _16685_);
  and (_16690_, _16687_, _02851_);
  and (_16691_, _16690_, _16684_);
  nor (_16692_, _11751_, _08372_);
  or (_16693_, _16692_, _16648_);
  and (_16694_, _16693_, _02576_);
  or (_16695_, _16694_, _03014_);
  or (_16696_, _16695_, _16691_);
  and (_16697_, _11758_, _05038_);
  or (_16698_, _16697_, _16648_);
  or (_16699_, _16698_, _03884_);
  and (_16701_, _16699_, _16696_);
  or (_16702_, _16701_, _03021_);
  and (_16703_, _11646_, _04632_);
  or (_16704_, _16648_, _05279_);
  or (_16705_, _16704_, _16703_);
  and (_16706_, _16705_, _03131_);
  and (_16707_, _16706_, _16702_);
  or (_16708_, _16707_, _16651_);
  and (_16709_, _16708_, _05274_);
  or (_16710_, _16648_, _04838_);
  and (_16712_, _16698_, _03020_);
  and (_16713_, _16712_, _16710_);
  or (_16714_, _16713_, _16709_);
  and (_16715_, _16714_, _03140_);
  and (_16716_, _16660_, _03139_);
  and (_16717_, _16716_, _16710_);
  or (_16718_, _16717_, _03036_);
  or (_16719_, _16718_, _16715_);
  nor (_16720_, _11644_, _08328_);
  or (_16721_, _16648_, _05781_);
  or (_16723_, _16721_, _16720_);
  and (_16724_, _16723_, _05786_);
  and (_16725_, _16724_, _16719_);
  nor (_16726_, _11768_, _08328_);
  or (_16727_, _16726_, _16648_);
  and (_16728_, _16727_, _03127_);
  or (_16729_, _16728_, _03166_);
  or (_16730_, _16729_, _16725_);
  or (_16731_, _16657_, _03563_);
  and (_16732_, _16731_, _03178_);
  and (_16734_, _16732_, _16730_);
  and (_16735_, _11821_, _04632_);
  or (_16736_, _16735_, _16648_);
  and (_16737_, _16736_, _03174_);
  or (_16738_, _16737_, _34702_);
  or (_16739_, _16738_, _16734_);
  and (_35187_, _16739_, _16646_);
  and (_35188_, \oc8051_golden_model_1.IE [0], _36029_);
  and (_35189_, \oc8051_golden_model_1.IE [1], _36029_);
  and (_35190_, \oc8051_golden_model_1.IE [2], _36029_);
  and (_35191_, \oc8051_golden_model_1.IE [3], _36029_);
  and (_35193_, \oc8051_golden_model_1.IE [4], _36029_);
  and (_35194_, \oc8051_golden_model_1.IE [5], _36029_);
  and (_35195_, \oc8051_golden_model_1.IE [6], _36029_);
  and (_35196_, \oc8051_golden_model_1.IP [0], _36029_);
  and (_35197_, \oc8051_golden_model_1.IP [1], _36029_);
  and (_35198_, \oc8051_golden_model_1.IP [2], _36029_);
  and (_35199_, \oc8051_golden_model_1.IP [3], _36029_);
  and (_35200_, \oc8051_golden_model_1.IP [4], _36029_);
  and (_35201_, \oc8051_golden_model_1.IP [5], _36029_);
  and (_35202_, \oc8051_golden_model_1.IP [6], _36029_);
  not (_16742_, \oc8051_golden_model_1.P0 [0]);
  nor (_16743_, _34698_, _16742_);
  or (_16744_, _16743_, rst);
  and (_16745_, _05044_, _04716_);
  nor (_16746_, _04716_, _16742_);
  and (_16747_, _04716_, _05566_);
  or (_16748_, _16747_, _16746_);
  nand (_16749_, _16748_, _03020_);
  nor (_16750_, _16749_, _16745_);
  and (_16752_, _10546_, _04716_);
  or (_16753_, _16752_, _16746_);
  and (_16754_, _16753_, _03130_);
  and (_16755_, _04716_, _03817_);
  or (_16756_, _16755_, _16746_);
  or (_16757_, _16756_, _06241_);
  or (_16758_, _16746_, _16745_);
  and (_16759_, _16758_, _02952_);
  nor (_16760_, _03825_, _16742_);
  and (_16761_, _04716_, \oc8051_golden_model_1.ACC [0]);
  or (_16763_, _16761_, _16746_);
  and (_16764_, _16763_, _03825_);
  or (_16765_, _16764_, _16760_);
  and (_16766_, _16765_, _03821_);
  or (_16767_, _16766_, _02891_);
  or (_16768_, _16767_, _16759_);
  and (_16769_, _10429_, _04629_);
  nor (_16770_, _04629_, _16742_);
  or (_16771_, _16770_, _02892_);
  or (_16772_, _16771_, _16769_);
  and (_16774_, _16772_, _03327_);
  and (_16775_, _16774_, _16768_);
  and (_16776_, _16756_, _02947_);
  or (_16777_, _16776_, _02950_);
  or (_16778_, _16777_, _16775_);
  or (_16779_, _16763_, _02959_);
  and (_16780_, _16779_, _02888_);
  and (_16781_, _16780_, _16778_);
  and (_16782_, _16746_, _02887_);
  or (_16783_, _16782_, _02880_);
  or (_16785_, _16783_, _16781_);
  or (_16786_, _16758_, _02881_);
  and (_16787_, _16786_, _02875_);
  and (_16788_, _16787_, _16785_);
  or (_16789_, _10472_, _10452_);
  and (_16790_, _16789_, _04629_);
  or (_16791_, _16790_, _16770_);
  and (_16792_, _16791_, _02874_);
  or (_16793_, _16792_, _06793_);
  or (_16794_, _16793_, _16788_);
  and (_16796_, _16794_, _16757_);
  or (_16797_, _16796_, _02855_);
  and (_16798_, _06174_, _04716_);
  or (_16799_, _16746_, _02856_);
  or (_16800_, _16799_, _16798_);
  and (_16801_, _16800_, _02851_);
  and (_16802_, _16801_, _16797_);
  and (_16803_, _05733_, \oc8051_golden_model_1.P1 [0]);
  and (_16804_, _05736_, \oc8051_golden_model_1.P0 [0]);
  and (_16805_, _05739_, \oc8051_golden_model_1.P2 [0]);
  and (_16807_, _05741_, \oc8051_golden_model_1.P3 [0]);
  or (_16808_, _16807_, _16805_);
  or (_16809_, _16808_, _16804_);
  nor (_16810_, _16809_, _16803_);
  and (_16811_, _16810_, _10525_);
  and (_16812_, _16811_, _10513_);
  nand (_16813_, _16812_, _10506_);
  or (_16814_, _16813_, _10485_);
  and (_16815_, _16814_, _04716_);
  or (_16816_, _16815_, _16746_);
  and (_16818_, _16816_, _02576_);
  or (_16819_, _16818_, _03014_);
  or (_16820_, _16819_, _16802_);
  or (_16821_, _16748_, _03884_);
  and (_16822_, _16821_, _16820_);
  or (_16823_, _16822_, _03021_);
  and (_16824_, _10425_, _04716_);
  or (_16825_, _16746_, _05279_);
  or (_16826_, _16825_, _16824_);
  and (_16827_, _16826_, _03131_);
  and (_16829_, _16827_, _16823_);
  or (_16830_, _16829_, _16754_);
  and (_16831_, _16830_, _05274_);
  or (_16832_, _16831_, _16750_);
  and (_16833_, _16832_, _03140_);
  or (_16834_, _16746_, _09183_);
  and (_16835_, _16763_, _03139_);
  and (_16836_, _16835_, _16834_);
  or (_16837_, _16836_, _03036_);
  or (_16838_, _16837_, _16833_);
  nor (_16840_, _10423_, _08424_);
  or (_16841_, _16746_, _05781_);
  or (_16842_, _16841_, _16840_);
  and (_16843_, _16842_, _05786_);
  and (_16844_, _16843_, _16838_);
  nor (_16845_, _10421_, _08424_);
  or (_16846_, _16845_, _16746_);
  and (_16847_, _16846_, _03127_);
  or (_16848_, _16847_, _03166_);
  or (_16849_, _16848_, _16844_);
  or (_16851_, _16758_, _03563_);
  and (_16852_, _16851_, _02501_);
  and (_16853_, _16852_, _16849_);
  and (_16854_, _16746_, _02500_);
  or (_16855_, _16854_, _03174_);
  or (_16856_, _16855_, _16853_);
  or (_16857_, _16758_, _03178_);
  and (_16858_, _16857_, _34698_);
  and (_16859_, _16858_, _16856_);
  or (_35204_, _16859_, _16744_);
  not (_16861_, \oc8051_golden_model_1.P0 [1]);
  nor (_16862_, _34698_, _16861_);
  or (_16863_, _16862_, rst);
  nand (_16864_, _04716_, _03705_);
  or (_16865_, _04716_, \oc8051_golden_model_1.P0 [1]);
  and (_16866_, _16865_, _03014_);
  and (_16867_, _16866_, _16864_);
  and (_16868_, _10622_, _04716_);
  not (_16869_, _16868_);
  and (_16870_, _16869_, _16865_);
  or (_16872_, _16870_, _03821_);
  nand (_16873_, _04716_, _02618_);
  and (_16874_, _16873_, _16865_);
  and (_16875_, _16874_, _03825_);
  nor (_16876_, _03825_, _16861_);
  or (_16877_, _16876_, _02952_);
  or (_16878_, _16877_, _16875_);
  and (_16879_, _16878_, _02892_);
  and (_16880_, _16879_, _16872_);
  and (_16881_, _10617_, _04629_);
  nor (_16883_, _04629_, _16861_);
  or (_16884_, _16883_, _02947_);
  or (_16885_, _16884_, _16881_);
  and (_16886_, _16885_, _09918_);
  or (_16887_, _16886_, _16880_);
  nor (_16888_, _04716_, _16861_);
  and (_16889_, _04716_, _04005_);
  or (_16890_, _16889_, _16888_);
  or (_16891_, _16890_, _03327_);
  and (_16892_, _16891_, _16887_);
  or (_16894_, _16892_, _02950_);
  or (_16895_, _16874_, _02959_);
  and (_16896_, _16895_, _02888_);
  and (_16897_, _16896_, _16894_);
  and (_16898_, _10620_, _04629_);
  or (_16899_, _16898_, _16883_);
  and (_16900_, _16899_, _02887_);
  or (_16901_, _16900_, _02880_);
  or (_16902_, _16901_, _16897_);
  and (_16903_, _16881_, _10616_);
  or (_16905_, _16883_, _02881_);
  or (_16906_, _16905_, _16903_);
  and (_16907_, _16906_, _16902_);
  and (_16908_, _16907_, _02875_);
  or (_16909_, _10660_, _10620_);
  and (_16910_, _16909_, _04629_);
  or (_16911_, _16883_, _16910_);
  and (_16912_, _16911_, _02874_);
  or (_16913_, _16912_, _06793_);
  or (_16914_, _16913_, _16908_);
  or (_16916_, _16890_, _06241_);
  and (_16917_, _16916_, _16914_);
  or (_16918_, _16917_, _02855_);
  and (_16919_, _06173_, _04716_);
  or (_16920_, _16888_, _02856_);
  or (_16921_, _16920_, _16919_);
  and (_16922_, _16921_, _02851_);
  and (_16923_, _16922_, _16918_);
  and (_16924_, _05733_, \oc8051_golden_model_1.P1 [1]);
  and (_16925_, _05736_, \oc8051_golden_model_1.P0 [1]);
  and (_16927_, _05739_, \oc8051_golden_model_1.P2 [1]);
  and (_16928_, _05741_, \oc8051_golden_model_1.P3 [1]);
  or (_16929_, _16928_, _16927_);
  or (_16930_, _16929_, _16925_);
  nor (_16931_, _16930_, _16924_);
  and (_16932_, _16931_, _10685_);
  and (_16933_, _16932_, _10680_);
  nand (_16934_, _16933_, _10717_);
  or (_16935_, _16934_, _10673_);
  and (_16936_, _16935_, _04716_);
  or (_16938_, _16936_, _16888_);
  and (_16939_, _16938_, _02576_);
  or (_16940_, _16939_, _16923_);
  and (_16941_, _16940_, _03884_);
  or (_16942_, _16941_, _16867_);
  and (_16943_, _16942_, _05279_);
  or (_16944_, _10612_, _08424_);
  and (_16945_, _16865_, _03021_);
  and (_16946_, _16945_, _16944_);
  or (_16947_, _16946_, _16943_);
  and (_16949_, _16947_, _03131_);
  or (_16950_, _10739_, _08424_);
  and (_16951_, _16865_, _03130_);
  and (_16952_, _16951_, _16950_);
  or (_16953_, _16952_, _16949_);
  and (_16954_, _16953_, _05274_);
  or (_16955_, _10611_, _08424_);
  and (_16956_, _16865_, _03020_);
  and (_16957_, _16956_, _16955_);
  or (_16958_, _16957_, _16954_);
  and (_16960_, _16958_, _03140_);
  or (_16961_, _16888_, _12724_);
  and (_16962_, _16874_, _03139_);
  and (_16963_, _16962_, _16961_);
  or (_16964_, _16963_, _16960_);
  and (_16965_, _16964_, _03128_);
  or (_16966_, _16864_, _12724_);
  and (_16967_, _16865_, _03036_);
  and (_16968_, _16967_, _16966_);
  or (_16969_, _16873_, _12724_);
  and (_16971_, _16865_, _03127_);
  and (_16972_, _16971_, _16969_);
  or (_16973_, _16972_, _03166_);
  or (_16974_, _16973_, _16968_);
  or (_16975_, _16974_, _16965_);
  or (_16976_, _16870_, _03563_);
  and (_16977_, _16976_, _02501_);
  and (_16978_, _16977_, _16975_);
  and (_16979_, _16899_, _02500_);
  or (_16980_, _16979_, _03174_);
  or (_16982_, _16980_, _16978_);
  or (_16983_, _16888_, _03178_);
  or (_16984_, _16983_, _16868_);
  and (_16985_, _16984_, _34698_);
  and (_16986_, _16985_, _16982_);
  or (_35205_, _16986_, _16863_);
  not (_16987_, \oc8051_golden_model_1.P0 [2]);
  nor (_16988_, _34698_, _16987_);
  or (_16989_, _16988_, rst);
  nor (_16990_, _04716_, _16987_);
  and (_16992_, _10831_, _04716_);
  or (_16993_, _16992_, _16990_);
  and (_16994_, _16993_, _03130_);
  nor (_16995_, _08424_, _04440_);
  or (_16996_, _16995_, _16990_);
  or (_16997_, _16996_, _06241_);
  and (_16998_, _16996_, _02947_);
  nor (_16999_, _04629_, _16987_);
  and (_17000_, _10853_, _04629_);
  or (_17001_, _17000_, _16999_);
  or (_17003_, _17001_, _02892_);
  nor (_17004_, _10849_, _08424_);
  or (_17005_, _17004_, _16990_);
  and (_17006_, _17005_, _02952_);
  nor (_17007_, _03825_, _16987_);
  and (_17008_, _04716_, \oc8051_golden_model_1.ACC [2]);
  or (_17009_, _17008_, _16990_);
  and (_17010_, _17009_, _03825_);
  or (_17011_, _17010_, _17007_);
  and (_17012_, _17011_, _03821_);
  or (_17014_, _17012_, _02891_);
  or (_17015_, _17014_, _17006_);
  and (_17016_, _17015_, _17003_);
  and (_17017_, _17016_, _03327_);
  or (_17018_, _17017_, _16998_);
  or (_17019_, _17018_, _02950_);
  or (_17020_, _17009_, _02959_);
  and (_17021_, _17020_, _02888_);
  and (_17022_, _17021_, _17019_);
  and (_17023_, _10838_, _04629_);
  or (_17025_, _17023_, _16999_);
  and (_17026_, _17025_, _02887_);
  or (_17027_, _17026_, _02880_);
  or (_17028_, _17027_, _17022_);
  or (_17029_, _16999_, _10868_);
  and (_17030_, _17029_, _17001_);
  or (_17031_, _17030_, _02881_);
  and (_17032_, _17031_, _02875_);
  and (_17033_, _17032_, _17028_);
  or (_17034_, _10885_, _10838_);
  and (_17036_, _17034_, _04629_);
  or (_17037_, _17036_, _16999_);
  and (_17038_, _17037_, _02874_);
  or (_17039_, _17038_, _06793_);
  or (_17040_, _17039_, _17033_);
  and (_17041_, _17040_, _16997_);
  or (_17042_, _17041_, _02855_);
  and (_17043_, _06177_, _04716_);
  or (_17044_, _16990_, _02856_);
  or (_17045_, _17044_, _17043_);
  and (_17047_, _17045_, _02851_);
  and (_17048_, _17047_, _17042_);
  and (_17049_, _05736_, \oc8051_golden_model_1.P0 [2]);
  and (_17050_, _05733_, \oc8051_golden_model_1.P1 [2]);
  and (_17051_, _05739_, \oc8051_golden_model_1.P2 [2]);
  and (_17052_, _05741_, \oc8051_golden_model_1.P3 [2]);
  or (_17053_, _17052_, _17051_);
  or (_17054_, _17053_, _17050_);
  nor (_17055_, _17054_, _17049_);
  and (_17056_, _17055_, _10904_);
  and (_17058_, _17056_, _10925_);
  nand (_17059_, _17058_, _10941_);
  or (_17060_, _17059_, _10898_);
  and (_17061_, _17060_, _04716_);
  or (_17062_, _17061_, _16990_);
  and (_17063_, _17062_, _02576_);
  or (_17064_, _17063_, _03014_);
  or (_17065_, _17064_, _17048_);
  and (_17066_, _04716_, _05727_);
  or (_17067_, _17066_, _16990_);
  or (_17069_, _17067_, _03884_);
  and (_17070_, _17069_, _17065_);
  or (_17071_, _17070_, _03021_);
  and (_17072_, _10835_, _04716_);
  or (_17073_, _16990_, _05279_);
  or (_17074_, _17073_, _17072_);
  and (_17075_, _17074_, _03131_);
  and (_17076_, _17075_, _17071_);
  or (_17077_, _17076_, _16994_);
  and (_17078_, _17077_, _05274_);
  or (_17080_, _16990_, _05143_);
  and (_17081_, _17067_, _03020_);
  and (_17082_, _17081_, _17080_);
  or (_17083_, _17082_, _17078_);
  and (_17084_, _17083_, _03140_);
  and (_17085_, _17009_, _03139_);
  and (_17086_, _17085_, _17080_);
  or (_17087_, _17086_, _03036_);
  or (_17088_, _17087_, _17084_);
  nor (_17089_, _10833_, _08424_);
  or (_17091_, _16990_, _05781_);
  or (_17092_, _17091_, _17089_);
  and (_17093_, _17092_, _05786_);
  and (_17094_, _17093_, _17088_);
  nor (_17095_, _10830_, _08424_);
  or (_17096_, _17095_, _16990_);
  and (_17097_, _17096_, _03127_);
  or (_17098_, _17097_, _03166_);
  or (_17099_, _17098_, _17094_);
  or (_17100_, _17005_, _03563_);
  and (_17102_, _17100_, _02501_);
  and (_17103_, _17102_, _17099_);
  and (_17104_, _17025_, _02500_);
  or (_17105_, _17104_, _03174_);
  or (_17106_, _17105_, _17103_);
  and (_17107_, _11008_, _04716_);
  or (_17108_, _16990_, _03178_);
  or (_17109_, _17108_, _17107_);
  and (_17110_, _17109_, _34698_);
  and (_17111_, _17110_, _17106_);
  or (_35206_, _17111_, _16989_);
  not (_17113_, \oc8051_golden_model_1.P0 [3]);
  nor (_17114_, _34698_, _17113_);
  or (_17115_, _17114_, rst);
  nor (_17116_, _04716_, _17113_);
  and (_17117_, _11028_, _04716_);
  or (_17118_, _17117_, _17116_);
  and (_17119_, _17118_, _03130_);
  nor (_17120_, _08424_, _04242_);
  or (_17121_, _17120_, _17116_);
  or (_17123_, _17121_, _06241_);
  nor (_17124_, _11040_, _08424_);
  or (_17125_, _17124_, _17116_);
  or (_17126_, _17125_, _03821_);
  and (_17127_, _04716_, \oc8051_golden_model_1.ACC [3]);
  or (_17128_, _17127_, _17116_);
  and (_17129_, _17128_, _03825_);
  nor (_17130_, _03825_, _17113_);
  or (_17131_, _17130_, _02952_);
  or (_17132_, _17131_, _17129_);
  and (_17134_, _17132_, _02892_);
  and (_17135_, _17134_, _17126_);
  nor (_17136_, _04629_, _17113_);
  and (_17137_, _11037_, _04629_);
  or (_17138_, _17137_, _17136_);
  and (_17139_, _17138_, _02891_);
  or (_17140_, _17139_, _02947_);
  or (_17141_, _17140_, _17135_);
  or (_17142_, _17121_, _03327_);
  and (_17143_, _17142_, _17141_);
  or (_17145_, _17143_, _02950_);
  or (_17146_, _17128_, _02959_);
  and (_17147_, _17146_, _02888_);
  and (_17148_, _17147_, _17145_);
  and (_17149_, _11035_, _04629_);
  or (_17150_, _17149_, _17136_);
  and (_17151_, _17150_, _02887_);
  or (_17152_, _17151_, _02880_);
  or (_17153_, _17152_, _17148_);
  or (_17154_, _17136_, _11066_);
  and (_17156_, _17154_, _17138_);
  or (_17157_, _17156_, _02881_);
  and (_17158_, _17157_, _02875_);
  and (_17159_, _17158_, _17153_);
  or (_17160_, _11035_, _11081_);
  and (_17161_, _17160_, _04629_);
  or (_17162_, _17161_, _17136_);
  and (_17163_, _17162_, _02874_);
  or (_17164_, _17163_, _06793_);
  or (_17165_, _17164_, _17159_);
  and (_17167_, _17165_, _17123_);
  or (_17168_, _17167_, _02855_);
  and (_17169_, _06176_, _04716_);
  or (_17170_, _17116_, _02856_);
  or (_17171_, _17170_, _17169_);
  and (_17172_, _17171_, _02851_);
  and (_17173_, _17172_, _17168_);
  and (_17174_, _05733_, \oc8051_golden_model_1.P1 [3]);
  and (_17175_, _05736_, \oc8051_golden_model_1.P0 [3]);
  and (_17176_, _05739_, \oc8051_golden_model_1.P2 [3]);
  and (_17178_, _05741_, \oc8051_golden_model_1.P3 [3]);
  or (_17179_, _17178_, _17176_);
  or (_17180_, _17179_, _17175_);
  nor (_17181_, _17180_, _17174_);
  and (_17182_, _17181_, _11109_);
  and (_17183_, _17182_, _11104_);
  nand (_17184_, _17183_, _11141_);
  or (_17185_, _17184_, _11096_);
  and (_17186_, _17185_, _04716_);
  or (_17187_, _17186_, _17116_);
  and (_17189_, _17187_, _02576_);
  or (_17190_, _17189_, _03014_);
  or (_17191_, _17190_, _17173_);
  and (_17192_, _04716_, _05664_);
  or (_17193_, _17192_, _17116_);
  or (_17194_, _17193_, _03884_);
  and (_17195_, _17194_, _17191_);
  or (_17196_, _17195_, _03021_);
  and (_17197_, _11032_, _04716_);
  or (_17198_, _17116_, _05279_);
  or (_17200_, _17198_, _17197_);
  and (_17201_, _17200_, _03131_);
  and (_17202_, _17201_, _17196_);
  or (_17203_, _17202_, _17119_);
  and (_17204_, _17203_, _05274_);
  or (_17205_, _17116_, _04996_);
  and (_17206_, _17193_, _03020_);
  and (_17207_, _17206_, _17205_);
  or (_17208_, _17207_, _17204_);
  and (_17209_, _17208_, _03140_);
  and (_17211_, _17128_, _03139_);
  and (_17212_, _17211_, _17205_);
  or (_17213_, _17212_, _03036_);
  or (_17214_, _17213_, _17209_);
  nor (_17215_, _11030_, _08424_);
  or (_17216_, _17116_, _05781_);
  or (_17217_, _17216_, _17215_);
  and (_17218_, _17217_, _05786_);
  and (_17219_, _17218_, _17214_);
  nor (_17220_, _11027_, _08424_);
  or (_17222_, _17220_, _17116_);
  and (_17223_, _17222_, _03127_);
  or (_17224_, _17223_, _03166_);
  or (_17225_, _17224_, _17219_);
  or (_17226_, _17125_, _03563_);
  and (_17227_, _17226_, _02501_);
  and (_17228_, _17227_, _17225_);
  and (_17229_, _17150_, _02500_);
  or (_17230_, _17229_, _03174_);
  or (_17231_, _17230_, _17228_);
  and (_17233_, _11213_, _04716_);
  or (_17234_, _17116_, _03178_);
  or (_17235_, _17234_, _17233_);
  and (_17236_, _17235_, _34698_);
  and (_17237_, _17236_, _17231_);
  or (_35208_, _17237_, _17115_);
  not (_17238_, \oc8051_golden_model_1.P0 [4]);
  nor (_17239_, _34698_, _17238_);
  or (_17240_, _17239_, rst);
  nor (_17241_, _04716_, _17238_);
  and (_17243_, _11368_, _04716_);
  or (_17244_, _17243_, _17241_);
  and (_17245_, _17244_, _03130_);
  nor (_17246_, _05202_, _08424_);
  or (_17247_, _17246_, _17241_);
  or (_17248_, _17247_, _06241_);
  nor (_17249_, _04629_, _17238_);
  and (_17250_, _11243_, _04629_);
  or (_17251_, _17250_, _17249_);
  and (_17252_, _17251_, _02887_);
  nor (_17254_, _11259_, _08424_);
  or (_17255_, _17254_, _17241_);
  or (_17256_, _17255_, _03821_);
  and (_17257_, _04716_, \oc8051_golden_model_1.ACC [4]);
  or (_17258_, _17257_, _17241_);
  and (_17259_, _17258_, _03825_);
  nor (_17260_, _03825_, _17238_);
  or (_17261_, _17260_, _02952_);
  or (_17262_, _17261_, _17259_);
  and (_17263_, _17262_, _02892_);
  and (_17265_, _17263_, _17256_);
  and (_17266_, _11245_, _04629_);
  or (_17267_, _17266_, _17249_);
  and (_17268_, _17267_, _02891_);
  or (_17269_, _17268_, _02947_);
  or (_17270_, _17269_, _17265_);
  or (_17271_, _17247_, _03327_);
  and (_17272_, _17271_, _17270_);
  or (_17273_, _17272_, _02950_);
  or (_17274_, _17258_, _02959_);
  and (_17276_, _17274_, _02888_);
  and (_17277_, _17276_, _17273_);
  or (_17278_, _17277_, _17252_);
  and (_17279_, _17278_, _02881_);
  or (_17280_, _17249_, _11276_);
  and (_17281_, _17280_, _02880_);
  and (_17282_, _17281_, _17267_);
  or (_17283_, _17282_, _17279_);
  and (_17284_, _17283_, _02875_);
  or (_17285_, _11243_, _11240_);
  and (_17287_, _17285_, _04629_);
  or (_17288_, _17287_, _17249_);
  and (_17289_, _17288_, _02874_);
  or (_17290_, _17289_, _06793_);
  or (_17291_, _17290_, _17284_);
  and (_17292_, _17291_, _17248_);
  or (_17293_, _17292_, _02855_);
  and (_17294_, _06181_, _04716_);
  or (_17295_, _17241_, _02856_);
  or (_17296_, _17295_, _17294_);
  and (_17298_, _17296_, _02851_);
  and (_17299_, _17298_, _17293_);
  and (_17300_, _05736_, \oc8051_golden_model_1.P0 [4]);
  and (_17301_, _05733_, \oc8051_golden_model_1.P1 [4]);
  and (_17302_, _05739_, \oc8051_golden_model_1.P2 [4]);
  and (_17303_, _05741_, \oc8051_golden_model_1.P3 [4]);
  or (_17304_, _17303_, _17302_);
  or (_17305_, _17304_, _17301_);
  nor (_17306_, _17305_, _17300_);
  and (_17307_, _17306_, _11344_);
  and (_17309_, _17307_, _11332_);
  nand (_17310_, _17309_, _11325_);
  or (_17311_, _17310_, _11303_);
  and (_17312_, _17311_, _04716_);
  or (_17313_, _17312_, _17241_);
  and (_17314_, _17313_, _02576_);
  or (_17315_, _17314_, _03014_);
  or (_17316_, _17315_, _17299_);
  and (_17317_, _05697_, _04716_);
  or (_17318_, _17317_, _17241_);
  or (_17320_, _17318_, _03884_);
  and (_17321_, _17320_, _17316_);
  or (_17322_, _17321_, _03021_);
  and (_17323_, _11362_, _04716_);
  or (_17324_, _17241_, _05279_);
  or (_17325_, _17324_, _17323_);
  and (_17326_, _17325_, _03131_);
  and (_17327_, _17326_, _17322_);
  or (_17328_, _17327_, _17245_);
  and (_17329_, _17328_, _05274_);
  or (_17331_, _17241_, _05251_);
  and (_17332_, _17318_, _03020_);
  and (_17333_, _17332_, _17331_);
  or (_17334_, _17333_, _17329_);
  and (_17335_, _17334_, _03140_);
  and (_17336_, _17258_, _03139_);
  and (_17337_, _17336_, _17331_);
  or (_17338_, _17337_, _03036_);
  or (_17339_, _17338_, _17335_);
  nor (_17340_, _11361_, _08424_);
  or (_17342_, _17241_, _05781_);
  or (_17343_, _17342_, _17340_);
  and (_17344_, _17343_, _05786_);
  and (_17345_, _17344_, _17339_);
  nor (_17346_, _11367_, _08424_);
  or (_17347_, _17346_, _17241_);
  and (_17348_, _17347_, _03127_);
  or (_17349_, _17348_, _03166_);
  or (_17350_, _17349_, _17345_);
  or (_17351_, _17255_, _03563_);
  and (_17353_, _17351_, _02501_);
  and (_17354_, _17353_, _17350_);
  and (_17355_, _17251_, _02500_);
  or (_17356_, _17355_, _03174_);
  or (_17357_, _17356_, _17354_);
  and (_17358_, _11417_, _04716_);
  or (_17359_, _17241_, _03178_);
  or (_17360_, _17359_, _17358_);
  and (_17361_, _17360_, _34698_);
  and (_17362_, _17361_, _17357_);
  or (_35209_, _17362_, _17240_);
  not (_17364_, \oc8051_golden_model_1.P0 [5]);
  nor (_17365_, _34698_, _17364_);
  or (_17366_, _17365_, rst);
  nor (_17367_, _04716_, _17364_);
  and (_17368_, _11436_, _04716_);
  or (_17369_, _17368_, _17367_);
  and (_17370_, _17369_, _03130_);
  nor (_17371_, _11445_, _08424_);
  or (_17372_, _17371_, _17367_);
  or (_17374_, _17372_, _03821_);
  and (_17375_, _04716_, \oc8051_golden_model_1.ACC [5]);
  or (_17376_, _17375_, _17367_);
  and (_17377_, _17376_, _03825_);
  nor (_17378_, _03825_, _17364_);
  or (_17379_, _17378_, _02952_);
  or (_17380_, _17379_, _17377_);
  and (_17381_, _17380_, _02892_);
  and (_17382_, _17381_, _17374_);
  nor (_17383_, _04629_, _17364_);
  and (_17384_, _11459_, _04629_);
  or (_17385_, _17384_, _17383_);
  and (_17386_, _17385_, _02891_);
  or (_17387_, _17386_, _02947_);
  or (_17388_, _17387_, _17382_);
  nor (_17389_, _04896_, _08424_);
  or (_17390_, _17389_, _17367_);
  or (_17391_, _17390_, _03327_);
  and (_17392_, _17391_, _17388_);
  or (_17393_, _17392_, _02950_);
  or (_17396_, _17376_, _02959_);
  and (_17397_, _17396_, _02888_);
  and (_17398_, _17397_, _17393_);
  and (_17399_, _11442_, _04629_);
  or (_17400_, _17399_, _17383_);
  and (_17401_, _17400_, _02887_);
  or (_17402_, _17401_, _02880_);
  or (_17403_, _17402_, _17398_);
  or (_17404_, _17383_, _11474_);
  and (_17405_, _17404_, _17385_);
  or (_17406_, _17405_, _02881_);
  and (_17407_, _17406_, _02875_);
  and (_17408_, _17407_, _17403_);
  or (_17409_, _11442_, _11439_);
  and (_17410_, _17409_, _04629_);
  or (_17411_, _17410_, _17383_);
  and (_17412_, _17411_, _02874_);
  or (_17413_, _17412_, _06793_);
  or (_17414_, _17413_, _17408_);
  or (_17415_, _17390_, _06241_);
  and (_17418_, _17415_, _17414_);
  or (_17419_, _17418_, _02855_);
  and (_17420_, _06180_, _04716_);
  or (_17421_, _17367_, _02856_);
  or (_17422_, _17421_, _17420_);
  and (_17423_, _17422_, _02851_);
  and (_17424_, _17423_, _17419_);
  and (_17425_, _05736_, \oc8051_golden_model_1.P0 [5]);
  and (_17426_, _05733_, \oc8051_golden_model_1.P1 [5]);
  and (_17427_, _05739_, \oc8051_golden_model_1.P2 [5]);
  and (_17429_, _05741_, \oc8051_golden_model_1.P3 [5]);
  or (_17430_, _17429_, _17427_);
  or (_17431_, _17430_, _17426_);
  nor (_17432_, _17431_, _17425_);
  and (_17433_, _17432_, _11542_);
  and (_17434_, _17433_, _11530_);
  nand (_17435_, _17434_, _11523_);
  or (_17436_, _17435_, _11501_);
  and (_17437_, _17436_, _04716_);
  or (_17438_, _17437_, _17367_);
  and (_17440_, _17438_, _02576_);
  or (_17441_, _17440_, _03014_);
  or (_17442_, _17441_, _17424_);
  and (_17443_, _05701_, _04716_);
  or (_17444_, _17443_, _17367_);
  or (_17445_, _17444_, _03884_);
  and (_17446_, _17445_, _17442_);
  or (_17447_, _17446_, _03021_);
  and (_17448_, _11562_, _04716_);
  or (_17449_, _17367_, _05279_);
  or (_17451_, _17449_, _17448_);
  and (_17452_, _17451_, _03131_);
  and (_17453_, _17452_, _17447_);
  or (_17454_, _17453_, _17370_);
  and (_17455_, _17454_, _05274_);
  or (_17456_, _17367_, _04944_);
  and (_17457_, _17444_, _03020_);
  and (_17458_, _17457_, _17456_);
  or (_17459_, _17458_, _17455_);
  and (_17460_, _17459_, _03140_);
  and (_17462_, _17376_, _03139_);
  and (_17463_, _17462_, _17456_);
  or (_17464_, _17463_, _03036_);
  or (_17465_, _17464_, _17460_);
  nor (_17466_, _11560_, _08424_);
  or (_17467_, _17367_, _05781_);
  or (_17468_, _17467_, _17466_);
  and (_17469_, _17468_, _05786_);
  and (_17470_, _17469_, _17465_);
  nor (_17471_, _11435_, _08424_);
  or (_17473_, _17471_, _17367_);
  and (_17474_, _17473_, _03127_);
  or (_17475_, _17474_, _03166_);
  or (_17476_, _17475_, _17470_);
  or (_17477_, _17372_, _03563_);
  and (_17478_, _17477_, _02501_);
  and (_17479_, _17478_, _17476_);
  and (_17480_, _17400_, _02500_);
  or (_17481_, _17480_, _03174_);
  or (_17482_, _17481_, _17479_);
  and (_17484_, _11619_, _04716_);
  or (_17485_, _17367_, _03178_);
  or (_17486_, _17485_, _17484_);
  and (_17487_, _17486_, _34698_);
  and (_17488_, _17487_, _17482_);
  or (_35210_, _17488_, _17366_);
  not (_17489_, \oc8051_golden_model_1.P0 [6]);
  nor (_17490_, _34698_, _17489_);
  or (_17491_, _17490_, rst);
  nor (_17492_, _04716_, _17489_);
  and (_17494_, _11769_, _04716_);
  or (_17495_, _17494_, _17492_);
  and (_17496_, _17495_, _03130_);
  nor (_17497_, _11636_, _08424_);
  or (_17498_, _17497_, _17492_);
  or (_17499_, _17498_, _03821_);
  and (_17500_, _04716_, \oc8051_golden_model_1.ACC [6]);
  or (_17501_, _17500_, _17492_);
  and (_17502_, _17501_, _03825_);
  nor (_17503_, _03825_, _17489_);
  or (_17505_, _17503_, _02952_);
  or (_17506_, _17505_, _17502_);
  and (_17507_, _17506_, _02892_);
  and (_17508_, _17507_, _17499_);
  nor (_17509_, _04629_, _17489_);
  and (_17510_, _11653_, _04629_);
  or (_17511_, _17510_, _17509_);
  and (_17512_, _17511_, _02891_);
  or (_17513_, _17512_, _02947_);
  or (_17514_, _17513_, _17508_);
  nor (_17516_, _04787_, _08424_);
  or (_17517_, _17516_, _17492_);
  or (_17518_, _17517_, _03327_);
  and (_17519_, _17518_, _17514_);
  or (_17520_, _17519_, _02950_);
  or (_17521_, _17501_, _02959_);
  and (_17522_, _17521_, _02888_);
  and (_17523_, _17522_, _17520_);
  and (_17524_, _11675_, _04629_);
  or (_17525_, _17524_, _17509_);
  and (_17527_, _17525_, _02887_);
  or (_17528_, _17527_, _02880_);
  or (_17529_, _17528_, _17523_);
  or (_17530_, _17509_, _11682_);
  and (_17531_, _17530_, _17511_);
  or (_17532_, _17531_, _02881_);
  and (_17533_, _17532_, _02875_);
  and (_17534_, _17533_, _17529_);
  or (_17535_, _11675_, _11649_);
  and (_17536_, _17535_, _04629_);
  or (_17538_, _17536_, _17509_);
  and (_17539_, _17538_, _02874_);
  or (_17540_, _17539_, _06793_);
  or (_17541_, _17540_, _17534_);
  or (_17542_, _17517_, _06241_);
  and (_17543_, _17542_, _17541_);
  or (_17544_, _17543_, _02855_);
  and (_17545_, _05847_, _04716_);
  or (_17546_, _17492_, _02856_);
  or (_17547_, _17546_, _17545_);
  and (_17549_, _17547_, _02851_);
  and (_17550_, _17549_, _17544_);
  and (_17551_, _05733_, \oc8051_golden_model_1.P1 [6]);
  and (_17552_, _05736_, \oc8051_golden_model_1.P0 [6]);
  and (_17553_, _05739_, \oc8051_golden_model_1.P2 [6]);
  and (_17554_, _05741_, \oc8051_golden_model_1.P3 [6]);
  or (_17555_, _17554_, _17553_);
  or (_17556_, _17555_, _17552_);
  or (_17557_, _17556_, _17551_);
  or (_17558_, _17557_, _11746_);
  or (_17560_, _17558_, _11736_);
  or (_17561_, _17560_, _11731_);
  or (_17562_, _17561_, _11724_);
  or (_17563_, _17562_, _11709_);
  and (_17564_, _17563_, _04716_);
  or (_17565_, _17564_, _17492_);
  and (_17566_, _17565_, _02576_);
  or (_17567_, _17566_, _03014_);
  or (_17568_, _17567_, _17550_);
  and (_17569_, _11758_, _04716_);
  or (_17571_, _17569_, _17492_);
  or (_17572_, _17571_, _03884_);
  and (_17573_, _17572_, _17568_);
  or (_17574_, _17573_, _03021_);
  and (_17575_, _11646_, _04716_);
  or (_17576_, _17492_, _05279_);
  or (_17577_, _17576_, _17575_);
  and (_17578_, _17577_, _03131_);
  and (_17579_, _17578_, _17574_);
  or (_17580_, _17579_, _17496_);
  and (_17582_, _17580_, _05274_);
  or (_17583_, _17492_, _04838_);
  and (_17584_, _17571_, _03020_);
  and (_17585_, _17584_, _17583_);
  or (_17586_, _17585_, _17582_);
  and (_17587_, _17586_, _03140_);
  and (_17588_, _17501_, _03139_);
  and (_17589_, _17588_, _17583_);
  or (_17590_, _17589_, _03036_);
  or (_17591_, _17590_, _17587_);
  nor (_17593_, _11644_, _08424_);
  or (_17594_, _17492_, _05781_);
  or (_17595_, _17594_, _17593_);
  and (_17596_, _17595_, _05786_);
  and (_17597_, _17596_, _17591_);
  nor (_17598_, _11768_, _08424_);
  or (_17599_, _17598_, _17492_);
  and (_17600_, _17599_, _03127_);
  or (_17601_, _17600_, _03166_);
  or (_17602_, _17601_, _17597_);
  or (_17604_, _17498_, _03563_);
  and (_17605_, _17604_, _02501_);
  and (_17606_, _17605_, _17602_);
  and (_17607_, _17525_, _02500_);
  or (_17608_, _17607_, _03174_);
  or (_17609_, _17608_, _17606_);
  and (_17610_, _11821_, _04716_);
  or (_17611_, _17492_, _03178_);
  or (_17612_, _17611_, _17610_);
  and (_17613_, _17612_, _34698_);
  and (_17615_, _17613_, _17609_);
  or (_35211_, _17615_, _17491_);
  not (_17616_, \oc8051_golden_model_1.P1 [0]);
  nor (_17617_, _34698_, _17616_);
  or (_17618_, _17617_, rst);
  nor (_17619_, _04719_, _17616_);
  and (_17620_, _10546_, _04719_);
  or (_17621_, _17620_, _17619_);
  and (_17622_, _17621_, _03130_);
  and (_17623_, _04719_, _03817_);
  or (_17625_, _17623_, _17619_);
  or (_17626_, _17625_, _06241_);
  and (_17627_, _05044_, _04719_);
  or (_17628_, _17627_, _17619_);
  or (_17629_, _17628_, _03821_);
  and (_17630_, _04719_, \oc8051_golden_model_1.ACC [0]);
  or (_17631_, _17630_, _17619_);
  and (_17632_, _17631_, _03825_);
  nor (_17633_, _03825_, _17616_);
  or (_17634_, _17633_, _02952_);
  or (_17636_, _17634_, _17632_);
  and (_17637_, _17636_, _02892_);
  and (_17638_, _17637_, _17629_);
  nor (_17639_, _05344_, _17616_);
  and (_17640_, _10429_, _05344_);
  or (_17641_, _17640_, _17639_);
  and (_17642_, _17641_, _02891_);
  or (_17643_, _17642_, _17638_);
  and (_17644_, _17643_, _03327_);
  and (_17645_, _17625_, _02947_);
  or (_17647_, _17645_, _02950_);
  or (_17648_, _17647_, _17644_);
  or (_17649_, _17631_, _02959_);
  and (_17650_, _17649_, _02888_);
  and (_17651_, _17650_, _17648_);
  and (_17652_, _17619_, _02887_);
  or (_17653_, _17652_, _02880_);
  or (_17654_, _17653_, _17651_);
  or (_17655_, _17628_, _02881_);
  and (_17656_, _17655_, _02875_);
  and (_17658_, _17656_, _17654_);
  and (_17659_, _16789_, _05344_);
  or (_17660_, _17659_, _17639_);
  and (_17661_, _17660_, _02874_);
  or (_17662_, _17661_, _06793_);
  or (_17663_, _17662_, _17658_);
  and (_17664_, _17663_, _17626_);
  or (_17665_, _17664_, _02855_);
  and (_17666_, _06174_, _04719_);
  or (_17667_, _17619_, _02856_);
  or (_17669_, _17667_, _17666_);
  and (_17670_, _17669_, _02851_);
  and (_17671_, _17670_, _17665_);
  and (_17672_, _16814_, _04719_);
  or (_17673_, _17672_, _17619_);
  and (_17674_, _17673_, _02576_);
  or (_17675_, _17674_, _03014_);
  or (_17676_, _17675_, _17671_);
  and (_17677_, _04719_, _05566_);
  or (_17678_, _17677_, _17619_);
  or (_17680_, _17678_, _03884_);
  and (_17681_, _17680_, _17676_);
  or (_17682_, _17681_, _03021_);
  and (_17683_, _10425_, _04719_);
  or (_17684_, _17619_, _05279_);
  or (_17685_, _17684_, _17683_);
  and (_17686_, _17685_, _03131_);
  and (_17687_, _17686_, _17682_);
  or (_17688_, _17687_, _17622_);
  and (_17689_, _17688_, _05274_);
  nand (_17691_, _17678_, _03020_);
  nor (_17692_, _17691_, _17627_);
  or (_17693_, _17692_, _17689_);
  and (_17694_, _17693_, _03140_);
  or (_17695_, _17619_, _09183_);
  and (_17696_, _17631_, _03139_);
  and (_17697_, _17696_, _17695_);
  or (_17698_, _17697_, _03036_);
  or (_17699_, _17698_, _17694_);
  nor (_17700_, _10423_, _08539_);
  or (_17702_, _17619_, _05781_);
  or (_17703_, _17702_, _17700_);
  and (_17704_, _17703_, _05786_);
  and (_17705_, _17704_, _17699_);
  nor (_17706_, _10421_, _08539_);
  or (_17707_, _17706_, _17619_);
  and (_17708_, _17707_, _03127_);
  or (_17709_, _17708_, _03166_);
  or (_17710_, _17709_, _17705_);
  or (_17711_, _17628_, _03563_);
  and (_17713_, _17711_, _02501_);
  and (_17714_, _17713_, _17710_);
  and (_17715_, _17619_, _02500_);
  or (_17716_, _17715_, _03174_);
  or (_17717_, _17716_, _17714_);
  or (_17718_, _17628_, _03178_);
  and (_17719_, _17718_, _34698_);
  and (_17720_, _17719_, _17717_);
  or (_35213_, _17720_, _17618_);
  not (_17721_, \oc8051_golden_model_1.P1 [1]);
  nor (_17723_, _34698_, _17721_);
  or (_17724_, _17723_, rst);
  nand (_17725_, _04719_, _03705_);
  or (_17726_, _04719_, \oc8051_golden_model_1.P1 [1]);
  and (_17727_, _17726_, _03014_);
  and (_17728_, _17727_, _17725_);
  or (_17729_, _16935_, _08539_);
  and (_17730_, _17726_, _02576_);
  and (_17731_, _17730_, _17729_);
  and (_17732_, _10622_, _04719_);
  not (_17734_, _17732_);
  and (_17735_, _17734_, _17726_);
  or (_17736_, _17735_, _03821_);
  nand (_17737_, _04719_, _02618_);
  and (_17738_, _17737_, _17726_);
  and (_17739_, _17738_, _03825_);
  nor (_17740_, _03825_, _17721_);
  or (_17741_, _17740_, _02952_);
  or (_17742_, _17741_, _17739_);
  and (_17743_, _17742_, _02892_);
  and (_17745_, _17743_, _17736_);
  nor (_17746_, _05344_, _17721_);
  and (_17747_, _10617_, _05344_);
  or (_17748_, _17747_, _17746_);
  and (_17749_, _17748_, _02891_);
  or (_17750_, _17749_, _02947_);
  or (_17751_, _17750_, _17745_);
  nor (_17752_, _04719_, _17721_);
  and (_17753_, _04719_, _04005_);
  or (_17754_, _17753_, _17752_);
  or (_17756_, _17754_, _03327_);
  and (_17757_, _17756_, _17751_);
  or (_17758_, _17757_, _02950_);
  or (_17759_, _17738_, _02959_);
  and (_17760_, _17759_, _02888_);
  and (_17761_, _17760_, _17758_);
  and (_17762_, _10620_, _05344_);
  or (_17763_, _17762_, _17746_);
  and (_17764_, _17763_, _02887_);
  or (_17765_, _17764_, _02880_);
  or (_17767_, _17765_, _17761_);
  and (_17768_, _17747_, _10616_);
  or (_17769_, _17746_, _02881_);
  or (_17770_, _17769_, _17768_);
  and (_17771_, _17770_, _17767_);
  and (_17772_, _17771_, _02875_);
  and (_17773_, _16909_, _05344_);
  or (_17774_, _17746_, _17773_);
  and (_17775_, _17774_, _02874_);
  or (_17776_, _17775_, _06793_);
  or (_17778_, _17776_, _17772_);
  or (_17779_, _17754_, _06241_);
  and (_17780_, _17779_, _17778_);
  or (_17781_, _17780_, _02855_);
  and (_17782_, _06173_, _04719_);
  or (_17783_, _17752_, _02856_);
  or (_17784_, _17783_, _17782_);
  and (_17785_, _17784_, _02851_);
  and (_17786_, _17785_, _17781_);
  or (_17787_, _17786_, _17731_);
  and (_17789_, _17787_, _03884_);
  or (_17790_, _17789_, _17728_);
  and (_17791_, _17790_, _05279_);
  or (_17792_, _10612_, _08539_);
  and (_17793_, _17726_, _03021_);
  and (_17794_, _17793_, _17792_);
  or (_17795_, _17794_, _17791_);
  and (_17796_, _17795_, _03131_);
  or (_17797_, _10739_, _08539_);
  and (_17798_, _17726_, _03130_);
  and (_17800_, _17798_, _17797_);
  or (_17801_, _17800_, _17796_);
  and (_17802_, _17801_, _05274_);
  or (_17803_, _10611_, _08539_);
  and (_17804_, _17726_, _03020_);
  and (_17805_, _17804_, _17803_);
  or (_17806_, _17805_, _17802_);
  and (_17807_, _17806_, _03140_);
  or (_17808_, _17752_, _12724_);
  and (_17809_, _17738_, _03139_);
  and (_17811_, _17809_, _17808_);
  or (_17812_, _17811_, _17807_);
  and (_17813_, _17812_, _03128_);
  or (_17814_, _17725_, _12724_);
  and (_17815_, _17726_, _03036_);
  and (_17816_, _17815_, _17814_);
  or (_17817_, _17737_, _12724_);
  and (_17818_, _17726_, _03127_);
  and (_17819_, _17818_, _17817_);
  or (_17820_, _17819_, _03166_);
  or (_17822_, _17820_, _17816_);
  or (_17823_, _17822_, _17813_);
  or (_17824_, _17735_, _03563_);
  and (_17825_, _17824_, _02501_);
  and (_17826_, _17825_, _17823_);
  and (_17827_, _17763_, _02500_);
  or (_17828_, _17827_, _03174_);
  or (_17829_, _17828_, _17826_);
  or (_17830_, _17752_, _03178_);
  or (_17831_, _17830_, _17732_);
  and (_17833_, _17831_, _34698_);
  and (_17834_, _17833_, _17829_);
  or (_35214_, _17834_, _17724_);
  not (_17835_, \oc8051_golden_model_1.P1 [2]);
  nor (_17836_, _34698_, _17835_);
  or (_17837_, _17836_, rst);
  nor (_17838_, _04719_, _17835_);
  and (_17839_, _10831_, _04719_);
  or (_17840_, _17839_, _17838_);
  and (_17841_, _17840_, _03130_);
  nor (_17843_, _08539_, _04440_);
  or (_17844_, _17843_, _17838_);
  or (_17845_, _17844_, _06241_);
  or (_17846_, _17844_, _03327_);
  nor (_17847_, _10849_, _08539_);
  or (_17848_, _17847_, _17838_);
  or (_17849_, _17848_, _03821_);
  and (_17850_, _04719_, \oc8051_golden_model_1.ACC [2]);
  or (_17851_, _17850_, _17838_);
  and (_17852_, _17851_, _03825_);
  nor (_17854_, _03825_, _17835_);
  or (_17855_, _17854_, _02952_);
  or (_17856_, _17855_, _17852_);
  and (_17857_, _17856_, _02892_);
  and (_17858_, _17857_, _17849_);
  nor (_17859_, _05344_, _17835_);
  and (_17860_, _10853_, _05344_);
  or (_17861_, _17860_, _17859_);
  and (_17862_, _17861_, _02891_);
  or (_17863_, _17862_, _02947_);
  or (_17865_, _17863_, _17858_);
  and (_17866_, _17865_, _17846_);
  or (_17867_, _17866_, _02950_);
  or (_17868_, _17851_, _02959_);
  and (_17869_, _17868_, _02888_);
  and (_17870_, _17869_, _17867_);
  and (_17871_, _10838_, _05344_);
  or (_17872_, _17871_, _17859_);
  and (_17873_, _17872_, _02887_);
  or (_17874_, _17873_, _02880_);
  or (_17876_, _17874_, _17870_);
  and (_17877_, _17860_, _10868_);
  or (_17878_, _17859_, _02881_);
  or (_17879_, _17878_, _17877_);
  and (_17880_, _17879_, _02875_);
  and (_17881_, _17880_, _17876_);
  and (_17882_, _17034_, _05344_);
  or (_17883_, _17882_, _17859_);
  and (_17884_, _17883_, _02874_);
  or (_17885_, _17884_, _06793_);
  or (_17887_, _17885_, _17881_);
  and (_17888_, _17887_, _17845_);
  or (_17889_, _17888_, _02855_);
  and (_17890_, _06177_, _04719_);
  or (_17891_, _17838_, _02856_);
  or (_17892_, _17891_, _17890_);
  and (_17893_, _17892_, _02851_);
  and (_17894_, _17893_, _17889_);
  and (_17895_, _17060_, _04719_);
  or (_17896_, _17895_, _17838_);
  and (_17898_, _17896_, _02576_);
  or (_17899_, _17898_, _03014_);
  or (_17900_, _17899_, _17894_);
  and (_17901_, _04719_, _05727_);
  or (_17902_, _17901_, _17838_);
  or (_17903_, _17902_, _03884_);
  and (_17904_, _17903_, _17900_);
  or (_17905_, _17904_, _03021_);
  and (_17906_, _10835_, _04719_);
  or (_17907_, _17838_, _05279_);
  or (_17909_, _17907_, _17906_);
  and (_17910_, _17909_, _03131_);
  and (_17911_, _17910_, _17905_);
  or (_17912_, _17911_, _17841_);
  and (_17913_, _17912_, _05274_);
  or (_17914_, _17838_, _05143_);
  and (_17915_, _17902_, _03020_);
  and (_17916_, _17915_, _17914_);
  or (_17917_, _17916_, _17913_);
  and (_17918_, _17917_, _03140_);
  and (_17920_, _17851_, _03139_);
  and (_17921_, _17920_, _17914_);
  or (_17922_, _17921_, _03036_);
  or (_17923_, _17922_, _17918_);
  nor (_17924_, _10833_, _08539_);
  or (_17925_, _17838_, _05781_);
  or (_17926_, _17925_, _17924_);
  and (_17927_, _17926_, _05786_);
  and (_17928_, _17927_, _17923_);
  nor (_17929_, _10830_, _08539_);
  or (_17931_, _17929_, _17838_);
  and (_17932_, _17931_, _03127_);
  or (_17933_, _17932_, _03166_);
  or (_17934_, _17933_, _17928_);
  or (_17935_, _17848_, _03563_);
  and (_17936_, _17935_, _02501_);
  and (_17937_, _17936_, _17934_);
  and (_17938_, _17872_, _02500_);
  or (_17939_, _17938_, _03174_);
  or (_17940_, _17939_, _17937_);
  and (_17942_, _11008_, _04719_);
  or (_17943_, _17838_, _03178_);
  or (_17944_, _17943_, _17942_);
  and (_17945_, _17944_, _34698_);
  and (_17946_, _17945_, _17940_);
  or (_35215_, _17946_, _17837_);
  nor (_17947_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_17948_, _17947_, _04548_);
  and (_17949_, _08539_, \oc8051_golden_model_1.P1 [3]);
  and (_17950_, _11028_, _04719_);
  or (_17952_, _17950_, _17949_);
  and (_17953_, _17952_, _03130_);
  nor (_17954_, _08539_, _04242_);
  or (_17955_, _17954_, _17949_);
  or (_17956_, _17955_, _06241_);
  nor (_17957_, _11040_, _08539_);
  or (_17958_, _17957_, _17949_);
  or (_17959_, _17958_, _03821_);
  and (_17960_, _04719_, \oc8051_golden_model_1.ACC [3]);
  or (_17961_, _17960_, _17949_);
  and (_17963_, _17961_, _03825_);
  and (_17964_, _03826_, \oc8051_golden_model_1.P1 [3]);
  or (_17965_, _17964_, _02952_);
  or (_17966_, _17965_, _17963_);
  and (_17967_, _17966_, _02892_);
  and (_17968_, _17967_, _17959_);
  not (_17969_, _05344_);
  and (_17970_, _17969_, \oc8051_golden_model_1.P1 [3]);
  and (_17971_, _11037_, _05344_);
  or (_17972_, _17971_, _17970_);
  and (_17974_, _17972_, _02891_);
  or (_17975_, _17974_, _02947_);
  or (_17976_, _17975_, _17968_);
  or (_17977_, _17955_, _03327_);
  and (_17978_, _17977_, _17976_);
  or (_17979_, _17978_, _02950_);
  or (_17980_, _17961_, _02959_);
  and (_17981_, _17980_, _02888_);
  and (_17982_, _17981_, _17979_);
  and (_17983_, _11035_, _05344_);
  or (_17985_, _17983_, _17970_);
  and (_17986_, _17985_, _02887_);
  or (_17987_, _17986_, _02880_);
  or (_17988_, _17987_, _17982_);
  or (_17989_, _17970_, _11066_);
  and (_17990_, _17989_, _17972_);
  or (_17991_, _17990_, _02881_);
  and (_17992_, _17991_, _02875_);
  and (_17993_, _17992_, _17988_);
  and (_17994_, _17160_, _05344_);
  or (_17996_, _17994_, _17970_);
  and (_17997_, _17996_, _02874_);
  or (_17998_, _17997_, _06793_);
  or (_17999_, _17998_, _17993_);
  and (_18000_, _17999_, _17956_);
  or (_18001_, _18000_, _02855_);
  and (_18002_, _06176_, _04719_);
  or (_18003_, _17949_, _02856_);
  or (_18004_, _18003_, _18002_);
  and (_18005_, _18004_, _02851_);
  and (_18007_, _18005_, _18001_);
  and (_18008_, _17185_, _04719_);
  or (_18009_, _18008_, _17949_);
  and (_18010_, _18009_, _02576_);
  or (_18011_, _18010_, _03014_);
  or (_18012_, _18011_, _18007_);
  and (_18013_, _04719_, _05664_);
  or (_18014_, _18013_, _17949_);
  or (_18015_, _18014_, _03884_);
  and (_18016_, _18015_, _18012_);
  or (_18018_, _18016_, _03021_);
  and (_18019_, _11032_, _04719_);
  or (_18020_, _17949_, _05279_);
  or (_18021_, _18020_, _18019_);
  and (_18022_, _18021_, _03131_);
  and (_18023_, _18022_, _18018_);
  or (_18024_, _18023_, _17953_);
  and (_18025_, _18024_, _05274_);
  or (_18026_, _17949_, _04996_);
  and (_18027_, _18014_, _03020_);
  and (_18029_, _18027_, _18026_);
  or (_18030_, _18029_, _18025_);
  and (_18031_, _18030_, _03140_);
  and (_18032_, _17961_, _03139_);
  and (_18033_, _18032_, _18026_);
  or (_18034_, _18033_, _03036_);
  or (_18035_, _18034_, _18031_);
  nor (_18036_, _11030_, _08539_);
  or (_18037_, _17949_, _05781_);
  or (_18038_, _18037_, _18036_);
  and (_18040_, _18038_, _05786_);
  and (_18041_, _18040_, _18035_);
  nor (_18042_, _11027_, _08539_);
  or (_18043_, _18042_, _17949_);
  and (_18044_, _18043_, _03127_);
  or (_18045_, _18044_, _03166_);
  or (_18046_, _18045_, _18041_);
  or (_18047_, _17958_, _03563_);
  and (_18048_, _18047_, _02501_);
  and (_18049_, _18048_, _18046_);
  and (_18051_, _17985_, _02500_);
  or (_18052_, _18051_, _03174_);
  or (_18053_, _18052_, _18049_);
  and (_18054_, _11213_, _04719_);
  or (_18055_, _17949_, _03178_);
  or (_18056_, _18055_, _18054_);
  and (_18057_, _18056_, _34698_);
  and (_18058_, _18057_, _18053_);
  or (_35216_, _18058_, _17948_);
  nor (_18059_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_18061_, _18059_, _04548_);
  and (_18062_, _08539_, \oc8051_golden_model_1.P1 [4]);
  and (_18063_, _11368_, _04719_);
  or (_18064_, _18063_, _18062_);
  and (_18065_, _18064_, _03130_);
  nor (_18066_, _05202_, _08539_);
  or (_18067_, _18066_, _18062_);
  or (_18068_, _18067_, _06241_);
  and (_18069_, _17969_, \oc8051_golden_model_1.P1 [4]);
  and (_18070_, _11243_, _05344_);
  or (_18072_, _18070_, _18069_);
  and (_18073_, _18072_, _02887_);
  nor (_18074_, _11259_, _08539_);
  or (_18075_, _18074_, _18062_);
  or (_18076_, _18075_, _03821_);
  and (_18077_, _04719_, \oc8051_golden_model_1.ACC [4]);
  or (_18078_, _18077_, _18062_);
  and (_18079_, _18078_, _03825_);
  and (_18080_, _03826_, \oc8051_golden_model_1.P1 [4]);
  or (_18081_, _18080_, _02952_);
  or (_18083_, _18081_, _18079_);
  and (_18084_, _18083_, _02892_);
  and (_18085_, _18084_, _18076_);
  and (_18086_, _11245_, _05344_);
  or (_18087_, _18086_, _18069_);
  and (_18088_, _18087_, _02891_);
  or (_18089_, _18088_, _02947_);
  or (_18090_, _18089_, _18085_);
  or (_18091_, _18067_, _03327_);
  and (_18092_, _18091_, _18090_);
  or (_18094_, _18092_, _02950_);
  or (_18095_, _18078_, _02959_);
  and (_18096_, _18095_, _02888_);
  and (_18097_, _18096_, _18094_);
  or (_18098_, _18097_, _18073_);
  and (_18099_, _18098_, _02881_);
  and (_18100_, _11277_, _05344_);
  or (_18101_, _18100_, _18069_);
  and (_18102_, _18101_, _02880_);
  or (_18103_, _18102_, _18099_);
  and (_18105_, _18103_, _02875_);
  and (_18106_, _17285_, _05344_);
  or (_18107_, _18106_, _18069_);
  and (_18108_, _18107_, _02874_);
  or (_18109_, _18108_, _06793_);
  or (_18110_, _18109_, _18105_);
  and (_18111_, _18110_, _18068_);
  or (_18112_, _18111_, _02855_);
  and (_18113_, _06181_, _04719_);
  or (_18114_, _18062_, _02856_);
  or (_18116_, _18114_, _18113_);
  and (_18117_, _18116_, _02851_);
  and (_18118_, _18117_, _18112_);
  and (_18119_, _17311_, _04719_);
  or (_18120_, _18119_, _18062_);
  and (_18121_, _18120_, _02576_);
  or (_18122_, _18121_, _03014_);
  or (_18123_, _18122_, _18118_);
  and (_18124_, _05697_, _04719_);
  or (_18125_, _18124_, _18062_);
  or (_18127_, _18125_, _03884_);
  and (_18128_, _18127_, _18123_);
  or (_18129_, _18128_, _03021_);
  and (_18130_, _11362_, _04719_);
  or (_18131_, _18062_, _05279_);
  or (_18132_, _18131_, _18130_);
  and (_18133_, _18132_, _03131_);
  and (_18134_, _18133_, _18129_);
  or (_18135_, _18134_, _18065_);
  and (_18136_, _18135_, _05274_);
  or (_18138_, _18062_, _05251_);
  and (_18139_, _18125_, _03020_);
  and (_18140_, _18139_, _18138_);
  or (_18141_, _18140_, _18136_);
  and (_18142_, _18141_, _03140_);
  and (_18143_, _18078_, _03139_);
  and (_18144_, _18143_, _18138_);
  or (_18145_, _18144_, _03036_);
  or (_18146_, _18145_, _18142_);
  nor (_18147_, _11361_, _08539_);
  or (_18149_, _18062_, _05781_);
  or (_18150_, _18149_, _18147_);
  and (_18151_, _18150_, _05786_);
  and (_18152_, _18151_, _18146_);
  nor (_18153_, _11367_, _08539_);
  or (_18154_, _18153_, _18062_);
  and (_18155_, _18154_, _03127_);
  or (_18156_, _18155_, _03166_);
  or (_18157_, _18156_, _18152_);
  or (_18158_, _18075_, _03563_);
  and (_18160_, _18158_, _02501_);
  and (_18161_, _18160_, _18157_);
  and (_18162_, _18072_, _02500_);
  or (_18163_, _18162_, _03174_);
  or (_18164_, _18163_, _18161_);
  and (_18165_, _11417_, _04719_);
  or (_18166_, _18062_, _03178_);
  or (_18167_, _18166_, _18165_);
  and (_18168_, _18167_, _34698_);
  and (_18169_, _18168_, _18164_);
  or (_35217_, _18169_, _18061_);
  nor (_18171_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_18172_, _18171_, _04548_);
  and (_18173_, _08539_, \oc8051_golden_model_1.P1 [5]);
  and (_18174_, _11436_, _04719_);
  or (_18175_, _18174_, _18173_);
  and (_18176_, _18175_, _03130_);
  nor (_18177_, _11445_, _08539_);
  or (_18178_, _18177_, _18173_);
  or (_18179_, _18178_, _03821_);
  and (_18181_, _04719_, \oc8051_golden_model_1.ACC [5]);
  or (_18182_, _18181_, _18173_);
  and (_18183_, _18182_, _03825_);
  and (_18184_, _03826_, \oc8051_golden_model_1.P1 [5]);
  or (_18185_, _18184_, _02952_);
  or (_18186_, _18185_, _18183_);
  and (_18187_, _18186_, _02892_);
  and (_18188_, _18187_, _18179_);
  and (_18189_, _17969_, \oc8051_golden_model_1.P1 [5]);
  and (_18190_, _11459_, _05344_);
  or (_18192_, _18190_, _18189_);
  and (_18193_, _18192_, _02891_);
  or (_18194_, _18193_, _02947_);
  or (_18195_, _18194_, _18188_);
  nor (_18196_, _04896_, _08539_);
  or (_18197_, _18196_, _18173_);
  or (_18198_, _18197_, _03327_);
  and (_18199_, _18198_, _18195_);
  or (_18200_, _18199_, _02950_);
  or (_18201_, _18182_, _02959_);
  and (_18203_, _18201_, _02888_);
  and (_18204_, _18203_, _18200_);
  and (_18205_, _11442_, _05344_);
  or (_18206_, _18205_, _18189_);
  and (_18207_, _18206_, _02887_);
  or (_18208_, _18207_, _02880_);
  or (_18209_, _18208_, _18204_);
  or (_18210_, _18189_, _11474_);
  and (_18211_, _18210_, _18192_);
  or (_18212_, _18211_, _02881_);
  and (_18214_, _18212_, _02875_);
  and (_18215_, _18214_, _18209_);
  and (_18216_, _17409_, _05344_);
  or (_18217_, _18216_, _18189_);
  and (_18218_, _18217_, _02874_);
  or (_18219_, _18218_, _06793_);
  or (_18220_, _18219_, _18215_);
  or (_18221_, _18197_, _06241_);
  and (_18222_, _18221_, _18220_);
  or (_18223_, _18222_, _02855_);
  and (_18225_, _06180_, _04719_);
  or (_18226_, _18173_, _02856_);
  or (_18227_, _18226_, _18225_);
  and (_18228_, _18227_, _02851_);
  and (_18229_, _18228_, _18223_);
  and (_18230_, _17436_, _04719_);
  or (_18231_, _18230_, _18173_);
  and (_18232_, _18231_, _02576_);
  or (_18233_, _18232_, _03014_);
  or (_18234_, _18233_, _18229_);
  and (_18236_, _05701_, _04719_);
  or (_18237_, _18236_, _18173_);
  or (_18238_, _18237_, _03884_);
  and (_18239_, _18238_, _18234_);
  or (_18240_, _18239_, _03021_);
  and (_18241_, _11562_, _04719_);
  or (_18242_, _18173_, _05279_);
  or (_18243_, _18242_, _18241_);
  and (_18244_, _18243_, _03131_);
  and (_18245_, _18244_, _18240_);
  or (_18247_, _18245_, _18176_);
  and (_18248_, _18247_, _05274_);
  or (_18249_, _18173_, _04944_);
  and (_18250_, _18237_, _03020_);
  and (_18251_, _18250_, _18249_);
  or (_18252_, _18251_, _18248_);
  and (_18253_, _18252_, _03140_);
  and (_18254_, _18182_, _03139_);
  and (_18255_, _18254_, _18249_);
  or (_18256_, _18255_, _03036_);
  or (_18258_, _18256_, _18253_);
  nor (_18259_, _11560_, _08539_);
  or (_18260_, _18173_, _05781_);
  or (_18261_, _18260_, _18259_);
  and (_18262_, _18261_, _05786_);
  and (_18263_, _18262_, _18258_);
  nor (_18264_, _11435_, _08539_);
  or (_18265_, _18264_, _18173_);
  and (_18266_, _18265_, _03127_);
  or (_18267_, _18266_, _03166_);
  or (_18269_, _18267_, _18263_);
  or (_18270_, _18178_, _03563_);
  and (_18271_, _18270_, _02501_);
  and (_18272_, _18271_, _18269_);
  and (_18273_, _18206_, _02500_);
  or (_18274_, _18273_, _03174_);
  or (_18275_, _18274_, _18272_);
  and (_18276_, _11619_, _04719_);
  or (_18277_, _18173_, _03178_);
  or (_18278_, _18277_, _18276_);
  and (_18280_, _18278_, _34698_);
  and (_18281_, _18280_, _18275_);
  or (_35218_, _18281_, _18172_);
  not (_18282_, \oc8051_golden_model_1.P1 [6]);
  nor (_18283_, _34698_, _18282_);
  or (_18284_, _18283_, rst);
  nor (_18285_, _04719_, _18282_);
  and (_18286_, _11769_, _04719_);
  or (_18287_, _18286_, _18285_);
  and (_18288_, _18287_, _03130_);
  nor (_18290_, _11636_, _08539_);
  or (_18291_, _18290_, _18285_);
  or (_18292_, _18291_, _03821_);
  and (_18293_, _04719_, \oc8051_golden_model_1.ACC [6]);
  or (_18294_, _18293_, _18285_);
  and (_18295_, _18294_, _03825_);
  nor (_18296_, _03825_, _18282_);
  or (_18297_, _18296_, _02952_);
  or (_18298_, _18297_, _18295_);
  and (_18299_, _18298_, _02892_);
  and (_18301_, _18299_, _18292_);
  nor (_18302_, _05344_, _18282_);
  and (_18303_, _11653_, _05344_);
  or (_18304_, _18303_, _18302_);
  and (_18305_, _18304_, _02891_);
  or (_18306_, _18305_, _02947_);
  or (_18307_, _18306_, _18301_);
  nor (_18308_, _04787_, _08539_);
  or (_18309_, _18308_, _18285_);
  or (_18310_, _18309_, _03327_);
  and (_18312_, _18310_, _18307_);
  or (_18313_, _18312_, _02950_);
  or (_18314_, _18294_, _02959_);
  and (_18315_, _18314_, _02888_);
  and (_18316_, _18315_, _18313_);
  and (_18317_, _11675_, _05344_);
  or (_18318_, _18317_, _18302_);
  and (_18319_, _18318_, _02887_);
  or (_18320_, _18319_, _02880_);
  or (_18321_, _18320_, _18316_);
  or (_18323_, _18302_, _11682_);
  and (_18324_, _18323_, _18304_);
  or (_18325_, _18324_, _02881_);
  and (_18326_, _18325_, _02875_);
  and (_18327_, _18326_, _18321_);
  and (_18328_, _17535_, _05344_);
  or (_18329_, _18328_, _18302_);
  and (_18330_, _18329_, _02874_);
  or (_18331_, _18330_, _06793_);
  or (_18332_, _18331_, _18327_);
  or (_18334_, _18309_, _06241_);
  and (_18335_, _18334_, _18332_);
  or (_18336_, _18335_, _02855_);
  and (_18337_, _05847_, _04719_);
  or (_18338_, _18285_, _02856_);
  or (_18339_, _18338_, _18337_);
  and (_18340_, _18339_, _02851_);
  and (_18341_, _18340_, _18336_);
  and (_18342_, _17563_, _04719_);
  or (_18343_, _18342_, _18285_);
  and (_18345_, _18343_, _02576_);
  or (_18346_, _18345_, _03014_);
  or (_18347_, _18346_, _18341_);
  and (_18348_, _11758_, _04719_);
  or (_18349_, _18348_, _18285_);
  or (_18350_, _18349_, _03884_);
  and (_18351_, _18350_, _18347_);
  or (_18352_, _18351_, _03021_);
  and (_18353_, _11646_, _04719_);
  or (_18354_, _18285_, _05279_);
  or (_18356_, _18354_, _18353_);
  and (_18357_, _18356_, _03131_);
  and (_18358_, _18357_, _18352_);
  or (_18359_, _18358_, _18288_);
  and (_18360_, _18359_, _05274_);
  or (_18361_, _18285_, _04838_);
  and (_18362_, _18349_, _03020_);
  and (_18363_, _18362_, _18361_);
  or (_18364_, _18363_, _18360_);
  and (_18365_, _18364_, _03140_);
  and (_18367_, _18294_, _03139_);
  and (_18368_, _18367_, _18361_);
  or (_18369_, _18368_, _03036_);
  or (_18370_, _18369_, _18365_);
  nor (_18371_, _11644_, _08539_);
  or (_18372_, _18285_, _05781_);
  or (_18373_, _18372_, _18371_);
  and (_18374_, _18373_, _05786_);
  and (_18375_, _18374_, _18370_);
  nor (_18376_, _11768_, _08539_);
  or (_18378_, _18376_, _18285_);
  and (_18379_, _18378_, _03127_);
  or (_18380_, _18379_, _03166_);
  or (_18381_, _18380_, _18375_);
  or (_18382_, _18291_, _03563_);
  and (_18383_, _18382_, _02501_);
  and (_18384_, _18383_, _18381_);
  and (_18385_, _18318_, _02500_);
  or (_18386_, _18385_, _03174_);
  or (_18387_, _18386_, _18384_);
  and (_18389_, _11821_, _04719_);
  or (_18390_, _18285_, _03178_);
  or (_18391_, _18390_, _18389_);
  and (_18392_, _18391_, _34698_);
  and (_18393_, _18392_, _18387_);
  or (_35219_, _18393_, _18284_);
  not (_18394_, \oc8051_golden_model_1.P2 [0]);
  nor (_18395_, _34698_, _18394_);
  or (_18396_, _18395_, rst);
  nor (_18397_, _04722_, _18394_);
  and (_18399_, _10546_, _04722_);
  or (_18400_, _18399_, _18397_);
  and (_18401_, _18400_, _03130_);
  and (_18402_, _04722_, _03817_);
  or (_18403_, _18402_, _18397_);
  or (_18404_, _18403_, _06241_);
  and (_18405_, _05044_, _04722_);
  or (_18406_, _18405_, _18397_);
  and (_18407_, _18406_, _02952_);
  nor (_18408_, _03825_, _18394_);
  and (_18410_, _04722_, \oc8051_golden_model_1.ACC [0]);
  or (_18411_, _18410_, _18397_);
  and (_18412_, _18411_, _03825_);
  or (_18413_, _18412_, _18408_);
  and (_18414_, _18413_, _03821_);
  or (_18415_, _18414_, _02891_);
  or (_18416_, _18415_, _18407_);
  and (_18417_, _10429_, _05346_);
  nor (_18418_, _05346_, _18394_);
  or (_18419_, _18418_, _02892_);
  or (_18421_, _18419_, _18417_);
  and (_18422_, _18421_, _03327_);
  and (_18423_, _18422_, _18416_);
  and (_18424_, _18403_, _02947_);
  or (_18425_, _18424_, _02950_);
  or (_18426_, _18425_, _18423_);
  or (_18427_, _18411_, _02959_);
  and (_18428_, _18427_, _02888_);
  and (_18429_, _18428_, _18426_);
  and (_18430_, _18397_, _02887_);
  or (_18432_, _18430_, _02880_);
  or (_18433_, _18432_, _18429_);
  or (_18434_, _18406_, _02881_);
  and (_18435_, _18434_, _02875_);
  and (_18436_, _18435_, _18433_);
  and (_18437_, _16789_, _05346_);
  or (_18438_, _18437_, _18418_);
  and (_18439_, _18438_, _02874_);
  or (_18440_, _18439_, _06793_);
  or (_18441_, _18440_, _18436_);
  and (_18443_, _18441_, _18404_);
  or (_18444_, _18443_, _02855_);
  and (_18445_, _06174_, _04722_);
  or (_18446_, _18397_, _02856_);
  or (_18447_, _18446_, _18445_);
  and (_18448_, _18447_, _02851_);
  and (_18449_, _18448_, _18444_);
  and (_18450_, _16814_, _04722_);
  or (_18451_, _18450_, _18397_);
  and (_18452_, _18451_, _02576_);
  or (_18454_, _18452_, _03014_);
  or (_18455_, _18454_, _18449_);
  and (_18456_, _04722_, _05566_);
  or (_18457_, _18456_, _18397_);
  or (_18458_, _18457_, _03884_);
  and (_18459_, _18458_, _18455_);
  or (_18460_, _18459_, _03021_);
  and (_18461_, _10425_, _04722_);
  or (_18462_, _18397_, _05279_);
  or (_18463_, _18462_, _18461_);
  and (_18465_, _18463_, _03131_);
  and (_18466_, _18465_, _18460_);
  or (_18467_, _18466_, _18401_);
  and (_18468_, _18467_, _05274_);
  nand (_18469_, _18457_, _03020_);
  nor (_18470_, _18469_, _18405_);
  or (_18471_, _18470_, _18468_);
  and (_18472_, _18471_, _03140_);
  or (_18473_, _18397_, _09183_);
  and (_18474_, _18411_, _03139_);
  and (_18476_, _18474_, _18473_);
  or (_18477_, _18476_, _03036_);
  or (_18478_, _18477_, _18472_);
  nor (_18479_, _10423_, _08642_);
  or (_18480_, _18397_, _05781_);
  or (_18481_, _18480_, _18479_);
  and (_18482_, _18481_, _05786_);
  and (_18483_, _18482_, _18478_);
  nor (_18484_, _10421_, _08642_);
  or (_18485_, _18484_, _18397_);
  and (_18487_, _18485_, _03127_);
  or (_18488_, _18487_, _03166_);
  or (_18489_, _18488_, _18483_);
  or (_18490_, _18406_, _03563_);
  and (_18491_, _18490_, _02501_);
  and (_18492_, _18491_, _18489_);
  and (_18493_, _18397_, _02500_);
  or (_18494_, _18493_, _03174_);
  or (_18495_, _18494_, _18492_);
  or (_18496_, _18406_, _03178_);
  and (_18498_, _18496_, _34698_);
  and (_18499_, _18498_, _18495_);
  or (_35221_, _18499_, _18396_);
  not (_18500_, \oc8051_golden_model_1.P2 [1]);
  nor (_18501_, _34698_, _18500_);
  or (_18502_, _18501_, rst);
  nand (_18503_, _04722_, _03705_);
  or (_18504_, _04722_, \oc8051_golden_model_1.P2 [1]);
  and (_18505_, _18504_, _03014_);
  and (_18506_, _18505_, _18503_);
  and (_18508_, _10622_, _04722_);
  not (_18509_, _18508_);
  and (_18510_, _18509_, _18504_);
  or (_18511_, _18510_, _03821_);
  nand (_18512_, _04722_, _02618_);
  and (_18513_, _18512_, _18504_);
  and (_18514_, _18513_, _03825_);
  nor (_18515_, _03825_, _18500_);
  or (_18516_, _18515_, _02952_);
  or (_18517_, _18516_, _18514_);
  and (_18519_, _18517_, _02892_);
  and (_18520_, _18519_, _18511_);
  and (_18521_, _10617_, _05346_);
  nor (_18522_, _05346_, _18500_);
  or (_18523_, _18522_, _02947_);
  or (_18524_, _18523_, _18521_);
  and (_18525_, _18524_, _09918_);
  or (_18526_, _18525_, _18520_);
  nor (_18527_, _04722_, _18500_);
  and (_18528_, _04722_, _04005_);
  or (_18530_, _18528_, _18527_);
  or (_18531_, _18530_, _03327_);
  and (_18532_, _18531_, _18526_);
  or (_18533_, _18532_, _02950_);
  or (_18534_, _18513_, _02959_);
  and (_18535_, _18534_, _02888_);
  and (_18536_, _18535_, _18533_);
  and (_18537_, _10620_, _05346_);
  or (_18538_, _18537_, _18522_);
  and (_18539_, _18538_, _02887_);
  or (_18541_, _18539_, _02880_);
  or (_18542_, _18541_, _18536_);
  and (_18543_, _18521_, _10616_);
  or (_18544_, _18522_, _02881_);
  or (_18545_, _18544_, _18543_);
  and (_18546_, _18545_, _18542_);
  and (_18547_, _18546_, _02875_);
  and (_18548_, _16909_, _05346_);
  or (_18549_, _18522_, _18548_);
  and (_18550_, _18549_, _02874_);
  or (_18552_, _18550_, _06793_);
  or (_18553_, _18552_, _18547_);
  or (_18554_, _18530_, _06241_);
  and (_18555_, _18554_, _18553_);
  or (_18556_, _18555_, _02855_);
  and (_18557_, _06173_, _04722_);
  or (_18558_, _18527_, _02856_);
  or (_18559_, _18558_, _18557_);
  and (_18560_, _18559_, _02851_);
  and (_18561_, _18560_, _18556_);
  and (_18563_, _16935_, _04722_);
  or (_18564_, _18563_, _18527_);
  and (_18565_, _18564_, _02576_);
  or (_18566_, _18565_, _18561_);
  and (_18567_, _18566_, _03884_);
  or (_18568_, _18567_, _18506_);
  and (_18569_, _18568_, _05279_);
  or (_18570_, _10612_, _08642_);
  and (_18571_, _18504_, _03021_);
  and (_18572_, _18571_, _18570_);
  or (_18574_, _18572_, _18569_);
  and (_18575_, _18574_, _03131_);
  or (_18576_, _10739_, _08642_);
  and (_18577_, _18504_, _03130_);
  and (_18578_, _18577_, _18576_);
  or (_18579_, _18578_, _18575_);
  and (_18580_, _18579_, _05274_);
  or (_18581_, _10611_, _08642_);
  and (_18582_, _18504_, _03020_);
  and (_18583_, _18582_, _18581_);
  or (_18585_, _18583_, _18580_);
  and (_18586_, _18585_, _03140_);
  or (_18587_, _18527_, _12724_);
  and (_18588_, _18513_, _03139_);
  and (_18589_, _18588_, _18587_);
  or (_18590_, _18589_, _18586_);
  and (_18591_, _18590_, _03128_);
  or (_18592_, _18503_, _12724_);
  and (_18593_, _18504_, _03036_);
  and (_18594_, _18593_, _18592_);
  or (_18596_, _18512_, _12724_);
  and (_18597_, _18504_, _03127_);
  and (_18598_, _18597_, _18596_);
  or (_18599_, _18598_, _03166_);
  or (_18600_, _18599_, _18594_);
  or (_18601_, _18600_, _18591_);
  or (_18602_, _18510_, _03563_);
  and (_18603_, _18602_, _02501_);
  and (_18604_, _18603_, _18601_);
  and (_18605_, _18538_, _02500_);
  or (_18607_, _18605_, _03174_);
  or (_18608_, _18607_, _18604_);
  or (_18609_, _18527_, _03178_);
  or (_18610_, _18609_, _18508_);
  and (_18611_, _18610_, _34698_);
  and (_18612_, _18611_, _18608_);
  or (_35222_, _18612_, _18502_);
  not (_18613_, \oc8051_golden_model_1.P2 [2]);
  nor (_18614_, _34698_, _18613_);
  or (_18615_, _18614_, rst);
  nor (_18617_, _04722_, _18613_);
  and (_18618_, _10831_, _04722_);
  or (_18619_, _18618_, _18617_);
  and (_18620_, _18619_, _03130_);
  nor (_18621_, _08642_, _04440_);
  or (_18622_, _18621_, _18617_);
  or (_18623_, _18622_, _06241_);
  or (_18624_, _18622_, _03327_);
  nor (_18625_, _10849_, _08642_);
  or (_18626_, _18625_, _18617_);
  or (_18628_, _18626_, _03821_);
  and (_18629_, _04722_, \oc8051_golden_model_1.ACC [2]);
  or (_18630_, _18629_, _18617_);
  and (_18631_, _18630_, _03825_);
  nor (_18632_, _03825_, _18613_);
  or (_18633_, _18632_, _02952_);
  or (_18634_, _18633_, _18631_);
  and (_18635_, _18634_, _02892_);
  and (_18636_, _18635_, _18628_);
  nor (_18637_, _05346_, _18613_);
  and (_18639_, _10853_, _05346_);
  or (_18640_, _18639_, _18637_);
  and (_18641_, _18640_, _02891_);
  or (_18642_, _18641_, _02947_);
  or (_18643_, _18642_, _18636_);
  and (_18644_, _18643_, _18624_);
  or (_18645_, _18644_, _02950_);
  or (_18646_, _18630_, _02959_);
  and (_18647_, _18646_, _02888_);
  and (_18648_, _18647_, _18645_);
  and (_18650_, _10838_, _05346_);
  or (_18651_, _18650_, _18637_);
  and (_18652_, _18651_, _02887_);
  or (_18653_, _18652_, _02880_);
  or (_18654_, _18653_, _18648_);
  and (_18655_, _18639_, _10868_);
  or (_18656_, _18637_, _02881_);
  or (_18657_, _18656_, _18655_);
  and (_18658_, _18657_, _02875_);
  and (_18659_, _18658_, _18654_);
  and (_18661_, _17034_, _05346_);
  or (_18662_, _18661_, _18637_);
  and (_18663_, _18662_, _02874_);
  or (_18664_, _18663_, _06793_);
  or (_18665_, _18664_, _18659_);
  and (_18666_, _18665_, _18623_);
  or (_18667_, _18666_, _02855_);
  and (_18668_, _06177_, _04722_);
  or (_18669_, _18617_, _02856_);
  or (_18670_, _18669_, _18668_);
  and (_18672_, _18670_, _02851_);
  and (_18673_, _18672_, _18667_);
  and (_18674_, _17060_, _04722_);
  or (_18675_, _18674_, _18617_);
  and (_18676_, _18675_, _02576_);
  or (_18677_, _18676_, _03014_);
  or (_18678_, _18677_, _18673_);
  and (_18679_, _04722_, _05727_);
  or (_18680_, _18679_, _18617_);
  or (_18681_, _18680_, _03884_);
  and (_18683_, _18681_, _18678_);
  or (_18684_, _18683_, _03021_);
  and (_18685_, _10835_, _04722_);
  or (_18686_, _18617_, _05279_);
  or (_18687_, _18686_, _18685_);
  and (_18688_, _18687_, _03131_);
  and (_18689_, _18688_, _18684_);
  or (_18690_, _18689_, _18620_);
  and (_18691_, _18690_, _05274_);
  or (_18692_, _18617_, _05143_);
  and (_18694_, _18680_, _03020_);
  and (_18695_, _18694_, _18692_);
  or (_18696_, _18695_, _18691_);
  and (_18697_, _18696_, _03140_);
  and (_18698_, _18630_, _03139_);
  and (_18699_, _18698_, _18692_);
  or (_18700_, _18699_, _03036_);
  or (_18701_, _18700_, _18697_);
  nor (_18702_, _10833_, _08642_);
  or (_18703_, _18617_, _05781_);
  or (_18705_, _18703_, _18702_);
  and (_18706_, _18705_, _05786_);
  and (_18707_, _18706_, _18701_);
  nor (_18708_, _10830_, _08642_);
  or (_18709_, _18708_, _18617_);
  and (_18710_, _18709_, _03127_);
  or (_18711_, _18710_, _03166_);
  or (_18712_, _18711_, _18707_);
  or (_18713_, _18626_, _03563_);
  and (_18714_, _18713_, _02501_);
  and (_18716_, _18714_, _18712_);
  and (_18717_, _18651_, _02500_);
  or (_18718_, _18717_, _03174_);
  or (_18719_, _18718_, _18716_);
  and (_18720_, _11008_, _04722_);
  or (_18721_, _18617_, _03178_);
  or (_18722_, _18721_, _18720_);
  and (_18723_, _18722_, _34698_);
  and (_18724_, _18723_, _18719_);
  or (_35223_, _18724_, _18615_);
  nor (_18726_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_18727_, _18726_, _04548_);
  and (_18728_, _08642_, \oc8051_golden_model_1.P2 [3]);
  and (_18729_, _11028_, _04722_);
  or (_18730_, _18729_, _18728_);
  and (_18731_, _18730_, _03130_);
  nor (_18732_, _08642_, _04242_);
  or (_18733_, _18732_, _18728_);
  or (_18734_, _18733_, _06241_);
  nor (_18735_, _11040_, _08642_);
  or (_18737_, _18735_, _18728_);
  or (_18738_, _18737_, _03821_);
  and (_18739_, _04722_, \oc8051_golden_model_1.ACC [3]);
  or (_18740_, _18739_, _18728_);
  and (_18741_, _18740_, _03825_);
  and (_18742_, _03826_, \oc8051_golden_model_1.P2 [3]);
  or (_18743_, _18742_, _02952_);
  or (_18744_, _18743_, _18741_);
  and (_18745_, _18744_, _02892_);
  and (_18746_, _18745_, _18738_);
  not (_18748_, _05346_);
  and (_18749_, _18748_, \oc8051_golden_model_1.P2 [3]);
  and (_18750_, _11037_, _05346_);
  or (_18751_, _18750_, _18749_);
  and (_18752_, _18751_, _02891_);
  or (_18753_, _18752_, _02947_);
  or (_18754_, _18753_, _18746_);
  or (_18755_, _18733_, _03327_);
  and (_18756_, _18755_, _18754_);
  or (_18757_, _18756_, _02950_);
  or (_18759_, _18740_, _02959_);
  and (_18760_, _18759_, _02888_);
  and (_18761_, _18760_, _18757_);
  and (_18762_, _11035_, _05346_);
  or (_18763_, _18762_, _18749_);
  and (_18764_, _18763_, _02887_);
  or (_18765_, _18764_, _02880_);
  or (_18766_, _18765_, _18761_);
  or (_18767_, _18749_, _11066_);
  and (_18768_, _18767_, _18751_);
  or (_18770_, _18768_, _02881_);
  and (_18771_, _18770_, _02875_);
  and (_18772_, _18771_, _18766_);
  and (_18773_, _17160_, _05346_);
  or (_18774_, _18773_, _18749_);
  and (_18775_, _18774_, _02874_);
  or (_18776_, _18775_, _06793_);
  or (_18777_, _18776_, _18772_);
  and (_18778_, _18777_, _18734_);
  or (_18779_, _18778_, _02855_);
  and (_18781_, _06176_, _04722_);
  or (_18782_, _18728_, _02856_);
  or (_18783_, _18782_, _18781_);
  and (_18784_, _18783_, _02851_);
  and (_18785_, _18784_, _18779_);
  and (_18786_, _17185_, _04722_);
  or (_18787_, _18786_, _18728_);
  and (_18788_, _18787_, _02576_);
  or (_18789_, _18788_, _03014_);
  or (_18790_, _18789_, _18785_);
  and (_18792_, _04722_, _05664_);
  or (_18793_, _18792_, _18728_);
  or (_18794_, _18793_, _03884_);
  and (_18795_, _18794_, _18790_);
  or (_18796_, _18795_, _03021_);
  and (_18797_, _11032_, _04722_);
  or (_18798_, _18728_, _05279_);
  or (_18799_, _18798_, _18797_);
  and (_18800_, _18799_, _03131_);
  and (_18801_, _18800_, _18796_);
  or (_18803_, _18801_, _18731_);
  and (_18804_, _18803_, _05274_);
  or (_18805_, _18728_, _04996_);
  and (_18806_, _18793_, _03020_);
  and (_18807_, _18806_, _18805_);
  or (_18808_, _18807_, _18804_);
  and (_18809_, _18808_, _03140_);
  and (_18810_, _18740_, _03139_);
  and (_18811_, _18810_, _18805_);
  or (_18812_, _18811_, _03036_);
  or (_18814_, _18812_, _18809_);
  nor (_18815_, _11030_, _08642_);
  or (_18816_, _18728_, _05781_);
  or (_18817_, _18816_, _18815_);
  and (_18818_, _18817_, _05786_);
  and (_18819_, _18818_, _18814_);
  nor (_18820_, _11027_, _08642_);
  or (_18821_, _18820_, _18728_);
  and (_18822_, _18821_, _03127_);
  or (_18823_, _18822_, _03166_);
  or (_18825_, _18823_, _18819_);
  or (_18826_, _18737_, _03563_);
  and (_18827_, _18826_, _02501_);
  and (_18828_, _18827_, _18825_);
  and (_18829_, _18763_, _02500_);
  or (_18830_, _18829_, _03174_);
  or (_18831_, _18830_, _18828_);
  and (_18832_, _11213_, _04722_);
  or (_18833_, _18728_, _03178_);
  or (_18834_, _18833_, _18832_);
  and (_18836_, _18834_, _34698_);
  and (_18837_, _18836_, _18831_);
  or (_35224_, _18837_, _18727_);
  nor (_18838_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_18839_, _18838_, _04548_);
  and (_18840_, _08642_, \oc8051_golden_model_1.P2 [4]);
  and (_18841_, _11368_, _04722_);
  or (_18842_, _18841_, _18840_);
  and (_18843_, _18842_, _03130_);
  nor (_18844_, _05202_, _08642_);
  or (_18846_, _18844_, _18840_);
  or (_18847_, _18846_, _06241_);
  and (_18848_, _18748_, \oc8051_golden_model_1.P2 [4]);
  and (_18849_, _11243_, _05346_);
  or (_18850_, _18849_, _18848_);
  and (_18851_, _18850_, _02887_);
  nor (_18852_, _11259_, _08642_);
  or (_18853_, _18852_, _18840_);
  or (_18854_, _18853_, _03821_);
  and (_18855_, _04722_, \oc8051_golden_model_1.ACC [4]);
  or (_18857_, _18855_, _18840_);
  and (_18858_, _18857_, _03825_);
  and (_18859_, _03826_, \oc8051_golden_model_1.P2 [4]);
  or (_18860_, _18859_, _02952_);
  or (_18861_, _18860_, _18858_);
  and (_18862_, _18861_, _02892_);
  and (_18863_, _18862_, _18854_);
  and (_18864_, _11245_, _05346_);
  or (_18865_, _18864_, _18848_);
  and (_18866_, _18865_, _02891_);
  or (_18868_, _18866_, _02947_);
  or (_18869_, _18868_, _18863_);
  or (_18870_, _18846_, _03327_);
  and (_18871_, _18870_, _18869_);
  or (_18872_, _18871_, _02950_);
  or (_18873_, _18857_, _02959_);
  and (_18874_, _18873_, _02888_);
  and (_18875_, _18874_, _18872_);
  or (_18876_, _18875_, _18851_);
  and (_18877_, _18876_, _02881_);
  or (_18879_, _18848_, _11276_);
  and (_18880_, _18879_, _02880_);
  and (_18881_, _18880_, _18865_);
  or (_18882_, _18881_, _18877_);
  and (_18883_, _18882_, _02875_);
  and (_18884_, _17285_, _05346_);
  or (_18885_, _18884_, _18848_);
  and (_18886_, _18885_, _02874_);
  or (_18887_, _18886_, _06793_);
  or (_18888_, _18887_, _18883_);
  and (_18890_, _18888_, _18847_);
  or (_18891_, _18890_, _02855_);
  and (_18892_, _06181_, _04722_);
  or (_18893_, _18840_, _02856_);
  or (_18894_, _18893_, _18892_);
  and (_18895_, _18894_, _02851_);
  and (_18896_, _18895_, _18891_);
  and (_18897_, _17311_, _04722_);
  or (_18898_, _18897_, _18840_);
  and (_18899_, _18898_, _02576_);
  or (_18901_, _18899_, _03014_);
  or (_18902_, _18901_, _18896_);
  and (_18903_, _05697_, _04722_);
  or (_18904_, _18903_, _18840_);
  or (_18905_, _18904_, _03884_);
  and (_18906_, _18905_, _18902_);
  or (_18907_, _18906_, _03021_);
  and (_18908_, _11362_, _04722_);
  or (_18909_, _18840_, _05279_);
  or (_18910_, _18909_, _18908_);
  and (_18912_, _18910_, _03131_);
  and (_18913_, _18912_, _18907_);
  or (_18914_, _18913_, _18843_);
  and (_18915_, _18914_, _05274_);
  or (_18916_, _18840_, _05251_);
  and (_18917_, _18904_, _03020_);
  and (_18918_, _18917_, _18916_);
  or (_18919_, _18918_, _18915_);
  and (_18920_, _18919_, _03140_);
  and (_18921_, _18857_, _03139_);
  and (_18923_, _18921_, _18916_);
  or (_18924_, _18923_, _03036_);
  or (_18925_, _18924_, _18920_);
  nor (_18926_, _11361_, _08642_);
  or (_18927_, _18840_, _05781_);
  or (_18928_, _18927_, _18926_);
  and (_18929_, _18928_, _05786_);
  and (_18930_, _18929_, _18925_);
  nor (_18931_, _11367_, _08642_);
  or (_18932_, _18931_, _18840_);
  and (_18934_, _18932_, _03127_);
  or (_18935_, _18934_, _03166_);
  or (_18936_, _18935_, _18930_);
  or (_18937_, _18853_, _03563_);
  and (_18938_, _18937_, _02501_);
  and (_18939_, _18938_, _18936_);
  and (_18940_, _18850_, _02500_);
  or (_18941_, _18940_, _03174_);
  or (_18942_, _18941_, _18939_);
  and (_18943_, _11417_, _04722_);
  or (_18945_, _18840_, _03178_);
  or (_18946_, _18945_, _18943_);
  and (_18947_, _18946_, _34698_);
  and (_18948_, _18947_, _18942_);
  or (_35225_, _18948_, _18839_);
  nor (_18949_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_18950_, _18949_, _04548_);
  and (_18951_, _08642_, \oc8051_golden_model_1.P2 [5]);
  and (_18952_, _11436_, _04722_);
  or (_18953_, _18952_, _18951_);
  and (_18955_, _18953_, _03130_);
  nor (_18956_, _11445_, _08642_);
  or (_18957_, _18956_, _18951_);
  or (_18958_, _18957_, _03821_);
  and (_18959_, _04722_, \oc8051_golden_model_1.ACC [5]);
  or (_18960_, _18959_, _18951_);
  and (_18961_, _18960_, _03825_);
  and (_18962_, _03826_, \oc8051_golden_model_1.P2 [5]);
  or (_18963_, _18962_, _02952_);
  or (_18964_, _18963_, _18961_);
  and (_18966_, _18964_, _02892_);
  and (_18967_, _18966_, _18958_);
  and (_18968_, _18748_, \oc8051_golden_model_1.P2 [5]);
  and (_18969_, _11459_, _05346_);
  or (_18970_, _18969_, _18968_);
  and (_18971_, _18970_, _02891_);
  or (_18972_, _18971_, _02947_);
  or (_18973_, _18972_, _18967_);
  nor (_18974_, _04896_, _08642_);
  or (_18975_, _18974_, _18951_);
  or (_18977_, _18975_, _03327_);
  and (_18978_, _18977_, _18973_);
  or (_18979_, _18978_, _02950_);
  or (_18980_, _18960_, _02959_);
  and (_18981_, _18980_, _02888_);
  and (_18982_, _18981_, _18979_);
  and (_18983_, _11442_, _05346_);
  or (_18984_, _18983_, _18968_);
  and (_18985_, _18984_, _02887_);
  or (_18986_, _18985_, _02880_);
  or (_18988_, _18986_, _18982_);
  or (_18989_, _18968_, _11474_);
  and (_18990_, _18989_, _18970_);
  or (_18991_, _18990_, _02881_);
  and (_18992_, _18991_, _02875_);
  and (_18993_, _18992_, _18988_);
  and (_18994_, _17409_, _05346_);
  or (_18995_, _18994_, _18968_);
  and (_18996_, _18995_, _02874_);
  or (_18997_, _18996_, _06793_);
  or (_18999_, _18997_, _18993_);
  or (_19000_, _18975_, _06241_);
  and (_19001_, _19000_, _18999_);
  or (_19002_, _19001_, _02855_);
  and (_19003_, _06180_, _04722_);
  or (_19004_, _18951_, _02856_);
  or (_19005_, _19004_, _19003_);
  and (_19006_, _19005_, _02851_);
  and (_19007_, _19006_, _19002_);
  and (_19008_, _17436_, _04722_);
  or (_19010_, _19008_, _18951_);
  and (_19011_, _19010_, _02576_);
  or (_19012_, _19011_, _03014_);
  or (_19013_, _19012_, _19007_);
  and (_19014_, _05701_, _04722_);
  or (_19015_, _19014_, _18951_);
  or (_19016_, _19015_, _03884_);
  and (_19017_, _19016_, _19013_);
  or (_19018_, _19017_, _03021_);
  and (_19019_, _11562_, _04722_);
  or (_19021_, _18951_, _05279_);
  or (_19022_, _19021_, _19019_);
  and (_19023_, _19022_, _03131_);
  and (_19024_, _19023_, _19018_);
  or (_19025_, _19024_, _18955_);
  and (_19026_, _19025_, _05274_);
  or (_19027_, _18951_, _04944_);
  and (_19028_, _19015_, _03020_);
  and (_19029_, _19028_, _19027_);
  or (_19030_, _19029_, _19026_);
  and (_19032_, _19030_, _03140_);
  and (_19033_, _18960_, _03139_);
  and (_19034_, _19033_, _19027_);
  or (_19035_, _19034_, _03036_);
  or (_19036_, _19035_, _19032_);
  nor (_19037_, _11560_, _08642_);
  or (_19038_, _18951_, _05781_);
  or (_19039_, _19038_, _19037_);
  and (_19040_, _19039_, _05786_);
  and (_19041_, _19040_, _19036_);
  nor (_19043_, _11435_, _08642_);
  or (_19044_, _19043_, _18951_);
  and (_19045_, _19044_, _03127_);
  or (_19046_, _19045_, _03166_);
  or (_19047_, _19046_, _19041_);
  or (_19048_, _18957_, _03563_);
  and (_19049_, _19048_, _02501_);
  and (_19050_, _19049_, _19047_);
  and (_19051_, _18984_, _02500_);
  or (_19052_, _19051_, _03174_);
  or (_19054_, _19052_, _19050_);
  and (_19055_, _11619_, _04722_);
  or (_19056_, _18951_, _03178_);
  or (_19057_, _19056_, _19055_);
  and (_19058_, _19057_, _34698_);
  and (_19059_, _19058_, _19054_);
  or (_35227_, _19059_, _18950_);
  not (_19060_, \oc8051_golden_model_1.P2 [6]);
  nor (_19061_, _34698_, _19060_);
  or (_19062_, _19061_, rst);
  nor (_19064_, _04722_, _19060_);
  and (_19065_, _11769_, _04722_);
  or (_19066_, _19065_, _19064_);
  and (_19067_, _19066_, _03130_);
  nor (_19068_, _11636_, _08642_);
  or (_19069_, _19068_, _19064_);
  or (_19070_, _19069_, _03821_);
  and (_19071_, _04722_, \oc8051_golden_model_1.ACC [6]);
  or (_19072_, _19071_, _19064_);
  and (_19073_, _19072_, _03825_);
  nor (_19075_, _03825_, _19060_);
  or (_19076_, _19075_, _02952_);
  or (_19077_, _19076_, _19073_);
  and (_19078_, _19077_, _02892_);
  and (_19079_, _19078_, _19070_);
  nor (_19080_, _05346_, _19060_);
  and (_19081_, _11653_, _05346_);
  or (_19082_, _19081_, _19080_);
  and (_19083_, _19082_, _02891_);
  or (_19084_, _19083_, _02947_);
  or (_19086_, _19084_, _19079_);
  nor (_19087_, _04787_, _08642_);
  or (_19088_, _19087_, _19064_);
  or (_19089_, _19088_, _03327_);
  and (_19090_, _19089_, _19086_);
  or (_19091_, _19090_, _02950_);
  or (_19092_, _19072_, _02959_);
  and (_19093_, _19092_, _02888_);
  and (_19094_, _19093_, _19091_);
  and (_19095_, _11675_, _05346_);
  or (_19097_, _19095_, _19080_);
  and (_19098_, _19097_, _02887_);
  or (_19099_, _19098_, _02880_);
  or (_19100_, _19099_, _19094_);
  or (_19101_, _19080_, _11682_);
  and (_19102_, _19101_, _19082_);
  or (_19103_, _19102_, _02881_);
  and (_19104_, _19103_, _02875_);
  and (_19105_, _19104_, _19100_);
  and (_19106_, _17535_, _05346_);
  or (_19108_, _19106_, _19080_);
  and (_19109_, _19108_, _02874_);
  or (_19110_, _19109_, _06793_);
  or (_19111_, _19110_, _19105_);
  or (_19112_, _19088_, _06241_);
  and (_19113_, _19112_, _19111_);
  or (_19114_, _19113_, _02855_);
  and (_19115_, _05847_, _04722_);
  or (_19116_, _19064_, _02856_);
  or (_19117_, _19116_, _19115_);
  and (_19119_, _19117_, _02851_);
  and (_19120_, _19119_, _19114_);
  and (_19121_, _17563_, _04722_);
  or (_19122_, _19121_, _19064_);
  and (_19123_, _19122_, _02576_);
  or (_19124_, _19123_, _03014_);
  or (_19125_, _19124_, _19120_);
  and (_19126_, _11758_, _04722_);
  or (_19127_, _19126_, _19064_);
  or (_19128_, _19127_, _03884_);
  and (_19130_, _19128_, _19125_);
  or (_19131_, _19130_, _03021_);
  and (_19132_, _11646_, _04722_);
  or (_19133_, _19064_, _05279_);
  or (_19134_, _19133_, _19132_);
  and (_19135_, _19134_, _03131_);
  and (_19136_, _19135_, _19131_);
  or (_19137_, _19136_, _19067_);
  and (_19138_, _19137_, _05274_);
  or (_19139_, _19064_, _04838_);
  and (_19141_, _19127_, _03020_);
  and (_19142_, _19141_, _19139_);
  or (_19143_, _19142_, _19138_);
  and (_19144_, _19143_, _03140_);
  and (_19145_, _19072_, _03139_);
  and (_19146_, _19145_, _19139_);
  or (_19147_, _19146_, _03036_);
  or (_19148_, _19147_, _19144_);
  nor (_19149_, _11644_, _08642_);
  or (_19150_, _19064_, _05781_);
  or (_19152_, _19150_, _19149_);
  and (_19153_, _19152_, _05786_);
  and (_19154_, _19153_, _19148_);
  nor (_19155_, _11768_, _08642_);
  or (_19156_, _19155_, _19064_);
  and (_19157_, _19156_, _03127_);
  or (_19158_, _19157_, _03166_);
  or (_19159_, _19158_, _19154_);
  or (_19160_, _19069_, _03563_);
  and (_19161_, _19160_, _02501_);
  and (_19163_, _19161_, _19159_);
  and (_19164_, _19097_, _02500_);
  or (_19165_, _19164_, _03174_);
  or (_19166_, _19165_, _19163_);
  and (_19167_, _11821_, _04722_);
  or (_19168_, _19064_, _03178_);
  or (_19169_, _19168_, _19167_);
  and (_19170_, _19169_, _34698_);
  and (_19171_, _19170_, _19166_);
  or (_35228_, _19171_, _19062_);
  not (_19173_, \oc8051_golden_model_1.P3 [0]);
  nor (_19174_, _34698_, _19173_);
  or (_19175_, _19174_, rst);
  nor (_19176_, _04724_, _19173_);
  and (_19177_, _10546_, _04724_);
  or (_19178_, _19177_, _19176_);
  and (_19179_, _19178_, _03130_);
  and (_19180_, _04724_, _03817_);
  or (_19181_, _19180_, _19176_);
  or (_19182_, _19181_, _06241_);
  and (_19184_, _05044_, _04724_);
  or (_19185_, _19184_, _19176_);
  or (_19186_, _19185_, _03821_);
  and (_19187_, _04724_, \oc8051_golden_model_1.ACC [0]);
  or (_19188_, _19187_, _19176_);
  and (_19189_, _19188_, _03825_);
  nor (_19190_, _03825_, _19173_);
  or (_19191_, _19190_, _02952_);
  or (_19192_, _19191_, _19189_);
  and (_19193_, _19192_, _02892_);
  and (_19195_, _19193_, _19186_);
  nor (_19196_, _05357_, _19173_);
  and (_19197_, _10429_, _05357_);
  or (_19198_, _19197_, _19196_);
  and (_19199_, _19198_, _02891_);
  or (_19200_, _19199_, _19195_);
  and (_19201_, _19200_, _03327_);
  and (_19202_, _19181_, _02947_);
  or (_19203_, _19202_, _02950_);
  or (_19204_, _19203_, _19201_);
  or (_19206_, _19188_, _02959_);
  and (_19207_, _19206_, _02888_);
  and (_19208_, _19207_, _19204_);
  and (_19209_, _19176_, _02887_);
  or (_19210_, _19209_, _02880_);
  or (_19211_, _19210_, _19208_);
  or (_19212_, _19185_, _02881_);
  and (_19213_, _19212_, _02875_);
  and (_19214_, _19213_, _19211_);
  and (_19215_, _16789_, _05357_);
  or (_19217_, _19215_, _19196_);
  and (_19218_, _19217_, _02874_);
  or (_19219_, _19218_, _06793_);
  or (_19220_, _19219_, _19214_);
  and (_19221_, _19220_, _19182_);
  or (_19222_, _19221_, _02855_);
  and (_19223_, _06174_, _04724_);
  or (_19224_, _19176_, _02856_);
  or (_19225_, _19224_, _19223_);
  and (_19226_, _19225_, _02851_);
  and (_19228_, _19226_, _19222_);
  and (_19229_, _16814_, _04724_);
  or (_19230_, _19229_, _19176_);
  and (_19231_, _19230_, _02576_);
  or (_19232_, _19231_, _03014_);
  or (_19233_, _19232_, _19228_);
  and (_19234_, _04724_, _05566_);
  or (_19235_, _19234_, _19176_);
  or (_19236_, _19235_, _03884_);
  and (_19237_, _19236_, _19233_);
  or (_19239_, _19237_, _03021_);
  and (_19240_, _10425_, _04724_);
  or (_19241_, _19176_, _05279_);
  or (_19242_, _19241_, _19240_);
  and (_19243_, _19242_, _03131_);
  and (_19244_, _19243_, _19239_);
  or (_19245_, _19244_, _19179_);
  and (_19246_, _19245_, _05274_);
  nand (_19247_, _19235_, _03020_);
  nor (_19248_, _19247_, _19184_);
  or (_19250_, _19248_, _19246_);
  and (_19251_, _19250_, _03140_);
  or (_19252_, _19176_, _09183_);
  and (_19253_, _19188_, _03139_);
  and (_19254_, _19253_, _19252_);
  or (_19255_, _19254_, _03036_);
  or (_19256_, _19255_, _19251_);
  nor (_19257_, _10423_, _08745_);
  or (_19258_, _19176_, _05781_);
  or (_19259_, _19258_, _19257_);
  and (_19261_, _19259_, _05786_);
  and (_19262_, _19261_, _19256_);
  nor (_19263_, _10421_, _08745_);
  or (_19264_, _19263_, _19176_);
  and (_19265_, _19264_, _03127_);
  or (_19266_, _19265_, _03166_);
  or (_19267_, _19266_, _19262_);
  or (_19268_, _19185_, _03563_);
  and (_19269_, _19268_, _02501_);
  and (_19270_, _19269_, _19267_);
  and (_19272_, _19176_, _02500_);
  or (_19273_, _19272_, _03174_);
  or (_19274_, _19273_, _19270_);
  or (_19275_, _19185_, _03178_);
  and (_19276_, _19275_, _34698_);
  and (_19277_, _19276_, _19274_);
  or (_35229_, _19277_, _19175_);
  not (_19278_, \oc8051_golden_model_1.P3 [1]);
  nor (_19279_, _34698_, _19278_);
  or (_19280_, _19279_, rst);
  nand (_19282_, _04724_, _03705_);
  or (_19283_, _04724_, \oc8051_golden_model_1.P3 [1]);
  and (_19284_, _19283_, _03014_);
  and (_19285_, _19284_, _19282_);
  or (_19286_, _16935_, _08745_);
  and (_19287_, _19283_, _02576_);
  and (_19288_, _19287_, _19286_);
  and (_19289_, _10622_, _04724_);
  not (_19290_, _19289_);
  and (_19291_, _19290_, _19283_);
  or (_19293_, _19291_, _03821_);
  nand (_19294_, _04724_, _02618_);
  and (_19295_, _19294_, _19283_);
  and (_19296_, _19295_, _03825_);
  nor (_19297_, _03825_, _19278_);
  or (_19298_, _19297_, _02952_);
  or (_19299_, _19298_, _19296_);
  and (_19300_, _19299_, _02892_);
  and (_19301_, _19300_, _19293_);
  and (_19302_, _10617_, _05357_);
  nor (_19304_, _05357_, _19278_);
  or (_19305_, _19304_, _02947_);
  or (_19306_, _19305_, _19302_);
  and (_19307_, _19306_, _09918_);
  or (_19308_, _19307_, _19301_);
  nor (_19309_, _04724_, _19278_);
  and (_19310_, _04724_, _04005_);
  or (_19311_, _19310_, _19309_);
  or (_19312_, _19311_, _03327_);
  and (_19313_, _19312_, _19308_);
  or (_19315_, _19313_, _02950_);
  or (_19316_, _19295_, _02959_);
  and (_19317_, _19316_, _02888_);
  and (_19318_, _19317_, _19315_);
  and (_19319_, _10620_, _05357_);
  or (_19320_, _19319_, _19304_);
  and (_19321_, _19320_, _02887_);
  or (_19322_, _19321_, _02880_);
  or (_19323_, _19322_, _19318_);
  and (_19324_, _19302_, _10616_);
  or (_19326_, _19304_, _02881_);
  or (_19327_, _19326_, _19324_);
  and (_19328_, _19327_, _19323_);
  and (_19329_, _19328_, _02875_);
  and (_19330_, _16909_, _05357_);
  or (_19331_, _19304_, _19330_);
  and (_19332_, _19331_, _02874_);
  or (_19333_, _19332_, _06793_);
  or (_19334_, _19333_, _19329_);
  or (_19335_, _19311_, _06241_);
  and (_19337_, _19335_, _19334_);
  or (_19338_, _19337_, _02855_);
  and (_19339_, _06173_, _04724_);
  or (_19340_, _19309_, _02856_);
  or (_19341_, _19340_, _19339_);
  and (_19342_, _19341_, _02851_);
  and (_19343_, _19342_, _19338_);
  or (_19344_, _19343_, _19288_);
  and (_19345_, _19344_, _03884_);
  or (_19346_, _19345_, _19285_);
  and (_19348_, _19346_, _05279_);
  or (_19349_, _10612_, _08745_);
  and (_19350_, _19283_, _03021_);
  and (_19351_, _19350_, _19349_);
  or (_19352_, _19351_, _19348_);
  and (_19353_, _19352_, _03131_);
  or (_19354_, _10739_, _08745_);
  and (_19355_, _19283_, _03130_);
  and (_19356_, _19355_, _19354_);
  or (_19357_, _19356_, _19353_);
  and (_19359_, _19357_, _05274_);
  or (_19360_, _10611_, _08745_);
  and (_19361_, _19283_, _03020_);
  and (_19362_, _19361_, _19360_);
  or (_19363_, _19362_, _19359_);
  and (_19364_, _19363_, _03140_);
  or (_19365_, _19309_, _12724_);
  and (_19366_, _19295_, _03139_);
  and (_19367_, _19366_, _19365_);
  or (_19368_, _19367_, _19364_);
  and (_19370_, _19368_, _03128_);
  or (_19371_, _19294_, _12724_);
  and (_19372_, _19283_, _03127_);
  and (_19373_, _19372_, _19371_);
  or (_19374_, _19373_, _03166_);
  or (_19375_, _19282_, _12724_);
  and (_19376_, _19283_, _03036_);
  and (_19377_, _19376_, _19375_);
  or (_19378_, _19377_, _19374_);
  or (_19379_, _19378_, _19370_);
  or (_19381_, _19291_, _03563_);
  and (_19382_, _19381_, _02501_);
  and (_19383_, _19382_, _19379_);
  and (_19384_, _19320_, _02500_);
  or (_19385_, _19384_, _03174_);
  or (_19386_, _19385_, _19383_);
  or (_19387_, _19309_, _03178_);
  or (_19388_, _19387_, _19289_);
  and (_19389_, _19388_, _34698_);
  and (_19390_, _19389_, _19386_);
  or (_35231_, _19390_, _19280_);
  not (_19392_, \oc8051_golden_model_1.P3 [2]);
  nor (_19393_, _34698_, _19392_);
  or (_19394_, _19393_, rst);
  nor (_19395_, _04724_, _19392_);
  and (_19396_, _10831_, _04724_);
  or (_19397_, _19396_, _19395_);
  and (_19398_, _19397_, _03130_);
  nor (_19399_, _08745_, _04440_);
  or (_19400_, _19399_, _19395_);
  or (_19402_, _19400_, _06241_);
  or (_19403_, _19400_, _03327_);
  nor (_19404_, _10849_, _08745_);
  or (_19405_, _19404_, _19395_);
  or (_19406_, _19405_, _03821_);
  and (_19407_, _04724_, \oc8051_golden_model_1.ACC [2]);
  or (_19408_, _19407_, _19395_);
  and (_19409_, _19408_, _03825_);
  nor (_19410_, _03825_, _19392_);
  or (_19411_, _19410_, _02952_);
  or (_19413_, _19411_, _19409_);
  and (_19414_, _19413_, _02892_);
  and (_19415_, _19414_, _19406_);
  nor (_19416_, _05357_, _19392_);
  and (_19417_, _10853_, _05357_);
  or (_19418_, _19417_, _19416_);
  and (_19419_, _19418_, _02891_);
  or (_19420_, _19419_, _02947_);
  or (_19421_, _19420_, _19415_);
  and (_19422_, _19421_, _19403_);
  or (_19424_, _19422_, _02950_);
  or (_19425_, _19408_, _02959_);
  and (_19426_, _19425_, _02888_);
  and (_19427_, _19426_, _19424_);
  and (_19428_, _10838_, _05357_);
  or (_19429_, _19428_, _19416_);
  and (_19430_, _19429_, _02887_);
  or (_19431_, _19430_, _02880_);
  or (_19432_, _19431_, _19427_);
  and (_19433_, _19417_, _10868_);
  or (_19435_, _19416_, _02881_);
  or (_19436_, _19435_, _19433_);
  and (_19437_, _19436_, _02875_);
  and (_19438_, _19437_, _19432_);
  and (_19439_, _17034_, _05357_);
  or (_19440_, _19439_, _19416_);
  and (_19441_, _19440_, _02874_);
  or (_19442_, _19441_, _06793_);
  or (_19443_, _19442_, _19438_);
  and (_19444_, _19443_, _19402_);
  or (_19446_, _19444_, _02855_);
  and (_19447_, _06177_, _04724_);
  or (_19448_, _19395_, _02856_);
  or (_19449_, _19448_, _19447_);
  and (_19450_, _19449_, _02851_);
  and (_19451_, _19450_, _19446_);
  and (_19452_, _17060_, _04724_);
  or (_19453_, _19452_, _19395_);
  and (_19454_, _19453_, _02576_);
  or (_19455_, _19454_, _03014_);
  or (_19457_, _19455_, _19451_);
  and (_19458_, _04724_, _05727_);
  or (_19459_, _19458_, _19395_);
  or (_19460_, _19459_, _03884_);
  and (_19461_, _19460_, _19457_);
  or (_19462_, _19461_, _03021_);
  and (_19463_, _10835_, _04724_);
  or (_19464_, _19395_, _05279_);
  or (_19465_, _19464_, _19463_);
  and (_19466_, _19465_, _03131_);
  and (_19468_, _19466_, _19462_);
  or (_19469_, _19468_, _19398_);
  and (_19470_, _19469_, _05274_);
  or (_19471_, _19395_, _05143_);
  and (_19472_, _19459_, _03020_);
  and (_19473_, _19472_, _19471_);
  or (_19474_, _19473_, _19470_);
  and (_19475_, _19474_, _03140_);
  and (_19476_, _19408_, _03139_);
  and (_19477_, _19476_, _19471_);
  or (_19479_, _19477_, _03036_);
  or (_19480_, _19479_, _19475_);
  nor (_19481_, _10833_, _08745_);
  or (_19482_, _19395_, _05781_);
  or (_19483_, _19482_, _19481_);
  and (_19484_, _19483_, _05786_);
  and (_19485_, _19484_, _19480_);
  nor (_19486_, _10830_, _08745_);
  or (_19487_, _19486_, _19395_);
  and (_19488_, _19487_, _03127_);
  or (_19490_, _19488_, _03166_);
  or (_19491_, _19490_, _19485_);
  or (_19492_, _19405_, _03563_);
  and (_19493_, _19492_, _02501_);
  and (_19494_, _19493_, _19491_);
  and (_19495_, _19429_, _02500_);
  or (_19496_, _19495_, _03174_);
  or (_19497_, _19496_, _19494_);
  and (_19498_, _11008_, _04724_);
  or (_19499_, _19395_, _03178_);
  or (_19501_, _19499_, _19498_);
  and (_19502_, _19501_, _34698_);
  and (_19503_, _19502_, _19497_);
  or (_35232_, _19503_, _19394_);
  nor (_19504_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_19505_, _19504_, _04548_);
  and (_19506_, _08745_, \oc8051_golden_model_1.P3 [3]);
  and (_19507_, _11028_, _04724_);
  or (_19508_, _19507_, _19506_);
  and (_19509_, _19508_, _03130_);
  nor (_19510_, _08745_, _04242_);
  or (_19511_, _19510_, _19506_);
  or (_19512_, _19511_, _06241_);
  nor (_19513_, _11040_, _08745_);
  or (_19514_, _19513_, _19506_);
  or (_19515_, _19514_, _03821_);
  and (_19516_, _04724_, \oc8051_golden_model_1.ACC [3]);
  or (_19517_, _19516_, _19506_);
  and (_19518_, _19517_, _03825_);
  and (_19519_, _03826_, \oc8051_golden_model_1.P3 [3]);
  or (_19521_, _19519_, _02952_);
  or (_19522_, _19521_, _19518_);
  and (_19523_, _19522_, _02892_);
  and (_19524_, _19523_, _19515_);
  not (_19525_, _05357_);
  and (_19526_, _19525_, \oc8051_golden_model_1.P3 [3]);
  and (_19527_, _11037_, _05357_);
  or (_19528_, _19527_, _19526_);
  and (_19529_, _19528_, _02891_);
  or (_19530_, _19529_, _02947_);
  or (_19532_, _19530_, _19524_);
  or (_19533_, _19511_, _03327_);
  and (_19534_, _19533_, _19532_);
  or (_19535_, _19534_, _02950_);
  or (_19536_, _19517_, _02959_);
  and (_19537_, _19536_, _02888_);
  and (_19538_, _19537_, _19535_);
  and (_19539_, _11035_, _05357_);
  or (_19540_, _19539_, _19526_);
  and (_19541_, _19540_, _02887_);
  or (_19543_, _19541_, _02880_);
  or (_19544_, _19543_, _19538_);
  or (_19545_, _19526_, _11066_);
  and (_19546_, _19545_, _19528_);
  or (_19547_, _19546_, _02881_);
  and (_19548_, _19547_, _02875_);
  and (_19549_, _19548_, _19544_);
  and (_19550_, _17160_, _05357_);
  or (_19551_, _19550_, _19526_);
  and (_19552_, _19551_, _02874_);
  or (_19553_, _19552_, _06793_);
  or (_19554_, _19553_, _19549_);
  and (_19555_, _19554_, _19512_);
  or (_19556_, _19555_, _02855_);
  and (_19557_, _06176_, _04724_);
  or (_19558_, _19506_, _02856_);
  or (_19559_, _19558_, _19557_);
  and (_19560_, _19559_, _02851_);
  and (_19561_, _19560_, _19556_);
  and (_19562_, _17185_, _04724_);
  or (_19564_, _19562_, _19506_);
  and (_19565_, _19564_, _02576_);
  or (_19566_, _19565_, _03014_);
  or (_19567_, _19566_, _19561_);
  and (_19568_, _04724_, _05664_);
  or (_19569_, _19568_, _19506_);
  or (_19570_, _19569_, _03884_);
  and (_19571_, _19570_, _19567_);
  or (_19572_, _19571_, _03021_);
  and (_19573_, _11032_, _04724_);
  or (_19574_, _19506_, _05279_);
  or (_19575_, _19574_, _19573_);
  and (_19576_, _19575_, _03131_);
  and (_19577_, _19576_, _19572_);
  or (_19578_, _19577_, _19509_);
  and (_19579_, _19578_, _05274_);
  or (_19580_, _19506_, _04996_);
  and (_19581_, _19569_, _03020_);
  and (_19582_, _19581_, _19580_);
  or (_19583_, _19582_, _19579_);
  and (_19585_, _19583_, _03140_);
  and (_19586_, _19517_, _03139_);
  and (_19587_, _19586_, _19580_);
  or (_19588_, _19587_, _03036_);
  or (_19589_, _19588_, _19585_);
  nor (_19590_, _11030_, _08745_);
  or (_19591_, _19506_, _05781_);
  or (_19592_, _19591_, _19590_);
  and (_19593_, _19592_, _05786_);
  and (_19594_, _19593_, _19589_);
  nor (_19596_, _11027_, _08745_);
  or (_19597_, _19596_, _19506_);
  and (_19598_, _19597_, _03127_);
  or (_19599_, _19598_, _03166_);
  or (_19600_, _19599_, _19594_);
  or (_19601_, _19514_, _03563_);
  and (_19602_, _19601_, _02501_);
  and (_19603_, _19602_, _19600_);
  and (_19604_, _19540_, _02500_);
  or (_19605_, _19604_, _03174_);
  or (_19606_, _19605_, _19603_);
  and (_19607_, _11213_, _04724_);
  or (_19608_, _19506_, _03178_);
  or (_19609_, _19608_, _19607_);
  and (_19610_, _19609_, _34698_);
  and (_19611_, _19610_, _19606_);
  or (_35233_, _19611_, _19505_);
  nor (_19612_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_19613_, _19612_, _04548_);
  and (_19614_, _08745_, \oc8051_golden_model_1.P3 [4]);
  and (_19616_, _11368_, _04724_);
  or (_19617_, _19616_, _19614_);
  and (_19618_, _19617_, _03130_);
  nor (_19619_, _05202_, _08745_);
  or (_19620_, _19619_, _19614_);
  or (_19621_, _19620_, _06241_);
  and (_19622_, _19525_, \oc8051_golden_model_1.P3 [4]);
  and (_19623_, _11243_, _05357_);
  or (_19624_, _19623_, _19622_);
  and (_19625_, _19624_, _02887_);
  nor (_19627_, _11259_, _08745_);
  or (_19628_, _19627_, _19614_);
  or (_19629_, _19628_, _03821_);
  and (_19630_, _04724_, \oc8051_golden_model_1.ACC [4]);
  or (_19631_, _19630_, _19614_);
  and (_19632_, _19631_, _03825_);
  and (_19633_, _03826_, \oc8051_golden_model_1.P3 [4]);
  or (_19634_, _19633_, _02952_);
  or (_19635_, _19634_, _19632_);
  and (_19636_, _19635_, _02892_);
  and (_19637_, _19636_, _19629_);
  and (_19638_, _11245_, _05357_);
  or (_19639_, _19638_, _19622_);
  and (_19640_, _19639_, _02891_);
  or (_19641_, _19640_, _02947_);
  or (_19642_, _19641_, _19637_);
  or (_19643_, _19620_, _03327_);
  and (_19644_, _19643_, _19642_);
  or (_19645_, _19644_, _02950_);
  or (_19646_, _19631_, _02959_);
  and (_19648_, _19646_, _02888_);
  and (_19649_, _19648_, _19645_);
  or (_19650_, _19649_, _19625_);
  and (_19651_, _19650_, _02881_);
  or (_19652_, _19622_, _11276_);
  and (_19653_, _19652_, _02880_);
  and (_19654_, _19653_, _19639_);
  or (_19655_, _19654_, _19651_);
  and (_19656_, _19655_, _02875_);
  and (_19657_, _17285_, _05357_);
  or (_19659_, _19657_, _19622_);
  and (_19660_, _19659_, _02874_);
  or (_19661_, _19660_, _06793_);
  or (_19662_, _19661_, _19656_);
  and (_19663_, _19662_, _19621_);
  or (_19664_, _19663_, _02855_);
  and (_19665_, _06181_, _04724_);
  or (_19666_, _19614_, _02856_);
  or (_19667_, _19666_, _19665_);
  and (_19668_, _19667_, _02851_);
  and (_19669_, _19668_, _19664_);
  and (_19670_, _17311_, _04724_);
  or (_19671_, _19670_, _19614_);
  and (_19672_, _19671_, _02576_);
  or (_19673_, _19672_, _03014_);
  or (_19674_, _19673_, _19669_);
  and (_19675_, _05697_, _04724_);
  or (_19676_, _19675_, _19614_);
  or (_19677_, _19676_, _03884_);
  and (_19678_, _19677_, _19674_);
  or (_19680_, _19678_, _03021_);
  and (_19681_, _11362_, _04724_);
  or (_19682_, _19614_, _05279_);
  or (_19683_, _19682_, _19681_);
  and (_19684_, _19683_, _03131_);
  and (_19685_, _19684_, _19680_);
  or (_19686_, _19685_, _19618_);
  and (_19687_, _19686_, _05274_);
  or (_19688_, _19614_, _05251_);
  and (_19689_, _19676_, _03020_);
  and (_19691_, _19689_, _19688_);
  or (_19692_, _19691_, _19687_);
  and (_19693_, _19692_, _03140_);
  and (_19694_, _19631_, _03139_);
  and (_19695_, _19694_, _19688_);
  or (_19696_, _19695_, _03036_);
  or (_19697_, _19696_, _19693_);
  nor (_19698_, _11361_, _08745_);
  or (_19699_, _19614_, _05781_);
  or (_19700_, _19699_, _19698_);
  and (_19701_, _19700_, _05786_);
  and (_19702_, _19701_, _19697_);
  nor (_19703_, _11367_, _08745_);
  or (_19704_, _19703_, _19614_);
  and (_19705_, _19704_, _03127_);
  or (_19706_, _19705_, _03166_);
  or (_19707_, _19706_, _19702_);
  or (_19708_, _19628_, _03563_);
  and (_19709_, _19708_, _02501_);
  and (_19710_, _19709_, _19707_);
  and (_19712_, _19624_, _02500_);
  or (_19713_, _19712_, _03174_);
  or (_19714_, _19713_, _19710_);
  and (_19715_, _11417_, _04724_);
  or (_19716_, _19614_, _03178_);
  or (_19717_, _19716_, _19715_);
  and (_19718_, _19717_, _34698_);
  and (_19719_, _19718_, _19714_);
  or (_35234_, _19719_, _19613_);
  nor (_19720_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_19722_, _19720_, _04548_);
  and (_19723_, _08745_, \oc8051_golden_model_1.P3 [5]);
  and (_19724_, _11436_, _04724_);
  or (_19725_, _19724_, _19723_);
  and (_19726_, _19725_, _03130_);
  nor (_19727_, _11445_, _08745_);
  or (_19728_, _19727_, _19723_);
  or (_19729_, _19728_, _03821_);
  and (_19730_, _04724_, \oc8051_golden_model_1.ACC [5]);
  or (_19731_, _19730_, _19723_);
  and (_19732_, _19731_, _03825_);
  and (_19733_, _03826_, \oc8051_golden_model_1.P3 [5]);
  or (_19734_, _19733_, _02952_);
  or (_19735_, _19734_, _19732_);
  and (_19736_, _19735_, _02892_);
  and (_19737_, _19736_, _19729_);
  and (_19738_, _19525_, \oc8051_golden_model_1.P3 [5]);
  and (_19739_, _11459_, _05357_);
  or (_19740_, _19739_, _19738_);
  and (_19741_, _19740_, _02891_);
  or (_19743_, _19741_, _02947_);
  or (_19744_, _19743_, _19737_);
  nor (_19745_, _04896_, _08745_);
  or (_19746_, _19745_, _19723_);
  or (_19747_, _19746_, _03327_);
  and (_19748_, _19747_, _19744_);
  or (_19749_, _19748_, _02950_);
  or (_19750_, _19731_, _02959_);
  and (_19751_, _19750_, _02888_);
  and (_19752_, _19751_, _19749_);
  and (_19754_, _11442_, _05357_);
  or (_19755_, _19754_, _19738_);
  and (_19756_, _19755_, _02887_);
  or (_19757_, _19756_, _02880_);
  or (_19758_, _19757_, _19752_);
  or (_19759_, _19738_, _11474_);
  and (_19760_, _19759_, _19740_);
  or (_19761_, _19760_, _02881_);
  and (_19762_, _19761_, _02875_);
  and (_19763_, _19762_, _19758_);
  and (_19764_, _17409_, _05357_);
  or (_19765_, _19764_, _19738_);
  and (_19766_, _19765_, _02874_);
  or (_19767_, _19766_, _06793_);
  or (_19768_, _19767_, _19763_);
  or (_19769_, _19746_, _06241_);
  and (_19770_, _19769_, _19768_);
  or (_19771_, _19770_, _02855_);
  and (_19772_, _06180_, _04724_);
  or (_19773_, _19723_, _02856_);
  or (_19775_, _19773_, _19772_);
  and (_19776_, _19775_, _02851_);
  and (_19777_, _19776_, _19771_);
  and (_19778_, _17436_, _04724_);
  or (_19779_, _19778_, _19723_);
  and (_19780_, _19779_, _02576_);
  or (_19781_, _19780_, _03014_);
  or (_19782_, _19781_, _19777_);
  and (_19783_, _05701_, _04724_);
  or (_19784_, _19783_, _19723_);
  or (_19786_, _19784_, _03884_);
  and (_19787_, _19786_, _19782_);
  or (_19788_, _19787_, _03021_);
  and (_19789_, _11562_, _04724_);
  or (_19790_, _19723_, _05279_);
  or (_19791_, _19790_, _19789_);
  and (_19792_, _19791_, _03131_);
  and (_19793_, _19792_, _19788_);
  or (_19794_, _19793_, _19726_);
  and (_19795_, _19794_, _05274_);
  or (_19796_, _19723_, _04944_);
  and (_19797_, _19784_, _03020_);
  and (_19798_, _19797_, _19796_);
  or (_19799_, _19798_, _19795_);
  and (_19800_, _19799_, _03140_);
  and (_19801_, _19731_, _03139_);
  and (_19802_, _19801_, _19796_);
  or (_19803_, _19802_, _03036_);
  or (_19804_, _19803_, _19800_);
  nor (_19805_, _11560_, _08745_);
  or (_19807_, _19723_, _05781_);
  or (_19808_, _19807_, _19805_);
  and (_19809_, _19808_, _05786_);
  and (_19810_, _19809_, _19804_);
  nor (_19811_, _11435_, _08745_);
  or (_19812_, _19811_, _19723_);
  and (_19813_, _19812_, _03127_);
  or (_19814_, _19813_, _03166_);
  or (_19815_, _19814_, _19810_);
  or (_19816_, _19728_, _03563_);
  and (_19818_, _19816_, _02501_);
  and (_19819_, _19818_, _19815_);
  and (_19820_, _19755_, _02500_);
  or (_19821_, _19820_, _03174_);
  or (_19822_, _19821_, _19819_);
  and (_19823_, _11619_, _04724_);
  or (_19824_, _19723_, _03178_);
  or (_19825_, _19824_, _19823_);
  and (_19826_, _19825_, _34698_);
  and (_19827_, _19826_, _19822_);
  or (_35235_, _19827_, _19722_);
  not (_19828_, \oc8051_golden_model_1.P3 [6]);
  nor (_19829_, _34698_, _19828_);
  or (_19830_, _19829_, rst);
  nor (_19831_, _04724_, _19828_);
  and (_19832_, _11769_, _04724_);
  or (_19833_, _19832_, _19831_);
  and (_19834_, _19833_, _03130_);
  nor (_19835_, _11636_, _08745_);
  or (_19836_, _19835_, _19831_);
  or (_19838_, _19836_, _03821_);
  and (_19839_, _04724_, \oc8051_golden_model_1.ACC [6]);
  or (_19840_, _19839_, _19831_);
  and (_19841_, _19840_, _03825_);
  nor (_19842_, _03825_, _19828_);
  or (_19843_, _19842_, _02952_);
  or (_19844_, _19843_, _19841_);
  and (_19845_, _19844_, _02892_);
  and (_19846_, _19845_, _19838_);
  nor (_19847_, _05357_, _19828_);
  and (_19849_, _11653_, _05357_);
  or (_19850_, _19849_, _19847_);
  and (_19851_, _19850_, _02891_);
  or (_19852_, _19851_, _02947_);
  or (_19853_, _19852_, _19846_);
  nor (_19854_, _04787_, _08745_);
  or (_19855_, _19854_, _19831_);
  or (_19856_, _19855_, _03327_);
  and (_19857_, _19856_, _19853_);
  or (_19858_, _19857_, _02950_);
  or (_19859_, _19840_, _02959_);
  and (_19860_, _19859_, _02888_);
  and (_19861_, _19860_, _19858_);
  and (_19862_, _11675_, _05357_);
  or (_19863_, _19862_, _19847_);
  and (_19864_, _19863_, _02887_);
  or (_19865_, _19864_, _02880_);
  or (_19866_, _19865_, _19861_);
  or (_19867_, _19847_, _11682_);
  and (_19868_, _19867_, _19850_);
  or (_19870_, _19868_, _02881_);
  and (_19871_, _19870_, _02875_);
  and (_19872_, _19871_, _19866_);
  and (_19873_, _17535_, _05357_);
  or (_19874_, _19873_, _19847_);
  and (_19875_, _19874_, _02874_);
  or (_19876_, _19875_, _06793_);
  or (_19877_, _19876_, _19872_);
  or (_19878_, _19855_, _06241_);
  and (_19879_, _19878_, _19877_);
  or (_19881_, _19879_, _02855_);
  and (_19882_, _05847_, _04724_);
  or (_19883_, _19831_, _02856_);
  or (_19884_, _19883_, _19882_);
  and (_19885_, _19884_, _02851_);
  and (_19886_, _19885_, _19881_);
  and (_19887_, _17563_, _04724_);
  or (_19888_, _19887_, _19831_);
  and (_19889_, _19888_, _02576_);
  or (_19890_, _19889_, _03014_);
  or (_19891_, _19890_, _19886_);
  and (_19892_, _11758_, _04724_);
  or (_19893_, _19892_, _19831_);
  or (_19894_, _19893_, _03884_);
  and (_19895_, _19894_, _19891_);
  or (_19896_, _19895_, _03021_);
  and (_19897_, _11646_, _04724_);
  or (_19898_, _19831_, _05279_);
  or (_19899_, _19898_, _19897_);
  and (_19900_, _19899_, _03131_);
  and (_19902_, _19900_, _19896_);
  or (_19903_, _19902_, _19834_);
  and (_19904_, _19903_, _05274_);
  or (_19905_, _19831_, _04838_);
  and (_19906_, _19893_, _03020_);
  and (_19907_, _19906_, _19905_);
  or (_19908_, _19907_, _19904_);
  and (_19909_, _19908_, _03140_);
  and (_19910_, _19840_, _03139_);
  and (_19911_, _19910_, _19905_);
  or (_19913_, _19911_, _03036_);
  or (_19914_, _19913_, _19909_);
  nor (_19915_, _11644_, _08745_);
  or (_19916_, _19831_, _05781_);
  or (_19917_, _19916_, _19915_);
  and (_19918_, _19917_, _05786_);
  and (_19919_, _19918_, _19914_);
  nor (_19920_, _11768_, _08745_);
  or (_19921_, _19920_, _19831_);
  and (_19922_, _19921_, _03127_);
  or (_19924_, _19922_, _03166_);
  or (_19925_, _19924_, _19919_);
  or (_19926_, _19836_, _03563_);
  and (_19927_, _19926_, _02501_);
  and (_19928_, _19927_, _19925_);
  and (_19929_, _19863_, _02500_);
  or (_19930_, _19929_, _03174_);
  or (_19931_, _19930_, _19928_);
  and (_19932_, _11821_, _04724_);
  or (_19933_, _19831_, _03178_);
  or (_19934_, _19933_, _19932_);
  and (_19935_, _19934_, _34698_);
  and (_19936_, _19935_, _19931_);
  or (_35236_, _19936_, _19830_);
  nor (_19937_, _03006_, _02526_);
  not (_19938_, _19937_);
  and (_19939_, _19938_, _03492_);
  and (_19940_, _09758_, _09765_);
  nor (_19941_, _19940_, _02247_);
  and (_19942_, _09736_, _09743_);
  nor (_19944_, _19942_, _02247_);
  and (_19945_, _08858_, _08136_);
  nor (_19946_, _19945_, _02247_);
  and (_19947_, _07320_, \oc8051_golden_model_1.PC [0]);
  nor (_19948_, _07320_, \oc8051_golden_model_1.PC [0]);
  nor (_19949_, _19948_, _19947_);
  and (_19950_, _19949_, _08864_);
  not (_19951_, _02538_);
  and (_19952_, _08873_, _05781_);
  nor (_19953_, _19952_, _02247_);
  not (_19955_, _02533_);
  and (_19956_, _09473_, _05274_);
  nor (_19957_, _19956_, _02247_);
  and (_19958_, _09448_, _05279_);
  nor (_19959_, _19958_, _02247_);
  and (_19960_, _03014_, _02247_);
  nor (_19961_, _03492_, _02566_);
  and (_19962_, _09169_, _02247_);
  and (_19963_, _03492_, \oc8051_golden_model_1.PC [0]);
  nor (_19964_, _19963_, _09084_);
  not (_19965_, _19964_);
  nor (_19966_, _19965_, _09169_);
  or (_19967_, _19966_, _09172_);
  nor (_19968_, _19967_, _19962_);
  nor (_19969_, _03492_, _02568_);
  and (_19970_, _09247_, _09239_);
  nor (_19971_, _19970_, _02247_);
  and (_19972_, _02563_, _02558_);
  or (_19973_, _19972_, _03492_);
  and (_19974_, _09203_, _09202_);
  nor (_19976_, _19974_, _02247_);
  or (_19977_, _19976_, _09224_);
  nor (_19978_, _09207_, _02247_);
  and (_19979_, _09207_, _02247_);
  nor (_19980_, _19979_, _19978_);
  and (_19981_, _19980_, _02558_);
  not (_19982_, _19981_);
  and (_19983_, _19982_, _19974_);
  or (_19984_, _19983_, _19977_);
  and (_19985_, _19984_, _05387_);
  and (_19987_, _19985_, _19973_);
  and (_19988_, _09196_, \oc8051_golden_model_1.PC [0]);
  and (_19989_, _02832_, _02247_);
  nor (_19990_, _19989_, _08943_);
  and (_19991_, _19990_, _09198_);
  or (_19992_, _19991_, _19988_);
  nor (_19993_, _19992_, _05387_);
  nor (_19994_, _19993_, _19987_);
  nor (_19995_, _19994_, _03818_);
  and (_19996_, _03818_, \oc8051_golden_model_1.PC [0]);
  nor (_19998_, _19996_, _02952_);
  not (_19999_, _19998_);
  nor (_20000_, _19999_, _19995_);
  not (_20001_, _20000_);
  and (_20002_, _19965_, _09186_);
  nor (_20003_, _09186_, _02247_);
  or (_20004_, _20003_, _03821_);
  or (_20005_, _20004_, _20002_);
  and (_20006_, _20005_, _09180_);
  and (_20007_, _20006_, _20001_);
  nor (_20008_, _09180_, _02247_);
  nor (_20009_, _20008_, _05382_);
  not (_20010_, _20009_);
  nor (_20011_, _20010_, _20007_);
  nor (_20012_, _03492_, _02556_);
  not (_20013_, _19970_);
  nor (_20014_, _20013_, _20012_);
  not (_20015_, _20014_);
  nor (_20016_, _20015_, _20011_);
  or (_20017_, _20016_, _09251_);
  nor (_20019_, _20017_, _19971_);
  nor (_20020_, _20019_, _19969_);
  or (_20021_, _20020_, _09299_);
  and (_20022_, _09297_, \oc8051_golden_model_1.PC [0]);
  nor (_20023_, _19964_, _09297_);
  or (_20024_, _20023_, _09263_);
  or (_20025_, _20024_, _20022_);
  and (_20026_, _20025_, _09172_);
  and (_20027_, _20026_, _20021_);
  nor (_20028_, _20027_, _02966_);
  not (_20030_, _20028_);
  nor (_20031_, _20030_, _19968_);
  and (_20032_, _09334_, _02247_);
  nor (_20033_, _19965_, _09334_);
  nor (_20034_, _20033_, _20032_);
  nor (_20035_, _20034_, _03377_);
  nor (_20036_, _20035_, _20031_);
  nor (_20037_, _20036_, _03025_);
  nor (_20038_, _19964_, _09325_);
  and (_20039_, _09325_, \oc8051_golden_model_1.PC [0]);
  or (_20040_, _20039_, _10029_);
  nor (_20041_, _20040_, _20038_);
  or (_20042_, _20041_, _20037_);
  and (_20043_, _20042_, _09306_);
  and (_20044_, _09305_, _02247_);
  or (_20045_, _20044_, _20043_);
  and (_20046_, _20045_, _02561_);
  not (_20047_, _09012_);
  nor (_20048_, _03492_, _02561_);
  nor (_20049_, _20048_, _20047_);
  not (_20051_, _20049_);
  nor (_20052_, _20051_, _20046_);
  nor (_20053_, _09012_, _02247_);
  nor (_20054_, _20053_, _09347_);
  not (_20055_, _20054_);
  nor (_20056_, _20055_, _20052_);
  and (_20057_, _09005_, _02586_);
  not (_20058_, _20057_);
  or (_20059_, _20058_, _20056_);
  nor (_20060_, _20059_, _19961_);
  nor (_20062_, _20057_, _02247_);
  nor (_20063_, _20062_, _02578_);
  not (_20064_, _20063_);
  nor (_20065_, _20064_, _20060_);
  nor (_20066_, _03492_, _05325_);
  nor (_20067_, _03023_, _02576_);
  and (_20068_, _20067_, _09376_);
  not (_20069_, _20068_);
  nor (_20070_, _20069_, _20066_);
  not (_20071_, _20070_);
  nor (_20073_, _20071_, _20065_);
  nor (_20074_, _20068_, _02247_);
  nor (_20075_, _20074_, _02521_);
  not (_20076_, _20075_);
  nor (_20077_, _20076_, _20073_);
  not (_20078_, _02521_);
  nor (_20079_, _03492_, _20078_);
  or (_20080_, _20079_, _09384_);
  nor (_20081_, _20080_, _20077_);
  nor (_20082_, _19990_, _09385_);
  nor (_20084_, _20082_, _20081_);
  and (_20085_, _20084_, _03884_);
  or (_20086_, _20085_, _19960_);
  and (_20087_, _20086_, _09401_);
  and (_20088_, _09400_, _02591_);
  or (_20089_, _20088_, _20087_);
  and (_20090_, _20089_, _04123_);
  nor (_20091_, _03492_, _04123_);
  or (_20092_, _20091_, _20090_);
  and (_20093_, _20092_, _09442_);
  not (_20095_, _19958_);
  and (_20096_, _08190_, \oc8051_golden_model_1.PC [0]);
  and (_20097_, _19990_, _08880_);
  or (_20098_, _20097_, _20096_);
  and (_20099_, _20098_, _09000_);
  nor (_20100_, _20099_, _20095_);
  not (_20101_, _20100_);
  nor (_20102_, _20101_, _20093_);
  nor (_20103_, _20102_, _19959_);
  and (_20104_, _20103_, _02513_);
  nor (_20106_, _03492_, _02513_);
  or (_20107_, _20106_, _20104_);
  and (_20108_, _20107_, _09462_);
  not (_20109_, _19956_);
  nor (_20110_, _19990_, _08880_);
  nor (_20111_, _08190_, \oc8051_golden_model_1.PC [0]);
  nor (_20112_, _20111_, _09462_);
  not (_20113_, _20112_);
  nor (_20114_, _20113_, _20110_);
  nor (_20115_, _20114_, _20109_);
  not (_20117_, _20115_);
  nor (_20118_, _20117_, _20108_);
  nor (_20119_, _20118_, _19957_);
  and (_20120_, _20119_, _19955_);
  nor (_20121_, _03492_, _19955_);
  or (_20122_, _20121_, _20120_);
  and (_20123_, _20122_, _08876_);
  not (_20124_, _19952_);
  and (_20125_, _07325_, \oc8051_golden_model_1.PC [0]);
  nor (_20126_, _07325_, \oc8051_golden_model_1.PC [0]);
  nor (_20128_, _20126_, _20125_);
  and (_20129_, _20128_, _08875_);
  nor (_20130_, _20129_, _20124_);
  not (_20131_, _20130_);
  nor (_20132_, _20131_, _20123_);
  nor (_20133_, _20132_, _19953_);
  and (_20134_, _20133_, _19951_);
  nor (_20135_, _03492_, _19951_);
  or (_20136_, _20135_, _20134_);
  and (_20137_, _20136_, _08865_);
  and (_20139_, _08862_, _08030_);
  not (_20140_, _20139_);
  or (_20141_, _20140_, _20137_);
  nor (_20142_, _20141_, _19950_);
  nor (_20143_, _20139_, _02247_);
  nor (_20144_, _20143_, _03148_);
  not (_20145_, _20144_);
  nor (_20146_, _20145_, _20142_);
  and (_20147_, _06174_, _03148_);
  or (_20148_, _20147_, _20146_);
  and (_20149_, _20148_, _05792_);
  nor (_20150_, _03492_, _05792_);
  or (_20151_, _20150_, _20149_);
  and (_20152_, _20151_, _03152_);
  and (_20153_, _19965_, _09709_);
  nor (_20154_, _09709_, _02247_);
  or (_20155_, _20154_, _03152_);
  or (_20156_, _20155_, _20153_);
  and (_20157_, _20156_, _19945_);
  not (_20158_, _20157_);
  nor (_20159_, _20158_, _20152_);
  nor (_20160_, _20159_, _19946_);
  and (_20161_, _20160_, _02898_);
  and (_20162_, _06174_, _02897_);
  or (_20163_, _20162_, _20161_);
  and (_20164_, _20163_, _09728_);
  nor (_20165_, _03492_, _09728_);
  nor (_20166_, _20165_, _20164_);
  nor (_20167_, _20166_, _02895_);
  not (_20168_, _19942_);
  and (_20170_, _09709_, \oc8051_golden_model_1.PC [0]);
  nor (_20171_, _19964_, _09709_);
  nor (_20172_, _20171_, _20170_);
  and (_20173_, _20172_, _02895_);
  nor (_20174_, _20173_, _20168_);
  not (_20175_, _20174_);
  nor (_20176_, _20175_, _20167_);
  nor (_20177_, _20176_, _19944_);
  nor (_20178_, _20177_, _04159_);
  and (_20179_, _04159_, _03492_);
  nor (_20181_, _20179_, _02500_);
  not (_20182_, _20181_);
  nor (_20183_, _20182_, _20178_);
  not (_20184_, _19940_);
  and (_20185_, _20172_, _02500_);
  nor (_20186_, _20185_, _20184_);
  not (_20187_, _20186_);
  nor (_20188_, _20187_, _20183_);
  nor (_20189_, _20188_, _19941_);
  nor (_20190_, _20189_, _19938_);
  or (_20192_, _20190_, _09777_);
  nor (_20193_, _20192_, _19939_);
  and (_20194_, _09777_, _02247_);
  nor (_20195_, _20194_, _20193_);
  nand (_20196_, _20195_, _34698_);
  or (_20197_, _34698_, \oc8051_golden_model_1.PC [0]);
  and (_20198_, _20197_, _36029_);
  and (_35239_, _20198_, _20196_);
  nor (_20199_, _09765_, _09082_);
  nor (_20200_, _03381_, _04141_);
  and (_20202_, _09709_, _09082_);
  nor (_20203_, _09086_, _09084_);
  nor (_20204_, _20203_, _09087_);
  nor (_20205_, _20204_, _09709_);
  nor (_20206_, _20205_, _20202_);
  and (_20207_, _20206_, _02500_);
  nor (_20208_, _09743_, _09082_);
  nor (_20209_, _05270_, _09082_);
  nor (_20210_, _08858_, _09082_);
  nor (_20211_, _08862_, _09082_);
  nor (_20213_, _08873_, _09082_);
  nor (_20214_, _09473_, _09082_);
  nor (_20215_, _09450_, _02218_);
  and (_20216_, _07791_, _02602_);
  nor (_20217_, _10050_, _09082_);
  and (_20218_, _09305_, _02602_);
  and (_20219_, _09297_, _02602_);
  not (_20220_, _20204_);
  nor (_20221_, _20220_, _09297_);
  or (_20222_, _20221_, _20219_);
  nor (_20224_, _20222_, _09263_);
  and (_20225_, _03705_, _09251_);
  or (_20226_, _20225_, _02886_);
  nor (_20227_, _03705_, _02563_);
  and (_20228_, _03382_, _02602_);
  nor (_20229_, _19978_, _03825_);
  and (_20230_, _20229_, _02218_);
  nor (_20231_, _20229_, _02218_);
  nor (_20232_, _20231_, _20230_);
  and (_20233_, _20232_, _02558_);
  nor (_20235_, _03705_, _02558_);
  and (_20236_, _02864_, _02953_);
  not (_20237_, _20236_);
  nor (_20238_, _03712_, _03325_);
  and (_20239_, _20238_, _20237_);
  not (_20240_, _20239_);
  or (_20241_, _20240_, _20235_);
  nor (_20242_, _20241_, _20233_);
  nor (_20243_, _20239_, _09082_);
  nor (_20244_, _20243_, _20242_);
  nor (_20246_, _20244_, _03382_);
  or (_20247_, _20246_, _02954_);
  nor (_20248_, _20247_, _20228_);
  and (_20249_, _02954_, _02218_);
  or (_20250_, _20249_, _20248_);
  and (_20251_, _20250_, _09202_);
  and (_20252_, _07452_, _09082_);
  or (_20253_, _20252_, _20251_);
  and (_20254_, _20253_, _02563_);
  or (_20255_, _20254_, _10433_);
  nor (_20257_, _20255_, _20227_);
  or (_20258_, _09198_, _02218_);
  nor (_20259_, _08945_, _08943_);
  nor (_20260_, _20259_, _08946_);
  or (_20261_, _20260_, _09196_);
  nand (_20262_, _20261_, _20258_);
  and (_20263_, _20262_, _10433_);
  or (_20264_, _20263_, _20257_);
  nand (_20265_, _20264_, _05402_);
  and (_20266_, _03818_, _02602_);
  nor (_20268_, _20266_, _02952_);
  and (_20269_, _20268_, _20265_);
  nand (_20270_, _20220_, _09186_);
  or (_20271_, _09186_, _02602_);
  and (_20272_, _20271_, _20270_);
  and (_20273_, _20272_, _02952_);
  nor (_20274_, _20273_, _20269_);
  nand (_20275_, _20274_, _09180_);
  nor (_20276_, _09180_, _09082_);
  nor (_20277_, _20276_, _02891_);
  nand (_20279_, _20277_, _20275_);
  and (_20280_, _02891_, _02218_);
  nor (_20281_, _20280_, _05382_);
  nand (_20282_, _20281_, _20279_);
  and (_20283_, _03705_, _05382_);
  nor (_20284_, _20283_, _02947_);
  nand (_20285_, _20284_, _20282_);
  and (_20286_, _02947_, _02218_);
  nor (_20287_, _20286_, _09240_);
  nand (_20288_, _20287_, _20285_);
  nor (_20290_, _09239_, _09082_);
  nor (_20291_, _20290_, _02950_);
  nand (_20292_, _20291_, _20288_);
  and (_20293_, _02950_, _02218_);
  nor (_20294_, _20293_, _09249_);
  nand (_20295_, _20294_, _20292_);
  nor (_20296_, _09247_, _09082_);
  nor (_20297_, _20296_, _02887_);
  nand (_20298_, _20297_, _20295_);
  and (_20299_, _02887_, _02218_);
  nor (_20301_, _20299_, _09251_);
  and (_20302_, _20301_, _20298_);
  or (_20303_, _20302_, _20226_);
  and (_20304_, _02886_, _02218_);
  nor (_20305_, _20304_, _09299_);
  and (_20306_, _20305_, _20303_);
  or (_20307_, _20306_, _20224_);
  and (_20308_, _20307_, _09172_);
  nor (_20309_, _20220_, _09169_);
  and (_20310_, _09169_, _02602_);
  or (_20312_, _20310_, _20309_);
  nor (_20313_, _20312_, _09172_);
  or (_20314_, _20313_, _20308_);
  or (_20315_, _20314_, _02966_);
  nor (_20316_, _20220_, _09334_);
  and (_20317_, _09334_, _02602_);
  nor (_20318_, _20317_, _20316_);
  or (_20319_, _20318_, _03377_);
  and (_20320_, _20319_, _20315_);
  or (_20321_, _20320_, _03025_);
  nor (_20323_, _20204_, _09325_);
  and (_20324_, _09325_, _09082_);
  or (_20325_, _20324_, _10029_);
  or (_20326_, _20325_, _20323_);
  and (_20327_, _20326_, _09306_);
  and (_20328_, _20327_, _20321_);
  or (_20329_, _20328_, _20218_);
  nand (_20330_, _20329_, _02881_);
  and (_20331_, _02880_, \oc8051_golden_model_1.PC [1]);
  nor (_20332_, _20331_, _04125_);
  nand (_20334_, _20332_, _20330_);
  nor (_20335_, _03705_, _02561_);
  nor (_20336_, _03867_, _02942_);
  and (_20337_, _20336_, _04118_);
  and (_20338_, _02843_, _02980_);
  nor (_20339_, _20338_, _02978_);
  and (_20340_, _20339_, _20337_);
  not (_20341_, _20340_);
  nor (_20342_, _20341_, _20335_);
  nand (_20343_, _20342_, _20334_);
  nor (_20345_, _20340_, _02218_);
  nor (_20346_, _20345_, _09009_);
  nand (_20347_, _20346_, _20343_);
  and (_20348_, _09011_, _02602_);
  or (_20349_, _20348_, _09012_);
  nand (_20350_, _20349_, _20347_);
  nor (_20351_, _09011_, _09082_);
  nor (_20352_, _20351_, _02987_);
  nand (_20353_, _20352_, _20350_);
  and (_20354_, _02987_, _02218_);
  nor (_20356_, _20354_, _09347_);
  nand (_20357_, _20356_, _20353_);
  and (_20358_, _03705_, _09347_);
  nor (_20359_, _20358_, _02986_);
  nand (_20360_, _20359_, _20357_);
  and (_20361_, _02986_, _02218_);
  not (_20362_, _20361_);
  and (_20363_, _20362_, _10050_);
  and (_20364_, _20363_, _20360_);
  or (_20365_, _20364_, _20217_);
  and (_20367_, _14648_, _02577_);
  not (_20368_, _20367_);
  and (_20369_, _20368_, _07424_);
  nand (_20370_, _20369_, _20365_);
  nor (_20371_, _20369_, _09082_);
  nor (_20372_, _20371_, _03442_);
  nand (_20373_, _20372_, _20370_);
  and (_20374_, _03442_, _09082_);
  nor (_20375_, _20374_, _07597_);
  nand (_20376_, _20375_, _20373_);
  nor (_20378_, _07596_, _02218_);
  nor (_20379_, _20378_, _02585_);
  and (_20380_, _20379_, _20376_);
  and (_20381_, _09082_, _02585_);
  or (_20382_, _20381_, _02874_);
  nor (_20383_, _20382_, _20380_);
  and (_20384_, _02874_, \oc8051_golden_model_1.PC [1]);
  or (_20385_, _20384_, _20383_);
  nand (_20386_, _20385_, _05325_);
  and (_20387_, _03705_, _02578_);
  nor (_20389_, _20387_, _03023_);
  nand (_20390_, _20389_, _20386_);
  not (_20391_, _09369_);
  and (_20392_, _03023_, _02602_);
  nor (_20393_, _20392_, _20391_);
  nand (_20394_, _20393_, _20390_);
  nor (_20395_, _09369_, _02218_);
  nor (_20396_, _20395_, _02576_);
  nand (_20397_, _20396_, _20394_);
  and (_20398_, _02602_, _02576_);
  nor (_20400_, _20398_, _09378_);
  nand (_20401_, _20400_, _20397_);
  nor (_20402_, _09376_, _09082_);
  nor (_20403_, _20402_, _02938_);
  nand (_20404_, _20403_, _20401_);
  and (_20405_, _02938_, _02218_);
  nor (_20406_, _20405_, _02521_);
  nand (_20407_, _20406_, _20404_);
  and (_20408_, _03705_, _02521_);
  nor (_20409_, _20408_, _09384_);
  nand (_20411_, _20409_, _20407_);
  and (_20412_, _20260_, _09384_);
  nor (_20413_, _20412_, _05562_);
  nand (_20414_, _20413_, _20411_);
  nor (_20415_, _05322_, _02218_);
  nor (_20416_, _20415_, _03014_);
  nand (_20417_, _20416_, _20414_);
  and (_20418_, _03014_, _02602_);
  nor (_20419_, _20418_, _07782_);
  and (_20420_, _20419_, _20417_);
  and (_20422_, _07782_, \oc8051_golden_model_1.PC [1]);
  or (_20423_, _20422_, _20420_);
  nand (_20424_, _20423_, _09401_);
  nor (_20425_, _09401_, _02611_);
  nor (_20426_, _20425_, _02937_);
  nand (_20427_, _20426_, _20424_);
  and (_20428_, _02937_, _02218_);
  nor (_20429_, _20428_, _02517_);
  nand (_20430_, _20429_, _20427_);
  and (_20431_, _03705_, _02517_);
  nor (_20433_, _20431_, _09000_);
  nand (_20434_, _20433_, _20430_);
  and (_20435_, _08190_, _02218_);
  and (_20436_, _20260_, _08880_);
  or (_20437_, _20436_, _20435_);
  and (_20438_, _20437_, _09000_);
  nor (_20439_, _20438_, _07791_);
  and (_20440_, _20439_, _20434_);
  or (_20441_, _20440_, _20216_);
  and (_20442_, _07802_, _02545_);
  not (_20444_, _20442_);
  and (_20445_, _20444_, _07797_);
  nand (_20446_, _20445_, _20441_);
  nor (_20447_, _20445_, _09082_);
  nor (_20448_, _20447_, _03504_);
  nand (_20449_, _20448_, _20446_);
  and (_20450_, _03504_, _09082_);
  nor (_20451_, _20450_, _09451_);
  and (_20452_, _20451_, _20449_);
  or (_20453_, _20452_, _20215_);
  nand (_20455_, _20453_, _05279_);
  and (_20456_, _03021_, _09082_);
  nor (_20457_, _20456_, _03130_);
  nand (_20458_, _20457_, _20455_);
  and (_20459_, _03130_, _02218_);
  nor (_20460_, _20459_, _02512_);
  nand (_20461_, _20460_, _20458_);
  and (_20462_, _03705_, _02512_);
  nor (_20463_, _20462_, _08994_);
  nand (_20464_, _20463_, _20461_);
  not (_20466_, _09473_);
  nor (_20467_, _20260_, _08880_);
  nor (_20468_, _08190_, _02218_);
  nor (_20469_, _20468_, _09462_);
  not (_20470_, _20469_);
  nor (_20471_, _20470_, _20467_);
  nor (_20472_, _20471_, _20466_);
  and (_20473_, _20472_, _20464_);
  or (_20474_, _20473_, _20214_);
  nand (_20475_, _20474_, _09475_);
  nor (_20477_, _09475_, _02218_);
  nor (_20478_, _20477_, _03020_);
  and (_20479_, _20478_, _20475_);
  and (_20480_, _03020_, _02602_);
  or (_20481_, _20480_, _03139_);
  nor (_20482_, _20481_, _20479_);
  and (_20483_, _03139_, \oc8051_golden_model_1.PC [1]);
  or (_20484_, _20483_, _20482_);
  nand (_20485_, _20484_, _19955_);
  and (_20486_, _03705_, _02533_);
  nor (_20488_, _20486_, _08875_);
  nand (_20489_, _20488_, _20485_);
  and (_20490_, \oc8051_golden_model_1.PSW [7], _02218_);
  and (_20491_, _20260_, _07319_);
  or (_20492_, _20491_, _20490_);
  and (_20493_, _20492_, _08875_);
  nor (_20494_, _20493_, _09487_);
  and (_20495_, _20494_, _20489_);
  or (_20496_, _20495_, _20213_);
  nand (_20497_, _20496_, _07866_);
  nor (_20499_, _07866_, _02218_);
  nor (_20500_, _20499_, _03036_);
  and (_20501_, _20500_, _20497_);
  and (_20502_, _03036_, _02602_);
  or (_20503_, _20502_, _03127_);
  nor (_20504_, _20503_, _20501_);
  and (_20505_, _03127_, \oc8051_golden_model_1.PC [1]);
  or (_20506_, _20505_, _20504_);
  nand (_20507_, _20506_, _19951_);
  and (_20508_, _03705_, _02538_);
  nor (_20510_, _20508_, _08864_);
  nand (_20511_, _20510_, _20507_);
  nor (_20512_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_20513_, _20260_, \oc8051_golden_model_1.PSW [7]);
  or (_20514_, _20513_, _20512_);
  and (_20515_, _20514_, _08864_);
  nor (_20516_, _20515_, _09503_);
  and (_20517_, _20516_, _20511_);
  or (_20518_, _20517_, _20211_);
  nand (_20519_, _20518_, _08860_);
  nor (_20521_, _08860_, _02218_);
  nor (_20522_, _20521_, _08029_);
  nand (_20523_, _20522_, _20519_);
  and (_20524_, _08029_, _09082_);
  nor (_20525_, _20524_, _03148_);
  and (_20526_, _20525_, _20523_);
  and (_20527_, _05893_, _03148_);
  or (_20528_, _20527_, _20526_);
  nand (_20529_, _20528_, _05792_);
  and (_20530_, _03705_, _02531_);
  nor (_20532_, _20530_, _03035_);
  nand (_20533_, _20532_, _20529_);
  nor (_20534_, _09709_, _02602_);
  not (_20535_, _20534_);
  and (_20536_, _20220_, _09709_);
  nor (_20537_, _20536_, _03152_);
  and (_20538_, _20537_, _20535_);
  nor (_20539_, _20538_, _09524_);
  and (_20540_, _20539_, _20533_);
  or (_20541_, _20540_, _20210_);
  nand (_20543_, _20541_, _08104_);
  nor (_20544_, _08104_, _02218_);
  nor (_20545_, _20544_, _08135_);
  and (_20546_, _20545_, _20543_);
  and (_20547_, _08135_, _09082_);
  or (_20548_, _20547_, _02897_);
  nor (_20549_, _20548_, _20546_);
  and (_20550_, _05893_, _02897_);
  or (_20551_, _20550_, _20549_);
  nand (_20552_, _20551_, _09728_);
  and (_20554_, _03705_, _02536_);
  nor (_20555_, _20554_, _02895_);
  nand (_20556_, _20555_, _20552_);
  and (_20557_, _20206_, _02895_);
  nor (_20558_, _20557_, _11177_);
  and (_20559_, _20558_, _20556_);
  or (_20560_, _20559_, _20209_);
  and (_20561_, _04084_, _03910_);
  nand (_20562_, _20561_, _20560_);
  nor (_20563_, _20561_, _09082_);
  nor (_20565_, _20563_, _03166_);
  nand (_20566_, _20565_, _20562_);
  and (_20567_, _03166_, _02218_);
  nor (_20568_, _20567_, _09744_);
  and (_20569_, _20568_, _20566_);
  or (_20570_, _20569_, _20208_);
  nand (_20571_, _20570_, _03916_);
  and (_20572_, _04159_, _03705_);
  nor (_20573_, _20572_, _02500_);
  and (_20574_, _20573_, _20571_);
  nor (_20576_, _20574_, _20207_);
  and (_20577_, _20576_, _10792_);
  nor (_20578_, _10792_, _09082_);
  nor (_20579_, _20578_, _20577_);
  or (_20580_, _20579_, _20200_);
  and (_20581_, _20200_, _02602_);
  nor (_20582_, _20581_, _03174_);
  nand (_20583_, _20582_, _20580_);
  and (_20584_, _03174_, _02218_);
  nor (_20585_, _20584_, _09766_);
  and (_20587_, _20585_, _20583_);
  or (_20588_, _20587_, _20199_);
  nand (_20589_, _20588_, _19937_);
  and (_20590_, _19938_, _03705_);
  nor (_20591_, _20590_, _09777_);
  and (_20592_, _20591_, _20589_);
  and (_20593_, _09777_, _09082_);
  or (_20594_, _20593_, _20592_);
  or (_20595_, _20594_, _34702_);
  or (_20596_, _34698_, \oc8051_golden_model_1.PC [1]);
  and (_20598_, _20596_, _36029_);
  and (_35240_, _20598_, _20595_);
  and (_20599_, _03174_, _02633_);
  and (_20600_, _03166_, _02633_);
  nor (_20601_, _08858_, _02638_);
  nor (_20602_, _08862_, _02638_);
  nor (_20603_, _08873_, _02638_);
  nor (_20604_, _09473_, _02638_);
  nor (_20605_, _09448_, _02638_);
  nor (_20606_, _06241_, _02633_);
  and (_20608_, _02874_, _02634_);
  nor (_20609_, _20340_, _02633_);
  and (_20610_, _09305_, _03054_);
  and (_20611_, _09091_, _09088_);
  nor (_20612_, _20611_, _09092_);
  nor (_20613_, _20612_, _09169_);
  and (_20614_, _09169_, _09080_);
  nor (_20615_, _20614_, _20613_);
  nor (_20616_, _20615_, _09172_);
  and (_20617_, _09196_, _02633_);
  and (_20619_, _08950_, _08947_);
  nor (_20620_, _20619_, _08951_);
  and (_20621_, _20620_, _09198_);
  nor (_20622_, _20621_, _20617_);
  and (_20623_, _20622_, _10433_);
  and (_20624_, _09206_, _02223_);
  nor (_20625_, _20624_, _03825_);
  and (_20626_, _03825_, _02633_);
  nor (_20627_, _20626_, _07442_);
  not (_20628_, _20627_);
  nor (_20630_, _20628_, _20625_);
  not (_20631_, _20630_);
  nor (_20632_, _09207_, _02638_);
  nor (_20633_, _20632_, _03824_);
  and (_20634_, _20633_, _20631_);
  not (_20635_, _09203_);
  nor (_20636_, _03302_, _02558_);
  or (_20637_, _20636_, _20635_);
  nor (_20638_, _20637_, _20634_);
  nor (_20639_, _09203_, _02638_);
  nor (_20641_, _20639_, _02954_);
  not (_20642_, _20641_);
  nor (_20643_, _20642_, _20638_);
  and (_20644_, _02954_, _02633_);
  or (_20645_, _20644_, _20643_);
  and (_20646_, _20645_, _09202_);
  and (_20647_, _07452_, _02638_);
  or (_20648_, _20647_, _20646_);
  and (_20649_, _20648_, _02563_);
  nor (_20650_, _03302_, _02563_);
  nor (_20652_, _20650_, _10433_);
  not (_20653_, _20652_);
  nor (_20654_, _20653_, _20649_);
  or (_20655_, _20654_, _20623_);
  nand (_20656_, _20655_, _05402_);
  and (_20657_, _03818_, _03054_);
  nor (_20658_, _20657_, _02952_);
  and (_20659_, _20658_, _20656_);
  not (_20660_, _20612_);
  nand (_20661_, _20660_, _09186_);
  or (_20663_, _09186_, _09079_);
  and (_20664_, _20663_, _20661_);
  and (_20665_, _20664_, _02952_);
  nor (_20666_, _20665_, _20659_);
  nand (_20667_, _20666_, _09180_);
  nor (_20668_, _09180_, _02638_);
  nor (_20669_, _20668_, _02891_);
  nand (_20670_, _20669_, _20667_);
  and (_20671_, _02891_, _02633_);
  nor (_20672_, _20671_, _05382_);
  nand (_20674_, _20672_, _20670_);
  and (_20675_, _03302_, _05382_);
  nor (_20676_, _20675_, _02947_);
  nand (_20677_, _20676_, _20674_);
  and (_20678_, _02947_, _02633_);
  nor (_20679_, _20678_, _09240_);
  nand (_20680_, _20679_, _20677_);
  nor (_20681_, _09239_, _02638_);
  nor (_20682_, _20681_, _02950_);
  nand (_20683_, _20682_, _20680_);
  and (_20685_, _02950_, _02633_);
  nor (_20686_, _20685_, _09249_);
  nand (_20687_, _20686_, _20683_);
  nor (_20688_, _09247_, _02638_);
  nor (_20689_, _20688_, _02887_);
  nand (_20690_, _20689_, _20687_);
  and (_20691_, _02887_, _02633_);
  nor (_20692_, _20691_, _09251_);
  nand (_20693_, _20692_, _20690_);
  and (_20694_, _03302_, _09251_);
  nor (_20696_, _20694_, _02886_);
  nand (_20697_, _20696_, _20693_);
  and (_20698_, _02886_, _02633_);
  nor (_20699_, _20698_, _09299_);
  and (_20700_, _20699_, _20697_);
  nor (_20701_, _20612_, _09297_);
  and (_20702_, _09297_, _09080_);
  nor (_20703_, _20702_, _20701_);
  nor (_20704_, _20703_, _09263_);
  or (_20705_, _20704_, _20700_);
  and (_20707_, _20705_, _09172_);
  or (_20708_, _20707_, _20616_);
  or (_20709_, _20708_, _02966_);
  and (_20710_, _09334_, _09079_);
  nor (_20711_, _20660_, _09334_);
  nor (_20712_, _20711_, _20710_);
  or (_20713_, _20712_, _03377_);
  and (_20714_, _20713_, _20709_);
  or (_20715_, _20714_, _03025_);
  nor (_20716_, _20612_, _09325_);
  and (_20718_, _09325_, _09080_);
  or (_20719_, _20718_, _10029_);
  or (_20720_, _20719_, _20716_);
  and (_20721_, _20720_, _09306_);
  and (_20722_, _20721_, _20715_);
  or (_20723_, _20722_, _20610_);
  nand (_20724_, _20723_, _02881_);
  and (_20725_, _02880_, _02634_);
  nor (_20726_, _20725_, _04125_);
  nand (_20727_, _20726_, _20724_);
  nor (_20729_, _03302_, _02561_);
  nor (_20730_, _20729_, _20341_);
  and (_20731_, _20730_, _20727_);
  or (_20732_, _20731_, _20609_);
  nand (_20733_, _20732_, _09012_);
  nor (_20734_, _09012_, _02638_);
  nor (_20735_, _20734_, _02987_);
  nand (_20736_, _20735_, _20733_);
  and (_20737_, _02987_, _02633_);
  nor (_20738_, _20737_, _09347_);
  nand (_20740_, _20738_, _20736_);
  and (_20741_, _03302_, _09347_);
  nor (_20742_, _20741_, _02986_);
  nand (_20743_, _20742_, _20740_);
  and (_20744_, _02986_, _02633_);
  nor (_20745_, _20744_, _13666_);
  and (_20746_, _20745_, _20743_);
  nor (_20747_, _09005_, _02638_);
  or (_20748_, _20747_, _20746_);
  nand (_20749_, _20748_, _07596_);
  nor (_20751_, _07596_, _02633_);
  nor (_20752_, _20751_, _02585_);
  nand (_20753_, _20752_, _20749_);
  and (_20754_, _02638_, _02585_);
  nor (_20755_, _20754_, _02874_);
  and (_20756_, _20755_, _20753_);
  or (_20757_, _20756_, _20608_);
  nand (_20758_, _20757_, _05325_);
  and (_20759_, _03302_, _02578_);
  nor (_20760_, _20759_, _03023_);
  nand (_20762_, _20760_, _20758_);
  and (_20763_, _09079_, _03023_);
  nor (_20764_, _20763_, _06793_);
  and (_20765_, _20764_, _20762_);
  or (_20766_, _20765_, _20606_);
  nand (_20767_, _20766_, _02856_);
  and (_20768_, _02855_, _02634_);
  nor (_20769_, _20768_, _02576_);
  nand (_20770_, _20769_, _20767_);
  and (_20771_, _09079_, _02576_);
  nor (_20773_, _20771_, _09378_);
  nand (_20774_, _20773_, _20770_);
  nor (_20775_, _09376_, _02638_);
  nor (_20776_, _20775_, _02938_);
  nand (_20777_, _20776_, _20774_);
  and (_20778_, _02938_, _02633_);
  nor (_20779_, _20778_, _02521_);
  and (_20780_, _20779_, _20777_);
  and (_20781_, _03302_, _02521_);
  or (_20782_, _20781_, _20780_);
  nand (_20784_, _20782_, _09385_);
  nor (_20785_, _20620_, _09385_);
  nor (_20786_, _20785_, _05562_);
  and (_20787_, _20786_, _20784_);
  nor (_20788_, _05322_, _02634_);
  or (_20789_, _20788_, _03014_);
  or (_20790_, _20789_, _20787_);
  and (_20791_, _09080_, _03014_);
  nor (_20792_, _20791_, _07782_);
  nand (_20793_, _20792_, _20790_);
  and (_20795_, _07782_, _02633_);
  nor (_20796_, _20795_, _09400_);
  nand (_20797_, _20796_, _20793_);
  and (_20798_, _09400_, _02649_);
  nor (_20799_, _20798_, _02937_);
  nand (_20800_, _20799_, _20797_);
  and (_20801_, _02937_, _02633_);
  nor (_20802_, _20801_, _02517_);
  nand (_20803_, _20802_, _20800_);
  and (_20804_, _03302_, _02517_);
  nor (_20806_, _20804_, _09000_);
  nand (_20807_, _20806_, _20803_);
  not (_20808_, _09448_);
  and (_20809_, _08190_, _02633_);
  and (_20810_, _20620_, _08880_);
  or (_20811_, _20810_, _20809_);
  and (_20812_, _20811_, _09000_);
  nor (_20813_, _20812_, _20808_);
  and (_20814_, _20813_, _20807_);
  or (_20815_, _20814_, _20605_);
  nand (_20817_, _20815_, _09450_);
  nor (_20818_, _09450_, _02633_);
  nor (_20819_, _20818_, _03021_);
  and (_20820_, _20819_, _20817_);
  and (_20821_, _09079_, _03021_);
  or (_20822_, _20821_, _03130_);
  nor (_20823_, _20822_, _20820_);
  and (_20824_, _03130_, _02634_);
  or (_20825_, _20824_, _20823_);
  nand (_20826_, _20825_, _02513_);
  and (_20828_, _03302_, _02512_);
  nor (_20829_, _20828_, _08994_);
  nand (_20830_, _20829_, _20826_);
  nor (_20831_, _20620_, _08880_);
  nor (_20832_, _08190_, _02633_);
  nor (_20833_, _20832_, _09462_);
  not (_20834_, _20833_);
  nor (_20835_, _20834_, _20831_);
  nor (_20836_, _20835_, _20466_);
  and (_20837_, _20836_, _20830_);
  or (_20839_, _20837_, _20604_);
  nand (_20840_, _20839_, _09475_);
  nor (_20841_, _09475_, _02633_);
  nor (_20842_, _20841_, _03020_);
  and (_20843_, _20842_, _20840_);
  and (_20844_, _09079_, _03020_);
  or (_20845_, _20844_, _03139_);
  nor (_20846_, _20845_, _20843_);
  and (_20847_, _03139_, _02634_);
  or (_20848_, _20847_, _20846_);
  nand (_20850_, _20848_, _19955_);
  and (_20851_, _03302_, _02533_);
  nor (_20852_, _20851_, _08875_);
  nand (_20853_, _20852_, _20850_);
  nor (_20854_, _20620_, \oc8051_golden_model_1.PSW [7]);
  nor (_20855_, _02633_, _07319_);
  nor (_20856_, _20855_, _08876_);
  not (_20857_, _20856_);
  nor (_20858_, _20857_, _20854_);
  nor (_20859_, _20858_, _09487_);
  and (_20861_, _20859_, _20853_);
  or (_20862_, _20861_, _20603_);
  nand (_20863_, _20862_, _07866_);
  nor (_20864_, _07866_, _02633_);
  nor (_20865_, _20864_, _03036_);
  nand (_20866_, _20865_, _20863_);
  and (_20867_, _09079_, _03036_);
  nor (_20868_, _20867_, _03127_);
  and (_20869_, _20868_, _20866_);
  and (_20870_, _03127_, _02634_);
  or (_20872_, _20870_, _20869_);
  nand (_20873_, _20872_, _19951_);
  and (_20874_, _03302_, _02538_);
  nor (_20875_, _20874_, _08864_);
  nand (_20876_, _20875_, _20873_);
  and (_20877_, _02633_, _07319_);
  and (_20878_, _20620_, \oc8051_golden_model_1.PSW [7]);
  or (_20879_, _20878_, _20877_);
  and (_20880_, _20879_, _08864_);
  nor (_20881_, _20880_, _09503_);
  and (_20883_, _20881_, _20876_);
  or (_20884_, _20883_, _20602_);
  nand (_20885_, _20884_, _08860_);
  nor (_20886_, _08860_, _02633_);
  nor (_20887_, _20886_, _08029_);
  and (_20888_, _20887_, _20885_);
  and (_20889_, _08029_, _02638_);
  or (_20890_, _20889_, _03148_);
  nor (_20891_, _20890_, _20888_);
  and (_20892_, _06029_, _03148_);
  or (_20894_, _20892_, _20891_);
  nand (_20895_, _20894_, _05792_);
  and (_20896_, _03302_, _02531_);
  nor (_20897_, _20896_, _03035_);
  nand (_20898_, _20897_, _20895_);
  nor (_20899_, _09709_, _09079_);
  and (_20900_, _20660_, _09709_);
  or (_20901_, _20900_, _03152_);
  or (_20902_, _20901_, _20899_);
  and (_20903_, _20902_, _08858_);
  and (_20905_, _20903_, _20898_);
  or (_20906_, _20905_, _20601_);
  nand (_20907_, _20906_, _08104_);
  nor (_20908_, _08104_, _02633_);
  nor (_20909_, _20908_, _08135_);
  and (_20910_, _20909_, _20907_);
  and (_20911_, _08135_, _02638_);
  or (_20912_, _20911_, _02897_);
  nor (_20913_, _20912_, _20910_);
  and (_20914_, _06029_, _02897_);
  or (_20916_, _20914_, _20913_);
  nand (_20917_, _20916_, _09728_);
  and (_20918_, _03302_, _02536_);
  nor (_20919_, _20918_, _02895_);
  nand (_20920_, _20919_, _20917_);
  nor (_20921_, _20612_, _09709_);
  and (_20922_, _09709_, _09080_);
  nor (_20923_, _20922_, _20921_);
  and (_20924_, _20923_, _02895_);
  nor (_20925_, _20924_, _09737_);
  nand (_20927_, _20925_, _20920_);
  nor (_20928_, _09736_, _02638_);
  nor (_20929_, _20928_, _03166_);
  and (_20930_, _20929_, _20927_);
  or (_20931_, _20930_, _20600_);
  nand (_20932_, _20931_, _09743_);
  nor (_20933_, _09743_, _03054_);
  nor (_20934_, _20933_, _04159_);
  nand (_20935_, _20934_, _20932_);
  and (_20936_, _04159_, _03302_);
  nor (_20938_, _20936_, _02500_);
  nand (_20939_, _20938_, _20935_);
  and (_20940_, _20923_, _02500_);
  nor (_20941_, _20940_, _09759_);
  nand (_20942_, _20941_, _20939_);
  nor (_20943_, _09758_, _02638_);
  nor (_20944_, _20943_, _03174_);
  and (_20945_, _20944_, _20942_);
  or (_20946_, _20945_, _20599_);
  nand (_20947_, _20946_, _09765_);
  nor (_20949_, _09765_, _03054_);
  nor (_20950_, _20949_, _19938_);
  nand (_20951_, _20950_, _20947_);
  and (_20952_, _19938_, _03302_);
  nor (_20953_, _20952_, _09777_);
  and (_20954_, _20953_, _20951_);
  and (_20955_, _09777_, _02638_);
  or (_20956_, _20955_, _20954_);
  or (_20957_, _20956_, _34702_);
  or (_20958_, _34698_, \oc8051_golden_model_1.PC [2]);
  and (_20960_, _20958_, _36029_);
  and (_35241_, _20960_, _20957_);
  and (_20961_, _09777_, _02693_);
  and (_20962_, _03174_, _02676_);
  and (_20963_, _03166_, _02676_);
  nor (_20964_, _08858_, _02693_);
  nor (_20965_, _08862_, _02693_);
  nor (_20966_, _08873_, _02693_);
  nor (_20967_, _09473_, _02693_);
  nor (_20968_, _09448_, _02693_);
  and (_20970_, _07782_, _02677_);
  and (_20971_, _02874_, _02677_);
  and (_20972_, _09305_, _02692_);
  or (_20973_, _09077_, _09076_);
  and (_20974_, _20973_, _09093_);
  nor (_20975_, _20973_, _09093_);
  nor (_20976_, _20975_, _20974_);
  nor (_20977_, _20976_, _09169_);
  and (_20978_, _09169_, _09075_);
  nor (_20979_, _20978_, _20977_);
  nor (_20981_, _20979_, _09172_);
  nor (_20982_, _09186_, _09074_);
  not (_20983_, _20976_);
  and (_20984_, _20983_, _09186_);
  nor (_20985_, _20984_, _20982_);
  nor (_20986_, _20985_, _03821_);
  and (_20987_, _09196_, _02676_);
  or (_20988_, _08940_, _08939_);
  and (_20989_, _20988_, _08952_);
  nor (_20990_, _20988_, _08952_);
  nor (_20992_, _20990_, _20989_);
  and (_20993_, _20992_, _09198_);
  or (_20994_, _20993_, _20987_);
  nor (_20995_, _20994_, _05387_);
  and (_20996_, _09206_, _02214_);
  nor (_20997_, _20996_, _03825_);
  and (_20998_, _03825_, _02676_);
  nor (_20999_, _20998_, _07442_);
  not (_21000_, _20999_);
  nor (_21001_, _21000_, _20997_);
  not (_21003_, _21001_);
  nor (_21004_, _09207_, _02693_);
  nor (_21005_, _21004_, _03824_);
  and (_21006_, _21005_, _21003_);
  nor (_21007_, _03120_, _02558_);
  or (_21008_, _21007_, _20635_);
  nor (_21009_, _21008_, _21006_);
  nor (_21010_, _09203_, _02693_);
  nor (_21011_, _21010_, _02954_);
  not (_21012_, _21011_);
  nor (_21014_, _21012_, _21009_);
  and (_21015_, _02954_, _02676_);
  or (_21016_, _21015_, _21014_);
  and (_21017_, _21016_, _09202_);
  and (_21018_, _07452_, _02693_);
  or (_21019_, _21018_, _21017_);
  and (_21020_, _21019_, _02563_);
  nor (_21021_, _03120_, _02563_);
  nor (_21022_, _21021_, _10433_);
  not (_21023_, _21022_);
  nor (_21025_, _21023_, _21020_);
  or (_21026_, _21025_, _03818_);
  or (_21027_, _21026_, _20995_);
  nand (_21028_, _03818_, _02693_);
  and (_21029_, _21028_, _03821_);
  and (_21030_, _21029_, _21027_);
  or (_21031_, _21030_, _20986_);
  nand (_21032_, _21031_, _09180_);
  nor (_21033_, _09180_, _02693_);
  nor (_21034_, _21033_, _02891_);
  nand (_21036_, _21034_, _21032_);
  and (_21037_, _02891_, _02676_);
  nor (_21038_, _21037_, _05382_);
  nand (_21039_, _21038_, _21036_);
  and (_21040_, _03120_, _05382_);
  nor (_21041_, _21040_, _02947_);
  nand (_21042_, _21041_, _21039_);
  and (_21043_, _02947_, _02676_);
  nor (_21044_, _21043_, _09240_);
  nand (_21045_, _21044_, _21042_);
  nor (_21047_, _09239_, _02693_);
  nor (_21048_, _21047_, _02950_);
  nand (_21049_, _21048_, _21045_);
  and (_21050_, _02950_, _02676_);
  nor (_21051_, _21050_, _09249_);
  nand (_21052_, _21051_, _21049_);
  nor (_21053_, _09247_, _02693_);
  nor (_21054_, _21053_, _02887_);
  nand (_21055_, _21054_, _21052_);
  and (_21056_, _02887_, _02676_);
  nor (_21058_, _21056_, _09251_);
  nand (_21059_, _21058_, _21055_);
  and (_21060_, _03120_, _09251_);
  nor (_21061_, _21060_, _02886_);
  nand (_21062_, _21061_, _21059_);
  and (_21063_, _02886_, _02676_);
  nor (_21064_, _21063_, _09299_);
  and (_21065_, _21064_, _21062_);
  and (_21066_, _09297_, _09074_);
  nor (_21067_, _20983_, _09297_);
  or (_21069_, _21067_, _21066_);
  nor (_21070_, _21069_, _09263_);
  or (_21071_, _21070_, _21065_);
  and (_21072_, _21071_, _09172_);
  or (_21073_, _21072_, _20981_);
  or (_21074_, _21073_, _02966_);
  nor (_21075_, _20983_, _09334_);
  and (_21076_, _09334_, _09074_);
  nor (_21077_, _21076_, _21075_);
  or (_21078_, _21077_, _03377_);
  and (_21080_, _21078_, _21074_);
  or (_21081_, _21080_, _03025_);
  and (_21082_, _09325_, _09074_);
  not (_21083_, _09325_);
  and (_21084_, _20976_, _21083_);
  or (_21085_, _21084_, _21082_);
  and (_21086_, _21085_, _03025_);
  nor (_21087_, _21086_, _09305_);
  and (_21088_, _21087_, _21081_);
  or (_21089_, _21088_, _20972_);
  nand (_21091_, _21089_, _02881_);
  and (_21092_, _02880_, _02677_);
  nor (_21093_, _21092_, _04125_);
  nand (_21094_, _21093_, _21091_);
  nor (_21095_, _03120_, _02561_);
  nor (_21096_, _21095_, _20341_);
  and (_21097_, _21096_, _21094_);
  nor (_21098_, _20340_, _02676_);
  or (_21099_, _21098_, _21097_);
  nand (_21100_, _21099_, _09012_);
  nor (_21102_, _09012_, _02693_);
  nor (_21103_, _21102_, _02987_);
  nand (_21104_, _21103_, _21100_);
  and (_21105_, _02987_, _02676_);
  nor (_21106_, _21105_, _09347_);
  nand (_21107_, _21106_, _21104_);
  and (_21108_, _03120_, _09347_);
  nor (_21109_, _21108_, _02986_);
  nand (_21110_, _21109_, _21107_);
  and (_21111_, _02986_, _02676_);
  nor (_21113_, _21111_, _13666_);
  and (_21114_, _21113_, _21110_);
  nor (_21115_, _09005_, _02693_);
  or (_21116_, _21115_, _21114_);
  nand (_21117_, _21116_, _07596_);
  nor (_21118_, _07596_, _02676_);
  nor (_21119_, _21118_, _02585_);
  nand (_21120_, _21119_, _21117_);
  and (_21121_, _02585_, _02693_);
  nor (_21122_, _21121_, _02874_);
  and (_21124_, _21122_, _21120_);
  or (_21125_, _21124_, _20971_);
  nand (_21126_, _21125_, _05325_);
  and (_21127_, _03120_, _02578_);
  nor (_21128_, _21127_, _03023_);
  nand (_21129_, _21128_, _21126_);
  and (_21130_, _09074_, _03023_);
  nor (_21131_, _21130_, _20391_);
  nand (_21132_, _21131_, _21129_);
  nor (_21133_, _09369_, _02676_);
  nor (_21135_, _21133_, _02576_);
  nand (_21136_, _21135_, _21132_);
  and (_21137_, _09074_, _02576_);
  nor (_21138_, _21137_, _09378_);
  nand (_21139_, _21138_, _21136_);
  nor (_21140_, _09376_, _02693_);
  nor (_21141_, _21140_, _02938_);
  nand (_21142_, _21141_, _21139_);
  and (_21143_, _02938_, _02676_);
  nor (_21144_, _21143_, _02521_);
  nand (_21146_, _21144_, _21142_);
  and (_21147_, _03120_, _02521_);
  nor (_21148_, _21147_, _09384_);
  nand (_21149_, _21148_, _21146_);
  and (_21150_, _20992_, _09384_);
  nor (_21151_, _21150_, _05562_);
  nand (_21152_, _21151_, _21149_);
  nor (_21153_, _05322_, _02676_);
  nor (_21154_, _21153_, _03014_);
  nand (_21155_, _21154_, _21152_);
  and (_21157_, _09074_, _03014_);
  nor (_21158_, _21157_, _07782_);
  and (_21159_, _21158_, _21155_);
  or (_21160_, _21159_, _20970_);
  nand (_21161_, _21160_, _09401_);
  and (_21162_, _09400_, _02688_);
  nor (_21163_, _21162_, _02937_);
  nand (_21164_, _21163_, _21161_);
  and (_21165_, _02937_, _02676_);
  nor (_21166_, _21165_, _02517_);
  nand (_21168_, _21166_, _21164_);
  and (_21169_, _03120_, _02517_);
  nor (_21170_, _21169_, _09000_);
  nand (_21171_, _21170_, _21168_);
  and (_21172_, _08190_, _02676_);
  and (_21173_, _20992_, _08880_);
  or (_21174_, _21173_, _21172_);
  and (_21175_, _21174_, _09000_);
  nor (_21176_, _21175_, _20808_);
  and (_21177_, _21176_, _21171_);
  or (_21179_, _21177_, _20968_);
  nand (_21180_, _21179_, _09450_);
  nor (_21181_, _09450_, _02676_);
  nor (_21182_, _21181_, _03021_);
  and (_21183_, _21182_, _21180_);
  and (_21184_, _09074_, _03021_);
  or (_21185_, _21184_, _03130_);
  nor (_21186_, _21185_, _21183_);
  and (_21187_, _03130_, _02677_);
  or (_21188_, _21187_, _21186_);
  nand (_21190_, _21188_, _02513_);
  and (_21191_, _03120_, _02512_);
  nor (_21192_, _21191_, _08994_);
  nand (_21193_, _21192_, _21190_);
  nor (_21194_, _08190_, _02677_);
  and (_21195_, _20992_, _08190_);
  or (_21196_, _21195_, _21194_);
  and (_21197_, _21196_, _08994_);
  nor (_21198_, _21197_, _20466_);
  and (_21199_, _21198_, _21193_);
  or (_21201_, _21199_, _20967_);
  nand (_21202_, _21201_, _09475_);
  nor (_21203_, _09475_, _02676_);
  nor (_21204_, _21203_, _03020_);
  and (_21205_, _21204_, _21202_);
  and (_21206_, _09074_, _03020_);
  or (_21207_, _21206_, _03139_);
  nor (_21208_, _21207_, _21205_);
  and (_21209_, _03139_, _02677_);
  or (_21210_, _21209_, _21208_);
  nand (_21212_, _21210_, _19955_);
  and (_21213_, _03120_, _02533_);
  nor (_21214_, _21213_, _08875_);
  nand (_21215_, _21214_, _21212_);
  nor (_21216_, _20992_, \oc8051_golden_model_1.PSW [7]);
  nor (_21217_, _02676_, _07319_);
  nor (_21218_, _21217_, _08876_);
  not (_21219_, _21218_);
  nor (_21220_, _21219_, _21216_);
  nor (_21221_, _21220_, _09487_);
  and (_21223_, _21221_, _21215_);
  or (_21224_, _21223_, _20966_);
  nand (_21225_, _21224_, _07866_);
  nor (_21226_, _07866_, _02676_);
  nor (_21227_, _21226_, _03036_);
  and (_21228_, _21227_, _21225_);
  and (_21229_, _09074_, _03036_);
  or (_21230_, _21229_, _03127_);
  nor (_21231_, _21230_, _21228_);
  and (_21232_, _03127_, _02677_);
  or (_21234_, _21232_, _21231_);
  nand (_21235_, _21234_, _19951_);
  and (_21236_, _03120_, _02538_);
  nor (_21237_, _21236_, _08864_);
  nand (_21238_, _21237_, _21235_);
  nor (_21239_, _20992_, _07319_);
  nor (_21240_, _02676_, \oc8051_golden_model_1.PSW [7]);
  nor (_21241_, _21240_, _08865_);
  not (_21242_, _21241_);
  nor (_21243_, _21242_, _21239_);
  nor (_21245_, _21243_, _09503_);
  and (_21246_, _21245_, _21238_);
  or (_21247_, _21246_, _20965_);
  nand (_21248_, _21247_, _08860_);
  nor (_21249_, _08860_, _02676_);
  nor (_21250_, _21249_, _08029_);
  and (_21251_, _21250_, _21248_);
  and (_21252_, _08029_, _02693_);
  or (_21253_, _21252_, _03148_);
  nor (_21254_, _21253_, _21251_);
  and (_21256_, _05984_, _03148_);
  or (_21257_, _21256_, _21254_);
  nand (_21258_, _21257_, _05792_);
  and (_21259_, _03120_, _02531_);
  nor (_21260_, _21259_, _03035_);
  nand (_21261_, _21260_, _21258_);
  and (_21262_, _20983_, _09709_);
  nor (_21263_, _09709_, _09074_);
  or (_21264_, _21263_, _03152_);
  or (_21265_, _21264_, _21262_);
  and (_21267_, _21265_, _08858_);
  and (_21268_, _21267_, _21261_);
  or (_21269_, _21268_, _20964_);
  nand (_21270_, _21269_, _08104_);
  nor (_21271_, _08104_, _02676_);
  nor (_21272_, _21271_, _08135_);
  and (_21273_, _21272_, _21270_);
  and (_21274_, _08135_, _02693_);
  or (_21275_, _21274_, _02897_);
  nor (_21276_, _21275_, _21273_);
  and (_21278_, _05984_, _02897_);
  or (_21279_, _21278_, _21276_);
  nand (_21280_, _21279_, _09728_);
  and (_21281_, _03120_, _02536_);
  nor (_21282_, _21281_, _02895_);
  nand (_21283_, _21282_, _21280_);
  nor (_21284_, _20976_, _09709_);
  and (_21285_, _09709_, _09075_);
  nor (_21286_, _21285_, _21284_);
  and (_21287_, _21286_, _02895_);
  nor (_21289_, _21287_, _09737_);
  nand (_21290_, _21289_, _21283_);
  nor (_21291_, _09736_, _02693_);
  nor (_21292_, _21291_, _03166_);
  and (_21293_, _21292_, _21290_);
  or (_21294_, _21293_, _20963_);
  nand (_21295_, _21294_, _09743_);
  nor (_21296_, _09743_, _02692_);
  nor (_21297_, _21296_, _04159_);
  nand (_21298_, _21297_, _21295_);
  and (_21300_, _04159_, _03120_);
  nor (_21301_, _21300_, _02500_);
  nand (_21302_, _21301_, _21298_);
  and (_21303_, _21286_, _02500_);
  nor (_21304_, _21303_, _09759_);
  nand (_21305_, _21304_, _21302_);
  nor (_21306_, _09758_, _02693_);
  nor (_21307_, _21306_, _03174_);
  and (_21308_, _21307_, _21305_);
  or (_21309_, _21308_, _20962_);
  nand (_21311_, _21309_, _09765_);
  nor (_21312_, _09765_, _02692_);
  nor (_21313_, _21312_, _19938_);
  nand (_21314_, _21313_, _21311_);
  and (_21315_, _19938_, _03120_);
  nor (_21316_, _21315_, _09777_);
  and (_21317_, _21316_, _21314_);
  or (_21318_, _21317_, _20961_);
  or (_21319_, _21318_, _34702_);
  or (_21320_, _34698_, \oc8051_golden_model_1.PC [3]);
  and (_21322_, _21320_, _36029_);
  and (_35242_, _21322_, _21319_);
  and (_21323_, _02233_, \oc8051_golden_model_1.PC [4]);
  nor (_21324_, _02233_, \oc8051_golden_model_1.PC [4]);
  nor (_21325_, _21324_, _21323_);
  and (_21326_, _21325_, _09777_);
  and (_21327_, _05630_, _04159_);
  and (_21328_, _06121_, _03148_);
  nor (_21329_, _08937_, _08190_);
  and (_21330_, _08957_, _08954_);
  nor (_21332_, _21330_, _08958_);
  and (_21333_, _21332_, _08190_);
  or (_21334_, _21333_, _21329_);
  and (_21335_, _21334_, _08994_);
  nor (_21336_, _20340_, _08936_);
  not (_21337_, _21325_);
  and (_21338_, _21337_, _09305_);
  and (_21339_, _09169_, _09069_);
  and (_21340_, _09098_, _09095_);
  nor (_21341_, _21340_, _09099_);
  not (_21343_, _21341_);
  nor (_21344_, _21343_, _09169_);
  nor (_21345_, _21344_, _21339_);
  nor (_21346_, _21345_, _09172_);
  and (_21347_, _08937_, _02887_);
  nor (_21348_, _21325_, _09234_);
  and (_21349_, _05630_, _03824_);
  and (_21350_, _08937_, _03825_);
  or (_21351_, _21350_, _07442_);
  nand (_21352_, _09206_, \oc8051_golden_model_1.PC [4]);
  and (_21354_, _21352_, _03826_);
  or (_21355_, _21354_, _21351_);
  or (_21356_, _21337_, _09207_);
  and (_21357_, _21356_, _02558_);
  and (_21358_, _21357_, _21355_);
  or (_21359_, _21358_, _20635_);
  or (_21360_, _21359_, _21349_);
  or (_21361_, _21337_, _09203_);
  and (_21362_, _21361_, _07433_);
  and (_21363_, _21362_, _21360_);
  and (_21365_, _08937_, _02954_);
  or (_21366_, _21365_, _21363_);
  nor (_21367_, _21366_, _07452_);
  and (_21368_, _21325_, _07452_);
  or (_21369_, _21368_, _21367_);
  and (_21370_, _21369_, _02563_);
  nor (_21371_, _05630_, _02563_);
  nor (_21372_, _21371_, _10433_);
  not (_21373_, _21372_);
  nor (_21374_, _21373_, _21370_);
  nand (_21376_, _21332_, _09198_);
  or (_21377_, _09198_, _08937_);
  and (_21378_, _21377_, _10433_);
  and (_21379_, _21378_, _21376_);
  or (_21380_, _21379_, _21374_);
  nand (_21381_, _21380_, _09228_);
  nand (_21382_, _21341_, _09186_);
  or (_21383_, _09186_, _09070_);
  and (_21384_, _21383_, _02952_);
  nand (_21385_, _21384_, _21382_);
  nand (_21387_, _21385_, _21381_);
  and (_21388_, _21387_, _09180_);
  or (_21389_, _21388_, _21348_);
  nand (_21390_, _21389_, _02892_);
  and (_21391_, _08937_, _02891_);
  nor (_21392_, _21391_, _05382_);
  and (_21393_, _21392_, _21390_);
  nor (_21394_, _05630_, _02556_);
  or (_21395_, _21394_, _02947_);
  nor (_21396_, _21395_, _21393_);
  and (_21398_, _08937_, _02947_);
  or (_21399_, _21398_, _21396_);
  and (_21400_, _21399_, _09239_);
  nor (_21401_, _21325_, _09239_);
  or (_21402_, _21401_, _21400_);
  nand (_21403_, _21402_, _02959_);
  and (_21404_, _08937_, _02950_);
  nor (_21405_, _21404_, _09249_);
  nand (_21406_, _21405_, _21403_);
  nor (_21407_, _21337_, _09247_);
  nor (_21409_, _21407_, _02887_);
  and (_21410_, _21409_, _21406_);
  or (_21411_, _21410_, _21347_);
  nand (_21412_, _21411_, _02568_);
  and (_21413_, _05630_, _09251_);
  nor (_21414_, _21413_, _02886_);
  nand (_21415_, _21414_, _21412_);
  and (_21416_, _08936_, _02886_);
  nor (_21417_, _21416_, _09299_);
  nand (_21418_, _21417_, _21415_);
  and (_21420_, _09297_, _09069_);
  nor (_21421_, _21343_, _09297_);
  or (_21422_, _21421_, _21420_);
  nor (_21423_, _21422_, _09263_);
  nor (_21424_, _21423_, _03038_);
  and (_21425_, _21424_, _21418_);
  nor (_21426_, _21425_, _21346_);
  nor (_21427_, _21426_, _02966_);
  and (_21428_, _09334_, _09069_);
  nor (_21429_, _21343_, _09334_);
  nor (_21431_, _21429_, _21428_);
  nor (_21432_, _21431_, _03377_);
  or (_21433_, _21432_, _21427_);
  nand (_21434_, _21433_, _10029_);
  and (_21435_, _09325_, _09069_);
  and (_21436_, _21341_, _21083_);
  or (_21437_, _21436_, _21435_);
  and (_21438_, _21437_, _03025_);
  nor (_21439_, _21438_, _09305_);
  and (_21440_, _21439_, _21434_);
  or (_21442_, _21440_, _21338_);
  nand (_21443_, _21442_, _02881_);
  and (_21444_, _08937_, _02880_);
  nor (_21445_, _21444_, _04125_);
  nand (_21446_, _21445_, _21443_);
  nor (_21447_, _05630_, _02561_);
  nor (_21448_, _21447_, _20341_);
  and (_21449_, _21448_, _21446_);
  or (_21450_, _21449_, _21336_);
  nand (_21451_, _21450_, _09012_);
  nor (_21453_, _21325_, _09012_);
  nor (_21454_, _21453_, _02987_);
  and (_21455_, _21454_, _21451_);
  and (_21456_, _08936_, _02987_);
  or (_21457_, _21456_, _21455_);
  and (_21458_, _21457_, _02566_);
  nor (_21459_, _05630_, _02566_);
  or (_21460_, _21459_, _02986_);
  or (_21461_, _21460_, _21458_);
  and (_21462_, _08937_, _02986_);
  nor (_21464_, _21462_, _13666_);
  nand (_21465_, _21464_, _21461_);
  nor (_21466_, _21337_, _09005_);
  nor (_21467_, _21466_, _07597_);
  nand (_21468_, _21467_, _21465_);
  nor (_21469_, _08936_, _07596_);
  nor (_21470_, _21469_, _02585_);
  and (_21471_, _21470_, _21468_);
  and (_21472_, _21325_, _02585_);
  or (_21473_, _21472_, _02874_);
  nor (_21475_, _21473_, _21471_);
  and (_21476_, _08937_, _02874_);
  or (_21477_, _21476_, _21475_);
  nand (_21478_, _21477_, _05325_);
  and (_21479_, _05630_, _02578_);
  nor (_21480_, _21479_, _03023_);
  nand (_21481_, _21480_, _21478_);
  and (_21482_, _09069_, _03023_);
  nor (_21483_, _21482_, _20391_);
  nand (_21484_, _21483_, _21481_);
  nor (_21486_, _09369_, _08936_);
  nor (_21487_, _21486_, _02576_);
  and (_21488_, _21487_, _21484_);
  and (_21489_, _09069_, _02576_);
  nor (_21490_, _21489_, _21488_);
  nand (_21491_, _21490_, _09376_);
  nor (_21492_, _21325_, _09376_);
  nor (_21493_, _21492_, _02938_);
  nand (_21494_, _21493_, _21491_);
  nor (_21495_, _08936_, _02521_);
  or (_21497_, _21495_, _09380_);
  nand (_21498_, _21497_, _21494_);
  and (_21499_, _05630_, _02521_);
  nor (_21500_, _21499_, _09384_);
  nand (_21501_, _21500_, _21498_);
  and (_21502_, _21332_, _09384_);
  nor (_21503_, _21502_, _05562_);
  nand (_21504_, _21503_, _21501_);
  nor (_21505_, _08936_, _05322_);
  nor (_21506_, _21505_, _03014_);
  nand (_21508_, _21506_, _21504_);
  and (_21509_, _09069_, _03014_);
  nor (_21510_, _21509_, _07782_);
  and (_21511_, _21510_, _21508_);
  and (_21512_, _08937_, _07782_);
  or (_21513_, _21512_, _21511_);
  nand (_21514_, _21513_, _09401_);
  and (_21515_, _09418_, _09415_);
  nor (_21516_, _21515_, _09419_);
  nor (_21517_, _21516_, _09401_);
  nor (_21519_, _21517_, _02937_);
  nand (_21520_, _21519_, _21514_);
  and (_21521_, _08936_, _02937_);
  nor (_21522_, _21521_, _02517_);
  nand (_21523_, _21522_, _21520_);
  and (_21524_, _05630_, _02517_);
  nor (_21525_, _21524_, _09000_);
  and (_21526_, _21525_, _21523_);
  and (_21527_, _08936_, _08190_);
  and (_21528_, _21332_, _08880_);
  or (_21530_, _21528_, _21527_);
  and (_21531_, _21530_, _09000_);
  or (_21532_, _21531_, _21526_);
  nand (_21533_, _21532_, _09448_);
  nor (_21534_, _21337_, _09448_);
  nor (_21535_, _21534_, _09451_);
  nand (_21536_, _21535_, _21533_);
  nor (_21537_, _08936_, _09450_);
  nor (_21538_, _21537_, _03021_);
  nand (_21539_, _21538_, _21536_);
  and (_21541_, _09069_, _03021_);
  nor (_21542_, _21541_, _03130_);
  and (_21543_, _21542_, _21539_);
  and (_21544_, _08937_, _03130_);
  or (_21545_, _21544_, _21543_);
  nand (_21546_, _21545_, _02513_);
  and (_21547_, _05630_, _02512_);
  nor (_21548_, _21547_, _08994_);
  and (_21549_, _21548_, _21546_);
  or (_21550_, _21549_, _21335_);
  nand (_21552_, _21550_, _09473_);
  nor (_21553_, _21337_, _09473_);
  nor (_21554_, _21553_, _09476_);
  nand (_21555_, _21554_, _21552_);
  nor (_21556_, _08936_, _09475_);
  nor (_21557_, _21556_, _03020_);
  nand (_21558_, _21557_, _21555_);
  and (_21559_, _09069_, _03020_);
  nor (_21560_, _21559_, _03139_);
  and (_21561_, _21560_, _21558_);
  and (_21563_, _08937_, _03139_);
  or (_21564_, _21563_, _21561_);
  nand (_21565_, _21564_, _19955_);
  and (_21566_, _05630_, _02533_);
  nor (_21567_, _21566_, _08875_);
  and (_21568_, _21567_, _21565_);
  and (_21569_, _08936_, \oc8051_golden_model_1.PSW [7]);
  and (_21570_, _21332_, _07319_);
  or (_21571_, _21570_, _21569_);
  and (_21572_, _21571_, _08875_);
  or (_21574_, _21572_, _21568_);
  nand (_21575_, _21574_, _08873_);
  nor (_21576_, _21337_, _08873_);
  nor (_21577_, _21576_, _07867_);
  nand (_21578_, _21577_, _21575_);
  nor (_21579_, _08936_, _07866_);
  nor (_21580_, _21579_, _03036_);
  and (_21581_, _21580_, _21578_);
  and (_21582_, _09069_, _03036_);
  or (_21583_, _21582_, _03127_);
  nor (_21585_, _21583_, _21581_);
  and (_21586_, _08937_, _03127_);
  or (_21587_, _21586_, _21585_);
  nand (_21588_, _21587_, _19951_);
  and (_21589_, _05630_, _02538_);
  nor (_21590_, _21589_, _08864_);
  nand (_21591_, _21590_, _21588_);
  nand (_21592_, _08936_, _07319_);
  nand (_21593_, _21332_, \oc8051_golden_model_1.PSW [7]);
  and (_21594_, _21593_, _21592_);
  or (_21596_, _21594_, _08865_);
  nand (_21597_, _21596_, _21591_);
  nand (_21598_, _21597_, _08862_);
  nor (_21599_, _21337_, _08862_);
  nor (_21600_, _21599_, _08861_);
  nand (_21601_, _21600_, _21598_);
  nor (_21602_, _08936_, _08860_);
  nor (_21603_, _21602_, _08029_);
  nand (_21604_, _21603_, _21601_);
  and (_21605_, _21325_, _08029_);
  nor (_21607_, _21605_, _03148_);
  and (_21608_, _21607_, _21604_);
  or (_21609_, _21608_, _21328_);
  nand (_21610_, _21609_, _05792_);
  and (_21611_, _05630_, _02531_);
  nor (_21612_, _21611_, _03035_);
  and (_21613_, _21612_, _21610_);
  nor (_21614_, _09709_, _09070_);
  and (_21615_, _21341_, _09709_);
  nor (_21616_, _21615_, _21614_);
  nor (_21619_, _21616_, _03152_);
  or (_21620_, _21619_, _21613_);
  nand (_21621_, _21620_, _08858_);
  nor (_21622_, _21337_, _08858_);
  nor (_21623_, _21622_, _08105_);
  nand (_21624_, _21623_, _21621_);
  nor (_21625_, _08936_, _08104_);
  nor (_21626_, _21625_, _08135_);
  nand (_21627_, _21626_, _21624_);
  and (_21628_, _21325_, _08135_);
  nor (_21631_, _21628_, _02897_);
  nand (_21632_, _21631_, _21627_);
  and (_21633_, _06121_, _02897_);
  nor (_21634_, _21633_, _02536_);
  and (_21635_, _21634_, _21632_);
  nor (_21636_, _05630_, _09728_);
  or (_21637_, _21636_, _02895_);
  or (_21638_, _21637_, _21635_);
  and (_21639_, _09709_, _09070_);
  nor (_21640_, _21341_, _09709_);
  nor (_21643_, _21640_, _21639_);
  nor (_21644_, _21643_, _02896_);
  nor (_21645_, _21644_, _09737_);
  nand (_21646_, _21645_, _21638_);
  nor (_21647_, _21337_, _09736_);
  nor (_21648_, _21647_, _03166_);
  nand (_21649_, _21648_, _21646_);
  and (_21650_, _08937_, _03166_);
  nor (_21651_, _21650_, _09744_);
  nand (_21652_, _21651_, _21649_);
  nor (_21655_, _21337_, _09743_);
  nor (_21656_, _21655_, _04159_);
  and (_21657_, _21656_, _21652_);
  or (_21658_, _21657_, _21327_);
  nand (_21659_, _21658_, _02501_);
  nor (_21660_, _21643_, _02501_);
  nor (_21661_, _21660_, _09759_);
  nand (_21662_, _21661_, _21659_);
  nor (_21663_, _21337_, _09758_);
  nor (_21664_, _21663_, _03174_);
  nand (_21667_, _21664_, _21662_);
  and (_21668_, _08937_, _03174_);
  nor (_21669_, _21668_, _09766_);
  nand (_21670_, _21669_, _21667_);
  nor (_21671_, _21337_, _09765_);
  nor (_21672_, _21671_, _19938_);
  nand (_21673_, _21672_, _21670_);
  and (_21674_, _19938_, _05630_);
  nor (_21675_, _21674_, _09777_);
  and (_21676_, _21675_, _21673_);
  or (_21679_, _21676_, _21326_);
  or (_21680_, _21679_, _34702_);
  or (_21681_, _34698_, \oc8051_golden_model_1.PC [4]);
  and (_21682_, _21681_, _36029_);
  and (_35243_, _21682_, _21680_);
  nor (_21683_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_21684_, _08931_, _02247_);
  nor (_21685_, _21684_, _21683_);
  and (_21686_, _21685_, _09777_);
  and (_21687_, _08931_, _03174_);
  nor (_21689_, _21685_, _09743_);
  nor (_21690_, _21685_, _08858_);
  nor (_21691_, _21685_, _08862_);
  nor (_21692_, _21685_, _08873_);
  nor (_21693_, _21685_, _09473_);
  nor (_21694_, _21685_, _09448_);
  and (_21695_, _08932_, _02874_);
  nor (_21696_, _21685_, _09005_);
  nor (_21697_, _20340_, _08931_);
  or (_21698_, _09067_, _09066_);
  not (_21700_, _21698_);
  nor (_21701_, _21700_, _09100_);
  and (_21702_, _21700_, _09100_);
  nor (_21703_, _21702_, _21701_);
  not (_21704_, _21703_);
  nor (_21705_, _21704_, _09169_);
  and (_21706_, _09169_, _09065_);
  nor (_21707_, _21706_, _21705_);
  nor (_21708_, _21707_, _09172_);
  not (_21709_, _09180_);
  and (_21711_, _21703_, _09186_);
  nor (_21712_, _09186_, _09064_);
  nor (_21713_, _21712_, _21711_);
  or (_21714_, _21713_, _03821_);
  and (_21715_, _09196_, _08931_);
  or (_21716_, _08934_, _08933_);
  not (_21717_, _21716_);
  nor (_21718_, _21717_, _08959_);
  and (_21719_, _21717_, _08959_);
  nor (_21720_, _21719_, _21718_);
  nor (_21722_, _21720_, _09196_);
  or (_21723_, _21722_, _21715_);
  nor (_21724_, _21723_, _05387_);
  not (_21725_, \oc8051_golden_model_1.PC [5]);
  and (_21726_, _09206_, _21725_);
  nor (_21727_, _21726_, _03825_);
  and (_21728_, _08931_, _03825_);
  nor (_21729_, _21728_, _07442_);
  not (_21730_, _21729_);
  nor (_21731_, _21730_, _21727_);
  not (_21733_, _21731_);
  nor (_21734_, _21685_, _09207_);
  nor (_21735_, _21734_, _03824_);
  and (_21736_, _21735_, _21733_);
  nor (_21737_, _05661_, _02558_);
  or (_21738_, _21737_, _20635_);
  nor (_21739_, _21738_, _21736_);
  nor (_21740_, _21685_, _09203_);
  nor (_21741_, _21740_, _02954_);
  not (_21742_, _21741_);
  nor (_21744_, _21742_, _21739_);
  and (_21745_, _08931_, _02954_);
  or (_21746_, _21745_, _21744_);
  and (_21747_, _21746_, _09202_);
  and (_21748_, _21685_, _07452_);
  or (_21749_, _21748_, _21747_);
  and (_21750_, _21749_, _02563_);
  nor (_21751_, _05661_, _02563_);
  nor (_21752_, _21751_, _10433_);
  not (_21753_, _21752_);
  nor (_21755_, _21753_, _21750_);
  or (_21756_, _21755_, _03818_);
  nor (_21757_, _21756_, _21724_);
  and (_21758_, _21685_, _03818_);
  or (_21759_, _21758_, _02952_);
  or (_21760_, _21759_, _21757_);
  and (_21761_, _21760_, _21714_);
  nor (_21762_, _21761_, _21709_);
  nor (_21763_, _21685_, _09180_);
  nor (_21764_, _21763_, _02891_);
  not (_21766_, _21764_);
  nor (_21767_, _21766_, _21762_);
  and (_21768_, _08931_, _02891_);
  nor (_21769_, _21768_, _21767_);
  or (_21770_, _21769_, _05382_);
  or (_21771_, _05661_, _02556_);
  and (_21772_, _21771_, _21770_);
  or (_21773_, _21772_, _02947_);
  and (_21774_, _08931_, _02947_);
  nor (_21775_, _21774_, _09240_);
  nand (_21777_, _21775_, _21773_);
  nor (_21778_, _21685_, _09239_);
  nor (_21779_, _21778_, _02950_);
  nand (_21780_, _21779_, _21777_);
  and (_21781_, _08931_, _02950_);
  nor (_21782_, _21781_, _09249_);
  nand (_21783_, _21782_, _21780_);
  nor (_21784_, _21685_, _09247_);
  nor (_21785_, _21784_, _02887_);
  nand (_21786_, _21785_, _21783_);
  and (_21788_, _08931_, _02887_);
  nor (_21789_, _21788_, _09251_);
  nand (_21790_, _21789_, _21786_);
  and (_21791_, _05661_, _09251_);
  nor (_21792_, _21791_, _02886_);
  nand (_21793_, _21792_, _21790_);
  and (_21794_, _08931_, _02886_);
  nor (_21795_, _21794_, _09299_);
  and (_21796_, _21795_, _21793_);
  and (_21797_, _09297_, _09064_);
  nor (_21799_, _21703_, _09297_);
  or (_21800_, _21799_, _21797_);
  nor (_21801_, _21800_, _09263_);
  or (_21802_, _21801_, _21796_);
  and (_21803_, _21802_, _09172_);
  or (_21804_, _21803_, _21708_);
  or (_21805_, _21804_, _02966_);
  nor (_21806_, _21703_, _09334_);
  and (_21807_, _09334_, _09064_);
  nor (_21808_, _21807_, _21806_);
  or (_21810_, _21808_, _03377_);
  and (_21811_, _21810_, _21805_);
  or (_21812_, _21811_, _03025_);
  nand (_21813_, _09325_, _09064_);
  or (_21814_, _21703_, _09325_);
  and (_21815_, _21814_, _21813_);
  or (_21816_, _21815_, _10029_);
  and (_21817_, _21816_, _21812_);
  or (_21818_, _21817_, _09305_);
  nand (_21819_, _21685_, _09305_);
  and (_21821_, _21819_, _21818_);
  nand (_21822_, _21821_, _02881_);
  and (_21823_, _08932_, _02880_);
  nor (_21824_, _21823_, _04125_);
  nand (_21825_, _21824_, _21822_);
  nor (_21826_, _05661_, _02561_);
  nor (_21827_, _21826_, _20341_);
  and (_21828_, _21827_, _21825_);
  or (_21829_, _21828_, _21697_);
  nand (_21830_, _21829_, _09012_);
  nor (_21832_, _21685_, _09012_);
  nor (_21833_, _21832_, _02987_);
  nand (_21834_, _21833_, _21830_);
  and (_21835_, _08931_, _02987_);
  nor (_21836_, _21835_, _09347_);
  nand (_21837_, _21836_, _21834_);
  and (_21838_, _05661_, _09347_);
  nor (_21839_, _21838_, _02986_);
  nand (_21840_, _21839_, _21837_);
  and (_21841_, _08931_, _02986_);
  nor (_21843_, _21841_, _13666_);
  and (_21844_, _21843_, _21840_);
  or (_21845_, _21844_, _21696_);
  nand (_21846_, _21845_, _07596_);
  nor (_21847_, _08931_, _07596_);
  nor (_21848_, _21847_, _02585_);
  nand (_21849_, _21848_, _21846_);
  and (_21850_, _21685_, _02585_);
  nor (_21851_, _21850_, _02874_);
  and (_21852_, _21851_, _21849_);
  or (_21854_, _21852_, _21695_);
  nand (_21855_, _21854_, _05325_);
  and (_21856_, _05661_, _02578_);
  nor (_21857_, _21856_, _03023_);
  nand (_21858_, _21857_, _21855_);
  and (_21859_, _09064_, _03023_);
  nor (_21860_, _21859_, _20391_);
  nand (_21861_, _21860_, _21858_);
  nor (_21862_, _09369_, _08931_);
  nor (_21863_, _21862_, _02576_);
  nand (_21865_, _21863_, _21861_);
  and (_21866_, _09064_, _02576_);
  nor (_21867_, _21866_, _09378_);
  nand (_21868_, _21867_, _21865_);
  nor (_21869_, _21685_, _09376_);
  nor (_21870_, _21869_, _02938_);
  nand (_21871_, _21870_, _21868_);
  and (_21872_, _08931_, _02938_);
  nor (_21873_, _21872_, _02521_);
  nand (_21874_, _21873_, _21871_);
  and (_21876_, _05661_, _02521_);
  nor (_21877_, _21876_, _09384_);
  nand (_21878_, _21877_, _21874_);
  nor (_21879_, _21720_, _09385_);
  nor (_21880_, _21879_, _05562_);
  nand (_21881_, _21880_, _21878_);
  nor (_21882_, _08931_, _05322_);
  nor (_21883_, _21882_, _03014_);
  nand (_21884_, _21883_, _21881_);
  and (_21885_, _09064_, _03014_);
  nor (_21887_, _21885_, _07782_);
  and (_21888_, _21887_, _21884_);
  and (_21889_, _08932_, _07782_);
  or (_21890_, _21889_, _21888_);
  nand (_21891_, _21890_, _09401_);
  and (_21892_, _09420_, _09413_);
  nor (_21893_, _21892_, _09421_);
  nor (_21894_, _21893_, _09401_);
  nor (_21895_, _21894_, _02937_);
  nand (_21896_, _21895_, _21891_);
  and (_21898_, _08931_, _02937_);
  nor (_21899_, _21898_, _02517_);
  nand (_21900_, _21899_, _21896_);
  and (_21901_, _05661_, _02517_);
  nor (_21902_, _21901_, _09000_);
  nand (_21903_, _21902_, _21900_);
  and (_21904_, _08931_, _08190_);
  nor (_21905_, _21720_, _08190_);
  or (_21906_, _21905_, _21904_);
  and (_21907_, _21906_, _09000_);
  nor (_21909_, _21907_, _20808_);
  and (_21910_, _21909_, _21903_);
  or (_21911_, _21910_, _21694_);
  nand (_21912_, _21911_, _09450_);
  nor (_21913_, _08931_, _09450_);
  nor (_21914_, _21913_, _03021_);
  and (_21915_, _21914_, _21912_);
  and (_21916_, _09064_, _03021_);
  or (_21917_, _21916_, _03130_);
  nor (_21918_, _21917_, _21915_);
  and (_21920_, _08932_, _03130_);
  or (_21921_, _21920_, _21918_);
  nand (_21922_, _21921_, _02513_);
  and (_21923_, _05661_, _02512_);
  nor (_21924_, _21923_, _08994_);
  nand (_21925_, _21924_, _21922_);
  and (_21926_, _08931_, _08880_);
  nor (_21927_, _21720_, _08880_);
  or (_21928_, _21927_, _21926_);
  and (_21929_, _21928_, _08994_);
  nor (_21931_, _21929_, _20466_);
  and (_21932_, _21931_, _21925_);
  or (_21933_, _21932_, _21693_);
  nand (_21934_, _21933_, _09475_);
  nor (_21935_, _08931_, _09475_);
  nor (_21936_, _21935_, _03020_);
  and (_21937_, _21936_, _21934_);
  and (_21938_, _09064_, _03020_);
  or (_21939_, _21938_, _03139_);
  nor (_21940_, _21939_, _21937_);
  and (_21942_, _08932_, _03139_);
  or (_21943_, _21942_, _21940_);
  nand (_21944_, _21943_, _19955_);
  and (_21945_, _05661_, _02533_);
  nor (_21946_, _21945_, _08875_);
  nand (_21947_, _21946_, _21944_);
  and (_21948_, _08931_, \oc8051_golden_model_1.PSW [7]);
  nor (_21949_, _21720_, \oc8051_golden_model_1.PSW [7]);
  or (_21950_, _21949_, _21948_);
  and (_21951_, _21950_, _08875_);
  nor (_21953_, _21951_, _09487_);
  and (_21954_, _21953_, _21947_);
  or (_21955_, _21954_, _21692_);
  nand (_21956_, _21955_, _07866_);
  nor (_21957_, _08931_, _07866_);
  nor (_21958_, _21957_, _03036_);
  nand (_21959_, _21958_, _21956_);
  and (_21960_, _09064_, _03036_);
  nor (_21961_, _21960_, _03127_);
  and (_21962_, _21961_, _21959_);
  and (_21964_, _08932_, _03127_);
  or (_21965_, _21964_, _21962_);
  nand (_21966_, _21965_, _19951_);
  and (_21967_, _05661_, _02538_);
  nor (_21968_, _21967_, _08864_);
  nand (_21969_, _21968_, _21966_);
  and (_21970_, _08931_, _07319_);
  nor (_21971_, _21720_, _07319_);
  or (_21972_, _21971_, _21970_);
  and (_21973_, _21972_, _08864_);
  nor (_21975_, _21973_, _09503_);
  and (_21976_, _21975_, _21969_);
  or (_21977_, _21976_, _21691_);
  nand (_21978_, _21977_, _08860_);
  nor (_21979_, _08931_, _08860_);
  nor (_21980_, _21979_, _08029_);
  and (_21981_, _21980_, _21978_);
  and (_21982_, _21685_, _08029_);
  or (_21983_, _21982_, _03148_);
  nor (_21984_, _21983_, _21981_);
  and (_21986_, _06076_, _03148_);
  or (_21987_, _21986_, _21984_);
  nand (_21988_, _21987_, _05792_);
  and (_21989_, _05661_, _02531_);
  nor (_21990_, _21989_, _03035_);
  nand (_21991_, _21990_, _21988_);
  nor (_21992_, _09709_, _09064_);
  and (_21993_, _21703_, _09709_);
  or (_21994_, _21993_, _03152_);
  or (_21995_, _21994_, _21992_);
  and (_21997_, _21995_, _08858_);
  and (_21998_, _21997_, _21991_);
  or (_21999_, _21998_, _21690_);
  nand (_22000_, _21999_, _08104_);
  nor (_22001_, _08931_, _08104_);
  nor (_22002_, _22001_, _08135_);
  nand (_22003_, _22002_, _22000_);
  and (_22004_, _21685_, _08135_);
  nor (_22005_, _22004_, _02897_);
  and (_22006_, _22005_, _22003_);
  and (_22008_, _06076_, _02897_);
  or (_22009_, _22008_, _22006_);
  nand (_22010_, _22009_, _09728_);
  and (_22011_, _05661_, _02536_);
  nor (_22012_, _22011_, _02895_);
  nand (_22013_, _22012_, _22010_);
  nor (_22014_, _21704_, _09709_);
  and (_22015_, _09709_, _09065_);
  nor (_22016_, _22015_, _22014_);
  and (_22017_, _22016_, _02895_);
  nor (_22019_, _22017_, _09737_);
  nand (_22020_, _22019_, _22013_);
  nor (_22021_, _21685_, _09736_);
  nor (_22022_, _22021_, _03166_);
  nand (_22023_, _22022_, _22020_);
  and (_22024_, _08931_, _03166_);
  nor (_22025_, _22024_, _09744_);
  and (_22026_, _22025_, _22023_);
  or (_22027_, _22026_, _21689_);
  nand (_22028_, _22027_, _03916_);
  and (_22030_, _05661_, _04159_);
  nor (_22031_, _22030_, _02500_);
  nand (_22032_, _22031_, _22028_);
  and (_22033_, _22016_, _02500_);
  nor (_22034_, _22033_, _09759_);
  nand (_22035_, _22034_, _22032_);
  nor (_22036_, _21685_, _09758_);
  nor (_22037_, _22036_, _03174_);
  and (_22038_, _22037_, _22035_);
  or (_22039_, _22038_, _21687_);
  nand (_22041_, _22039_, _09765_);
  and (_22042_, _21685_, _09766_);
  nor (_22043_, _22042_, _19938_);
  nand (_22044_, _22043_, _22041_);
  and (_22045_, _19938_, _05661_);
  nor (_22046_, _22045_, _09777_);
  and (_22047_, _22046_, _22044_);
  or (_22048_, _22047_, _21686_);
  or (_22049_, _22048_, _34702_);
  or (_22050_, _34698_, \oc8051_golden_model_1.PC [5]);
  and (_22052_, _22050_, _36029_);
  and (_35244_, _22052_, _22049_);
  and (_22053_, _05389_, _02233_);
  nor (_22054_, _22053_, \oc8051_golden_model_1.PC [6]);
  nor (_22055_, _22054_, _08841_);
  and (_22056_, _22055_, _09777_);
  and (_22057_, _05598_, _04159_);
  not (_22058_, _22055_);
  and (_22059_, _22058_, _08135_);
  and (_22060_, _09057_, _03036_);
  and (_22062_, _09057_, _03020_);
  and (_22063_, _09057_, _03021_);
  and (_22064_, _08961_, _08928_);
  nor (_22065_, _22064_, _08962_);
  and (_22066_, _22065_, _09384_);
  and (_22067_, _22058_, _02585_);
  and (_22068_, _22058_, _09305_);
  and (_22069_, _09102_, _09061_);
  nor (_22070_, _22069_, _09103_);
  not (_22071_, _22070_);
  nor (_22073_, _22071_, _09169_);
  and (_22074_, _09169_, _09056_);
  nor (_22075_, _22074_, _22073_);
  nor (_22076_, _22075_, _09172_);
  and (_22077_, _08924_, _02887_);
  nor (_22078_, _22055_, _09234_);
  and (_22079_, _05598_, _03824_);
  and (_22080_, _08924_, _03825_);
  or (_22081_, _22080_, _07442_);
  nand (_22082_, _09206_, \oc8051_golden_model_1.PC [6]);
  and (_22084_, _22082_, _03826_);
  or (_22085_, _22084_, _22081_);
  or (_22086_, _22058_, _09207_);
  and (_22087_, _22086_, _02558_);
  and (_22088_, _22087_, _22085_);
  or (_22089_, _22088_, _20635_);
  or (_22090_, _22089_, _22079_);
  or (_22091_, _22058_, _09203_);
  and (_22092_, _22091_, _07433_);
  and (_22093_, _22092_, _22090_);
  and (_22095_, _08924_, _02954_);
  or (_22096_, _22095_, _22093_);
  nor (_22097_, _22096_, _07452_);
  and (_22098_, _22055_, _07452_);
  or (_22099_, _22098_, _22097_);
  and (_22100_, _22099_, _02563_);
  nor (_22101_, _05598_, _02563_);
  nor (_22102_, _22101_, _10433_);
  not (_22103_, _22102_);
  nor (_22104_, _22103_, _22100_);
  nand (_22106_, _22065_, _09198_);
  or (_22107_, _09198_, _08924_);
  and (_22108_, _22107_, _10433_);
  and (_22109_, _22108_, _22106_);
  or (_22110_, _22109_, _22104_);
  nand (_22111_, _22110_, _09228_);
  nand (_22112_, _22070_, _09186_);
  or (_22113_, _09186_, _09057_);
  and (_22114_, _22113_, _02952_);
  nand (_22115_, _22114_, _22112_);
  nand (_22117_, _22115_, _22111_);
  and (_22118_, _22117_, _09180_);
  or (_22119_, _22118_, _22078_);
  nand (_22120_, _22119_, _02892_);
  and (_22121_, _08924_, _02891_);
  nor (_22122_, _22121_, _05382_);
  nand (_22123_, _22122_, _22120_);
  nor (_22124_, _05598_, _02556_);
  nor (_22125_, _22124_, _02947_);
  and (_22126_, _22125_, _22123_);
  and (_22128_, _08924_, _02947_);
  or (_22129_, _22128_, _22126_);
  or (_22130_, _22129_, _09240_);
  or (_22131_, _22058_, _09239_);
  and (_22132_, _22131_, _02959_);
  nand (_22133_, _22132_, _22130_);
  and (_22134_, _08924_, _02950_);
  nor (_22135_, _22134_, _09249_);
  nand (_22136_, _22135_, _22133_);
  nor (_22137_, _22058_, _09247_);
  nor (_22139_, _22137_, _02887_);
  and (_22140_, _22139_, _22136_);
  or (_22141_, _22140_, _22077_);
  nand (_22142_, _22141_, _02568_);
  and (_22143_, _05598_, _09251_);
  nor (_22144_, _22143_, _02886_);
  nand (_22145_, _22144_, _22142_);
  and (_22146_, _08923_, _02886_);
  nor (_22147_, _22146_, _09299_);
  nand (_22148_, _22147_, _22145_);
  and (_22150_, _09297_, _09056_);
  nor (_22151_, _22071_, _09297_);
  or (_22152_, _22151_, _22150_);
  nor (_22153_, _22152_, _09263_);
  nor (_22154_, _22153_, _03038_);
  and (_22155_, _22154_, _22148_);
  nor (_22156_, _22155_, _22076_);
  nor (_22157_, _22156_, _02966_);
  and (_22158_, _09334_, _09056_);
  nor (_22159_, _22071_, _09334_);
  nor (_22161_, _22159_, _22158_);
  nor (_22162_, _22161_, _03377_);
  or (_22163_, _22162_, _22157_);
  nand (_22164_, _22163_, _10029_);
  and (_22165_, _09325_, _09056_);
  and (_22166_, _22070_, _21083_);
  or (_22167_, _22166_, _22165_);
  and (_22168_, _22167_, _03025_);
  nor (_22169_, _22168_, _09305_);
  and (_22170_, _22169_, _22164_);
  or (_22172_, _22170_, _22068_);
  nand (_22173_, _22172_, _02881_);
  and (_22174_, _08924_, _02880_);
  nor (_22175_, _22174_, _04125_);
  nand (_22176_, _22175_, _22173_);
  nor (_22177_, _05598_, _02561_);
  nor (_22178_, _22177_, _20341_);
  and (_22179_, _22178_, _22176_);
  nor (_22180_, _20340_, _08923_);
  or (_22181_, _22180_, _22179_);
  nand (_22182_, _22181_, _09012_);
  nor (_22183_, _22055_, _09012_);
  nor (_22184_, _22183_, _02987_);
  nand (_22185_, _22184_, _22182_);
  and (_22186_, _08923_, _02987_);
  nor (_22187_, _22186_, _09347_);
  nand (_22188_, _22187_, _22185_);
  and (_22189_, _05598_, _09347_);
  nor (_22190_, _22189_, _02986_);
  and (_22191_, _22190_, _22188_);
  and (_22194_, _08923_, _02986_);
  nor (_22195_, _22194_, _22191_);
  nand (_22196_, _22195_, _09005_);
  nor (_22197_, _22055_, _09005_);
  nor (_22198_, _22197_, _07597_);
  nand (_22199_, _22198_, _22196_);
  nor (_22200_, _08924_, _07596_);
  nor (_22201_, _22200_, _02585_);
  and (_22202_, _22201_, _22199_);
  or (_22203_, _22202_, _22067_);
  nand (_22205_, _22203_, _02875_);
  and (_22206_, _08924_, _02874_);
  nor (_22207_, _22206_, _02578_);
  and (_22208_, _22207_, _22205_);
  nor (_22209_, _05598_, _05325_);
  or (_22210_, _22209_, _03023_);
  nor (_22211_, _22210_, _22208_);
  and (_22212_, _09057_, _03023_);
  or (_22213_, _22212_, _22211_);
  and (_22214_, _22213_, _09369_);
  nor (_22216_, _09369_, _08923_);
  or (_22217_, _22216_, _22214_);
  nand (_22218_, _22217_, _02851_);
  and (_22219_, _09057_, _02576_);
  nor (_22220_, _22219_, _09378_);
  nand (_22221_, _22220_, _22218_);
  nor (_22222_, _22058_, _09376_);
  nor (_22223_, _22222_, _02938_);
  nand (_22224_, _22223_, _22221_);
  and (_22225_, _08924_, _02938_);
  nor (_22227_, _22225_, _02521_);
  and (_22228_, _22227_, _22224_);
  nor (_22229_, _05598_, _20078_);
  or (_22230_, _22229_, _22228_);
  and (_22231_, _22230_, _09385_);
  nor (_22232_, _22231_, _22066_);
  or (_22233_, _22232_, _05562_);
  or (_22234_, _08924_, _05322_);
  and (_22235_, _22234_, _03884_);
  nand (_22236_, _22235_, _22233_);
  and (_22238_, _09057_, _03014_);
  nor (_22239_, _22238_, _07782_);
  nand (_22240_, _22239_, _22236_);
  and (_22241_, _08923_, _07782_);
  nor (_22242_, _22241_, _09400_);
  nand (_22243_, _22242_, _22240_);
  and (_22244_, _09422_, _09409_);
  nor (_22245_, _22244_, _09423_);
  nor (_22246_, _22245_, _09401_);
  nor (_22247_, _22246_, _02937_);
  nand (_22249_, _22247_, _22243_);
  and (_22250_, _08923_, _02937_);
  nor (_22251_, _22250_, _02517_);
  nand (_22252_, _22251_, _22249_);
  and (_22253_, _05598_, _02517_);
  nor (_22254_, _22253_, _09000_);
  nand (_22255_, _22254_, _22252_);
  and (_22256_, _08923_, _08190_);
  and (_22257_, _22065_, _08880_);
  or (_22258_, _22257_, _22256_);
  and (_22260_, _22258_, _09000_);
  nor (_22261_, _22260_, _20808_);
  nand (_22262_, _22261_, _22255_);
  nor (_22263_, _22055_, _09448_);
  nor (_22264_, _22263_, _09451_);
  nand (_22265_, _22264_, _22262_);
  nor (_22266_, _08924_, _09450_);
  nor (_22267_, _22266_, _03021_);
  and (_22268_, _22267_, _22265_);
  or (_22269_, _22268_, _22063_);
  nand (_22271_, _22269_, _03131_);
  and (_22272_, _08924_, _03130_);
  nor (_22273_, _22272_, _02512_);
  and (_22274_, _22273_, _22271_);
  nor (_22275_, _05598_, _02513_);
  or (_22276_, _22275_, _22274_);
  nand (_22277_, _22276_, _09462_);
  and (_22278_, _08923_, _08880_);
  and (_22279_, _22065_, _08190_);
  or (_22280_, _22279_, _22278_);
  and (_22282_, _22280_, _08994_);
  nor (_22283_, _22282_, _20466_);
  nand (_22284_, _22283_, _22277_);
  nor (_22285_, _22055_, _09473_);
  nor (_22286_, _22285_, _09476_);
  nand (_22287_, _22286_, _22284_);
  nor (_22288_, _08924_, _09475_);
  nor (_22289_, _22288_, _03020_);
  and (_22290_, _22289_, _22287_);
  or (_22291_, _22290_, _22062_);
  nand (_22293_, _22291_, _03140_);
  and (_22294_, _08924_, _03139_);
  nor (_22295_, _22294_, _02533_);
  and (_22296_, _22295_, _22293_);
  nor (_22297_, _05598_, _19955_);
  or (_22298_, _22297_, _22296_);
  nand (_22299_, _22298_, _08876_);
  nor (_22300_, _22065_, \oc8051_golden_model_1.PSW [7]);
  nor (_22301_, _08923_, _07319_);
  nor (_22302_, _22301_, _08876_);
  not (_22304_, _22302_);
  nor (_22305_, _22304_, _22300_);
  nor (_22306_, _22305_, _09487_);
  nand (_22307_, _22306_, _22299_);
  nor (_22308_, _22055_, _08873_);
  nor (_22309_, _22308_, _07867_);
  nand (_22310_, _22309_, _22307_);
  nor (_22311_, _08924_, _07866_);
  nor (_22312_, _22311_, _03036_);
  and (_22313_, _22312_, _22310_);
  or (_22315_, _22313_, _22060_);
  nand (_22316_, _22315_, _05786_);
  and (_22317_, _08924_, _03127_);
  nor (_22318_, _22317_, _02538_);
  and (_22319_, _22318_, _22316_);
  nor (_22320_, _05598_, _19951_);
  or (_22321_, _22320_, _22319_);
  nand (_22322_, _22321_, _08865_);
  nor (_22323_, _22065_, _07319_);
  nor (_22324_, _08923_, \oc8051_golden_model_1.PSW [7]);
  nor (_22326_, _22324_, _08865_);
  not (_22327_, _22326_);
  nor (_22328_, _22327_, _22323_);
  nor (_22329_, _22328_, _09503_);
  nand (_22330_, _22329_, _22322_);
  nor (_22331_, _22055_, _08862_);
  nor (_22332_, _22331_, _08861_);
  nand (_22333_, _22332_, _22330_);
  nor (_22334_, _08924_, _08860_);
  nor (_22335_, _22334_, _08029_);
  nand (_22337_, _22335_, _22333_);
  and (_22338_, _22058_, _08029_);
  nor (_22339_, _22338_, _03148_);
  and (_22340_, _22339_, _22337_);
  and (_22341_, _05847_, _03148_);
  or (_22342_, _22341_, _02531_);
  or (_22343_, _22342_, _22340_);
  and (_22344_, _05598_, _02531_);
  nor (_22345_, _22344_, _03035_);
  nand (_22346_, _22345_, _22343_);
  and (_22348_, _22071_, _09709_);
  nor (_22349_, _09709_, _09056_);
  or (_22350_, _22349_, _03152_);
  or (_22351_, _22350_, _22348_);
  and (_22352_, _22351_, _08858_);
  nand (_22353_, _22352_, _22346_);
  nor (_22354_, _22055_, _08858_);
  nor (_22355_, _22354_, _08105_);
  nand (_22356_, _22355_, _22353_);
  nor (_22357_, _08924_, _08104_);
  nor (_22359_, _22357_, _08135_);
  and (_22360_, _22359_, _22356_);
  or (_22361_, _22360_, _22059_);
  nand (_22362_, _22361_, _02898_);
  nor (_22363_, _05847_, _02898_);
  nor (_22364_, _22363_, _02536_);
  and (_22365_, _22364_, _22362_);
  nor (_22366_, _05598_, _09728_);
  or (_22367_, _22366_, _02895_);
  nor (_22368_, _22367_, _22365_);
  and (_22370_, _09709_, _09057_);
  nor (_22371_, _22070_, _09709_);
  nor (_22372_, _22371_, _22370_);
  nor (_22373_, _22372_, _02896_);
  or (_22374_, _22373_, _22368_);
  and (_22375_, _22374_, _09736_);
  nor (_22376_, _22055_, _09736_);
  or (_22377_, _22376_, _22375_);
  nand (_22378_, _22377_, _03563_);
  and (_22379_, _08924_, _03166_);
  nor (_22380_, _22379_, _09744_);
  nand (_22381_, _22380_, _22378_);
  nor (_22382_, _22058_, _09743_);
  nor (_22383_, _22382_, _04159_);
  and (_22384_, _22383_, _22381_);
  or (_22385_, _22384_, _22057_);
  nand (_22386_, _22385_, _02501_);
  nor (_22387_, _22372_, _02501_);
  nor (_22388_, _22387_, _09759_);
  nand (_22389_, _22388_, _22386_);
  nor (_22391_, _22058_, _09758_);
  nor (_22392_, _22391_, _03174_);
  nand (_22393_, _22392_, _22389_);
  and (_22394_, _08924_, _03174_);
  nor (_22395_, _22394_, _09766_);
  nand (_22396_, _22395_, _22393_);
  nor (_22397_, _22058_, _09765_);
  nor (_22398_, _22397_, _19938_);
  nand (_22399_, _22398_, _22396_);
  and (_22400_, _19938_, _05598_);
  nor (_22402_, _22400_, _09777_);
  and (_22403_, _22402_, _22399_);
  or (_22404_, _22403_, _22056_);
  or (_22405_, _22404_, _34702_);
  or (_22406_, _34698_, \oc8051_golden_model_1.PC [6]);
  and (_22407_, _22406_, _36029_);
  and (_35245_, _22407_, _22405_);
  nor (_22408_, _08841_, \oc8051_golden_model_1.PC [7]);
  nor (_22409_, _22408_, _08842_);
  and (_22410_, _22409_, _09777_);
  and (_22411_, _05394_, _03174_);
  and (_22412_, _05394_, _03166_);
  nor (_22413_, _22409_, _08858_);
  nor (_22414_, _22409_, _08862_);
  nor (_22415_, _22409_, _08873_);
  nor (_22416_, _22409_, _09473_);
  nor (_22417_, _22409_, _09448_);
  nor (_22418_, _20340_, _05394_);
  not (_22419_, _22409_);
  and (_22420_, _22419_, _09305_);
  or (_22421_, _09052_, _09053_);
  and (_22422_, _22421_, _09104_);
  nor (_22423_, _22421_, _09104_);
  nor (_22424_, _22423_, _22422_);
  nor (_22425_, _22424_, _09169_);
  and (_22426_, _09169_, _06139_);
  nor (_22427_, _22426_, _22425_);
  nor (_22428_, _22427_, _09172_);
  nor (_22429_, _09186_, _06138_);
  not (_22430_, _22424_);
  and (_22431_, _22430_, _09186_);
  nor (_22432_, _22431_, _22429_);
  or (_22433_, _22432_, _03821_);
  and (_22434_, _09196_, _05394_);
  or (_22435_, _08919_, _08920_);
  and (_22436_, _22435_, _08963_);
  nor (_22437_, _22435_, _08963_);
  nor (_22438_, _22437_, _22436_);
  and (_22439_, _22438_, _09198_);
  or (_22440_, _22439_, _22434_);
  nor (_22442_, _22440_, _05387_);
  not (_22443_, \oc8051_golden_model_1.PC [7]);
  and (_22444_, _09206_, _22443_);
  nor (_22445_, _22444_, _03825_);
  and (_22446_, _05394_, _03825_);
  nor (_22447_, _22446_, _07442_);
  not (_22448_, _22447_);
  nor (_22449_, _22448_, _22445_);
  not (_22450_, _22449_);
  nor (_22451_, _22409_, _09207_);
  nor (_22452_, _22451_, _03824_);
  and (_22453_, _22452_, _22450_);
  nor (_22454_, _05311_, _02558_);
  or (_22455_, _22454_, _20635_);
  nor (_22456_, _22455_, _22453_);
  nor (_22457_, _22409_, _09203_);
  nor (_22458_, _22457_, _02954_);
  not (_22459_, _22458_);
  nor (_22460_, _22459_, _22456_);
  and (_22461_, _05394_, _02954_);
  or (_22463_, _22461_, _22460_);
  and (_22464_, _22463_, _09202_);
  and (_22465_, _22409_, _07452_);
  or (_22466_, _22465_, _22464_);
  and (_22467_, _22466_, _02563_);
  nor (_22468_, _05311_, _02563_);
  nor (_22469_, _22468_, _10433_);
  not (_22470_, _22469_);
  nor (_22471_, _22470_, _22467_);
  or (_22472_, _22471_, _03818_);
  nor (_22474_, _22472_, _22442_);
  and (_22475_, _22409_, _03818_);
  or (_22476_, _22475_, _02952_);
  or (_22477_, _22476_, _22474_);
  and (_22478_, _22477_, _22433_);
  nor (_22479_, _22478_, _21709_);
  nor (_22480_, _22409_, _09180_);
  nor (_22481_, _22480_, _02891_);
  not (_22482_, _22481_);
  or (_22483_, _22482_, _22479_);
  and (_22484_, _05394_, _02891_);
  nor (_22485_, _22484_, _05382_);
  nand (_22486_, _22485_, _22483_);
  and (_22487_, _05311_, _05382_);
  nor (_22488_, _22487_, _02947_);
  nand (_22489_, _22488_, _22486_);
  and (_22490_, _05394_, _02947_);
  nor (_22491_, _22490_, _09240_);
  nand (_22492_, _22491_, _22489_);
  nor (_22493_, _22409_, _09239_);
  nor (_22495_, _22493_, _02950_);
  nand (_22496_, _22495_, _22492_);
  and (_22497_, _05394_, _02950_);
  nor (_22498_, _22497_, _09249_);
  nand (_22499_, _22498_, _22496_);
  nor (_22500_, _22409_, _09247_);
  nor (_22501_, _22500_, _02887_);
  nand (_22502_, _22501_, _22499_);
  and (_22503_, _05394_, _02887_);
  nor (_22504_, _22503_, _09251_);
  nand (_22506_, _22504_, _22502_);
  and (_22507_, _05311_, _09251_);
  nor (_22508_, _22507_, _02886_);
  nand (_22509_, _22508_, _22506_);
  and (_22510_, _05394_, _02886_);
  nor (_22511_, _22510_, _09299_);
  and (_22512_, _22511_, _22509_);
  and (_22513_, _09297_, _06138_);
  nor (_22514_, _22430_, _09297_);
  or (_22515_, _22514_, _22513_);
  nor (_22517_, _22515_, _09263_);
  or (_22518_, _22517_, _22512_);
  and (_22519_, _22518_, _09172_);
  or (_22520_, _22519_, _22428_);
  or (_22521_, _22520_, _02966_);
  nor (_22522_, _22430_, _09334_);
  and (_22523_, _09334_, _06138_);
  nor (_22524_, _22523_, _22522_);
  or (_22525_, _22524_, _03377_);
  and (_22526_, _22525_, _22521_);
  or (_22528_, _22526_, _03025_);
  and (_22529_, _09325_, _06138_);
  and (_22530_, _22424_, _21083_);
  or (_22531_, _22530_, _22529_);
  and (_22532_, _22531_, _03025_);
  nor (_22533_, _22532_, _09305_);
  and (_22534_, _22533_, _22528_);
  or (_22535_, _22534_, _22420_);
  nand (_22536_, _22535_, _02881_);
  and (_22537_, _05395_, _02880_);
  nor (_22538_, _22537_, _04125_);
  nand (_22539_, _22538_, _22536_);
  nor (_22540_, _05311_, _02561_);
  nor (_22541_, _22540_, _20341_);
  and (_22542_, _22541_, _22539_);
  or (_22543_, _22542_, _22418_);
  nand (_22544_, _22543_, _09012_);
  nor (_22545_, _22409_, _09012_);
  nor (_22546_, _22545_, _02987_);
  nand (_22547_, _22546_, _22544_);
  and (_22549_, _05394_, _02987_);
  nor (_22550_, _22549_, _09347_);
  nand (_22551_, _22550_, _22547_);
  and (_22552_, _05311_, _09347_);
  nor (_22553_, _22552_, _02986_);
  nand (_22554_, _22553_, _22551_);
  and (_22555_, _05394_, _02986_);
  nor (_22556_, _22555_, _13666_);
  and (_22557_, _22556_, _22554_);
  nor (_22558_, _22409_, _09005_);
  or (_22560_, _22558_, _22557_);
  nand (_22561_, _22560_, _07596_);
  nor (_22562_, _07596_, _05394_);
  nor (_22563_, _22562_, _02585_);
  and (_22564_, _22563_, _22561_);
  and (_22565_, _22409_, _02585_);
  or (_22566_, _22565_, _02874_);
  nor (_22567_, _22566_, _22564_);
  and (_22568_, _05395_, _02874_);
  or (_22569_, _22568_, _22567_);
  nand (_22571_, _22569_, _05325_);
  and (_22572_, _05311_, _02578_);
  nor (_22573_, _22572_, _03023_);
  nand (_22574_, _22573_, _22571_);
  and (_22575_, _06138_, _03023_);
  nor (_22576_, _22575_, _20391_);
  nand (_22577_, _22576_, _22574_);
  nor (_22578_, _09369_, _05394_);
  nor (_22579_, _22578_, _02576_);
  nand (_22580_, _22579_, _22577_);
  and (_22582_, _06138_, _02576_);
  nor (_22583_, _22582_, _09378_);
  nand (_22584_, _22583_, _22580_);
  nor (_22585_, _22409_, _09376_);
  nor (_22586_, _22585_, _02938_);
  nand (_22587_, _22586_, _22584_);
  nor (_22588_, _05394_, _02521_);
  or (_22589_, _22588_, _09380_);
  nand (_22590_, _22589_, _22587_);
  and (_22591_, _05311_, _02521_);
  nor (_22593_, _22591_, _09384_);
  nand (_22594_, _22593_, _22590_);
  and (_22595_, _22438_, _09384_);
  nor (_22596_, _22595_, _05562_);
  nand (_22597_, _22596_, _22594_);
  nor (_22598_, _05394_, _05322_);
  nor (_22599_, _22598_, _03014_);
  nand (_22600_, _22599_, _22597_);
  and (_22601_, _06138_, _03014_);
  nor (_22602_, _22601_, _07782_);
  and (_22603_, _22602_, _22600_);
  and (_22604_, _07782_, _05395_);
  or (_22605_, _22604_, _22603_);
  nand (_22606_, _22605_, _09401_);
  or (_22607_, _09405_, _09404_);
  and (_22608_, _22607_, _09424_);
  nor (_22609_, _22607_, _09424_);
  nor (_22610_, _22609_, _22608_);
  nor (_22611_, _22610_, _09401_);
  nor (_22612_, _22611_, _02937_);
  nand (_22614_, _22612_, _22606_);
  and (_22615_, _05394_, _02937_);
  nor (_22616_, _22615_, _02517_);
  nand (_22617_, _22616_, _22614_);
  and (_22618_, _05311_, _02517_);
  nor (_22619_, _22618_, _09000_);
  nand (_22620_, _22619_, _22617_);
  and (_22621_, _08190_, _05394_);
  and (_22622_, _22438_, _08880_);
  or (_22623_, _22622_, _22621_);
  and (_22625_, _22623_, _09000_);
  nor (_22626_, _22625_, _20808_);
  and (_22627_, _22626_, _22620_);
  or (_22628_, _22627_, _22417_);
  nand (_22629_, _22628_, _09450_);
  nor (_22630_, _09450_, _05394_);
  nor (_22631_, _22630_, _03021_);
  and (_22632_, _22631_, _22629_);
  and (_22633_, _06138_, _03021_);
  or (_22634_, _22633_, _03130_);
  nor (_22636_, _22634_, _22632_);
  and (_22637_, _05395_, _03130_);
  or (_22638_, _22637_, _22636_);
  nand (_22639_, _22638_, _02513_);
  and (_22640_, _05311_, _02512_);
  nor (_22641_, _22640_, _08994_);
  nand (_22642_, _22641_, _22639_);
  and (_22643_, _08880_, _05394_);
  and (_22644_, _22438_, _08190_);
  or (_22645_, _22644_, _22643_);
  and (_22647_, _22645_, _08994_);
  nor (_22648_, _22647_, _20466_);
  and (_22649_, _22648_, _22642_);
  or (_22650_, _22649_, _22416_);
  nand (_22651_, _22650_, _09475_);
  nor (_22652_, _09475_, _05394_);
  nor (_22653_, _22652_, _03020_);
  and (_22654_, _22653_, _22651_);
  and (_22655_, _06138_, _03020_);
  or (_22656_, _22655_, _03139_);
  nor (_22658_, _22656_, _22654_);
  and (_22659_, _05395_, _03139_);
  or (_22660_, _22659_, _22658_);
  nand (_22661_, _22660_, _19955_);
  and (_22662_, _05311_, _02533_);
  nor (_22663_, _22662_, _08875_);
  nand (_22664_, _22663_, _22661_);
  and (_22665_, _05394_, \oc8051_golden_model_1.PSW [7]);
  and (_22666_, _22438_, _07319_);
  or (_22667_, _22666_, _22665_);
  and (_22668_, _22667_, _08875_);
  nor (_22669_, _22668_, _09487_);
  and (_22670_, _22669_, _22664_);
  or (_22671_, _22670_, _22415_);
  nand (_22672_, _22671_, _07866_);
  nor (_22673_, _07866_, _05394_);
  nor (_22674_, _22673_, _03036_);
  nand (_22675_, _22674_, _22672_);
  and (_22676_, _06138_, _03036_);
  nor (_22677_, _22676_, _03127_);
  and (_22679_, _22677_, _22675_);
  and (_22680_, _05395_, _03127_);
  or (_22681_, _22680_, _22679_);
  nand (_22682_, _22681_, _19951_);
  and (_22683_, _05311_, _02538_);
  nor (_22684_, _22683_, _08864_);
  nand (_22685_, _22684_, _22682_);
  and (_22686_, _05394_, _07319_);
  and (_22687_, _22438_, \oc8051_golden_model_1.PSW [7]);
  or (_22688_, _22687_, _22686_);
  and (_22690_, _22688_, _08864_);
  nor (_22691_, _22690_, _09503_);
  and (_22692_, _22691_, _22685_);
  or (_22693_, _22692_, _22414_);
  nand (_22694_, _22693_, _08860_);
  nor (_22695_, _08860_, _05394_);
  nor (_22696_, _22695_, _08029_);
  nand (_22697_, _22696_, _22694_);
  and (_22698_, _22409_, _08029_);
  nor (_22699_, _22698_, _03148_);
  and (_22701_, _22699_, _22697_);
  nor (_22702_, _05490_, _10250_);
  or (_22703_, _22702_, _22701_);
  nand (_22704_, _22703_, _05792_);
  and (_22705_, _05311_, _02531_);
  nor (_22706_, _22705_, _03035_);
  nand (_22707_, _22706_, _22704_);
  and (_22708_, _22430_, _09709_);
  nor (_22709_, _09709_, _06138_);
  or (_22710_, _22709_, _03152_);
  or (_22712_, _22710_, _22708_);
  and (_22713_, _22712_, _08858_);
  and (_22714_, _22713_, _22707_);
  or (_22715_, _22714_, _22413_);
  nand (_22716_, _22715_, _08104_);
  nor (_22717_, _08104_, _05394_);
  nor (_22718_, _22717_, _08135_);
  nand (_22719_, _22718_, _22716_);
  and (_22720_, _22409_, _08135_);
  nor (_22721_, _22720_, _02897_);
  and (_22723_, _22721_, _22719_);
  nor (_22724_, _05490_, _02898_);
  or (_22725_, _22724_, _22723_);
  nand (_22726_, _22725_, _09728_);
  and (_22727_, _05311_, _02536_);
  nor (_22728_, _22727_, _02895_);
  nand (_22729_, _22728_, _22726_);
  and (_22730_, _09709_, _06139_);
  nor (_22731_, _22424_, _09709_);
  nor (_22732_, _22731_, _22730_);
  and (_22733_, _22732_, _02895_);
  nor (_22734_, _22733_, _09737_);
  nand (_22735_, _22734_, _22729_);
  nor (_22736_, _22409_, _09736_);
  nor (_22737_, _22736_, _03166_);
  and (_22738_, _22737_, _22735_);
  or (_22739_, _22738_, _22412_);
  nand (_22740_, _22739_, _09743_);
  nor (_22741_, _22419_, _09743_);
  nor (_22742_, _22741_, _04159_);
  nand (_22744_, _22742_, _22740_);
  and (_22745_, _05311_, _04159_);
  nor (_22746_, _22745_, _02500_);
  nand (_22747_, _22746_, _22744_);
  and (_22748_, _22732_, _02500_);
  nor (_22749_, _22748_, _09759_);
  nand (_22750_, _22749_, _22747_);
  nor (_22751_, _22409_, _09758_);
  nor (_22752_, _22751_, _03174_);
  and (_22753_, _22752_, _22750_);
  or (_22755_, _22753_, _22411_);
  nand (_22756_, _22755_, _09765_);
  nor (_22757_, _22419_, _09765_);
  nor (_22758_, _22757_, _19938_);
  nand (_22759_, _22758_, _22756_);
  and (_22760_, _19938_, _05311_);
  nor (_22761_, _22760_, _09777_);
  and (_22762_, _22761_, _22759_);
  or (_22763_, _22762_, _22410_);
  or (_22764_, _22763_, _34702_);
  or (_22766_, _34698_, \oc8051_golden_model_1.PC [7]);
  and (_22767_, _22766_, _36029_);
  and (_35246_, _22767_, _22764_);
  nor (_22768_, _02832_, _09770_);
  nor (_22769_, _02832_, _06195_);
  nor (_22770_, _08842_, \oc8051_golden_model_1.PC [8]);
  nor (_22771_, _22770_, _08849_);
  nor (_22772_, _22771_, _08858_);
  and (_22773_, _22771_, _08029_);
  nor (_22774_, _22771_, _08862_);
  nor (_22776_, _22771_, _08873_);
  nor (_22777_, _22771_, _09473_);
  and (_22778_, _09108_, _03021_);
  nor (_22779_, _22771_, _09448_);
  nor (_22780_, _09384_, _02521_);
  and (_22781_, _08917_, _02938_);
  nor (_22782_, _22771_, _09012_);
  nor (_22783_, _20340_, _08917_);
  not (_22784_, _09252_);
  and (_22785_, _08917_, _02887_);
  or (_22787_, _02947_, _05382_);
  nand (_22788_, _08917_, _02891_);
  nor (_22789_, _09186_, _09108_);
  nor (_22790_, _09112_, _09106_);
  nor (_22791_, _22790_, _09113_);
  not (_22792_, _22791_);
  and (_22793_, _22792_, _09186_);
  or (_22794_, _22793_, _22789_);
  and (_22795_, _22794_, _02952_);
  not (_22796_, _08917_);
  or (_22797_, _09198_, _22796_);
  nor (_22798_, _08967_, _08965_);
  nor (_22799_, _22798_, _08968_);
  nand (_22800_, _22799_, _09198_);
  and (_22801_, _22800_, _22797_);
  and (_22802_, _22801_, _10433_);
  nand (_22803_, _08917_, _02954_);
  nor (_22804_, _22771_, _09207_);
  and (_22805_, _22796_, _03825_);
  nor (_22806_, _03825_, \oc8051_golden_model_1.PC [8]);
  and (_22808_, _22806_, _09206_);
  or (_22809_, _22808_, _22805_);
  and (_22810_, _22809_, _09204_);
  and (_22811_, _22810_, _09203_);
  or (_22812_, _22811_, _22804_);
  and (_22813_, _22812_, _02558_);
  nor (_22814_, _22771_, _09203_);
  or (_22815_, _22814_, _02954_);
  or (_22816_, _22815_, _22813_);
  and (_22817_, _22816_, _22803_);
  or (_22819_, _22817_, _07452_);
  nand (_22820_, _22771_, _07452_);
  and (_22821_, _05387_, _02563_);
  and (_22822_, _22821_, _22820_);
  and (_22823_, _22822_, _22819_);
  or (_22824_, _22823_, _03818_);
  or (_22825_, _22824_, _22802_);
  nand (_22826_, _22771_, _03818_);
  and (_22827_, _22826_, _03821_);
  and (_22828_, _22827_, _22825_);
  or (_22830_, _22828_, _22795_);
  and (_22831_, _22830_, _09180_);
  nor (_22832_, _22771_, _09180_);
  or (_22833_, _22832_, _02891_);
  or (_22834_, _22833_, _22831_);
  and (_22835_, _22834_, _22788_);
  nor (_22836_, _22835_, _22787_);
  and (_22837_, _08917_, _02947_);
  nor (_22838_, _22837_, _09240_);
  not (_22839_, _22838_);
  nor (_22841_, _22839_, _22836_);
  nor (_22842_, _22771_, _09239_);
  nor (_22843_, _22842_, _02950_);
  not (_22844_, _22843_);
  nor (_22845_, _22844_, _22841_);
  and (_22846_, _08917_, _02950_);
  nor (_22847_, _22846_, _09249_);
  not (_22848_, _22847_);
  nor (_22849_, _22848_, _22845_);
  nor (_22850_, _22771_, _09247_);
  nor (_22852_, _22850_, _02887_);
  not (_22853_, _22852_);
  nor (_22854_, _22853_, _22849_);
  nor (_22855_, _22854_, _22785_);
  nor (_22856_, _22855_, _22784_);
  and (_22857_, _08917_, _02886_);
  nor (_22858_, _22857_, _09299_);
  not (_22859_, _22858_);
  nor (_22860_, _22859_, _22856_);
  and (_22861_, _09297_, _09108_);
  nor (_22862_, _22792_, _09297_);
  or (_22863_, _22862_, _22861_);
  nor (_22864_, _22863_, _09263_);
  nor (_22865_, _22864_, _22860_);
  nor (_22866_, _22865_, _03038_);
  nor (_22867_, _22791_, _09169_);
  and (_22868_, _09169_, _09109_);
  nor (_22869_, _22868_, _22867_);
  nor (_22870_, _22869_, _09172_);
  or (_22871_, _22870_, _02966_);
  nor (_22873_, _22871_, _22866_);
  nor (_22874_, _22792_, _09334_);
  and (_22875_, _09334_, _09108_);
  nor (_22876_, _22875_, _22874_);
  nor (_22877_, _22876_, _03377_);
  nor (_22878_, _22877_, _22873_);
  nor (_22879_, _22878_, _03025_);
  and (_22880_, _09325_, _09108_);
  and (_22881_, _22791_, _21083_);
  or (_22882_, _22881_, _22880_);
  and (_22884_, _22882_, _03025_);
  or (_22885_, _22884_, _22879_);
  and (_22886_, _22885_, _09306_);
  and (_22887_, _22771_, _09305_);
  or (_22888_, _22887_, _22886_);
  and (_22889_, _22888_, _02881_);
  and (_22890_, _08917_, _02880_);
  and (_22891_, _20340_, _02561_);
  not (_22892_, _22891_);
  nor (_22893_, _22892_, _22890_);
  not (_22895_, _22893_);
  nor (_22896_, _22895_, _22889_);
  nor (_22897_, _22896_, _22783_);
  nor (_22898_, _22897_, _20047_);
  or (_22899_, _22898_, _02987_);
  or (_22900_, _22899_, _22782_);
  and (_22901_, _08917_, _02987_);
  nor (_22902_, _22901_, _09347_);
  and (_22903_, _22902_, _22900_);
  or (_22904_, _22903_, _02986_);
  and (_22906_, _08917_, _02986_);
  nor (_22907_, _22906_, _13666_);
  and (_22908_, _22907_, _22904_);
  nor (_22909_, _22771_, _09005_);
  or (_22910_, _22909_, _22908_);
  and (_22911_, _22910_, _07596_);
  nor (_22912_, _08917_, _07596_);
  nor (_22913_, _22912_, _02585_);
  not (_22914_, _22913_);
  or (_22915_, _22914_, _22911_);
  and (_22917_, _22771_, _02585_);
  nor (_22918_, _22917_, _02874_);
  nand (_22919_, _22918_, _22915_);
  and (_22920_, _22796_, _02874_);
  nor (_22921_, _03023_, _02578_);
  not (_22922_, _22921_);
  nor (_22923_, _22922_, _22920_);
  nand (_22924_, _22923_, _22919_);
  and (_22925_, _09108_, _03023_);
  nor (_22926_, _22925_, _20391_);
  nand (_22927_, _22926_, _22924_);
  nor (_22928_, _09369_, _08917_);
  nor (_22929_, _22928_, _02576_);
  nand (_22930_, _22929_, _22927_);
  and (_22931_, _09108_, _02576_);
  nor (_22932_, _22931_, _09378_);
  nand (_22933_, _22932_, _22930_);
  nor (_22934_, _22771_, _09376_);
  nor (_22935_, _22934_, _02938_);
  and (_22936_, _22935_, _22933_);
  or (_22938_, _22936_, _22781_);
  nand (_22939_, _22938_, _22780_);
  and (_22940_, _22799_, _09384_);
  nor (_22941_, _22940_, _05562_);
  nand (_22942_, _22941_, _22939_);
  nor (_22943_, _08917_, _05322_);
  nor (_22944_, _22943_, _03014_);
  nand (_22945_, _22944_, _22942_);
  and (_22946_, _09108_, _03014_);
  nor (_22947_, _22946_, _07782_);
  and (_22949_, _22947_, _22945_);
  and (_22950_, _22796_, _07782_);
  or (_22951_, _22950_, _22949_);
  nand (_22952_, _22951_, _09401_);
  and (_22953_, _09426_, _09403_);
  nor (_22954_, _22953_, _09427_);
  nor (_22955_, _22954_, _09401_);
  nor (_22956_, _22955_, _02937_);
  nand (_22957_, _22956_, _22952_);
  and (_22958_, _08917_, _02937_);
  nor (_22960_, _22958_, _02517_);
  nand (_22961_, _22960_, _22957_);
  nand (_22962_, _22961_, _09442_);
  nor (_22963_, _22799_, _08190_);
  nor (_22964_, _08917_, _08880_);
  nor (_22965_, _22964_, _09442_);
  not (_22966_, _22965_);
  nor (_22967_, _22966_, _22963_);
  nor (_22968_, _22967_, _20808_);
  and (_22969_, _22968_, _22962_);
  or (_22971_, _22969_, _22779_);
  nand (_22972_, _22971_, _09450_);
  nor (_22973_, _08917_, _09450_);
  nor (_22974_, _22973_, _03021_);
  and (_22975_, _22974_, _22972_);
  or (_22976_, _22975_, _22778_);
  nand (_22977_, _22976_, _03131_);
  and (_22978_, _08917_, _03130_);
  nor (_22979_, _22978_, _02512_);
  nand (_22980_, _22979_, _22977_);
  nand (_22982_, _22980_, _09462_);
  and (_22983_, _08917_, _08880_);
  and (_22984_, _22799_, _08190_);
  or (_22985_, _22984_, _22983_);
  and (_22986_, _22985_, _08994_);
  nor (_22987_, _22986_, _20466_);
  and (_22988_, _22987_, _22982_);
  or (_22989_, _22988_, _22777_);
  nand (_22990_, _22989_, _09475_);
  nor (_22991_, _08917_, _09475_);
  nor (_22993_, _22991_, _03020_);
  nand (_22994_, _22993_, _22990_);
  and (_22995_, _09108_, _03020_);
  nor (_22996_, _22995_, _03139_);
  nand (_22997_, _22996_, _22994_);
  nor (_22998_, _08875_, _02533_);
  and (_22999_, _22796_, _03139_);
  not (_23000_, _22999_);
  and (_23001_, _23000_, _22998_);
  nand (_23002_, _23001_, _22997_);
  or (_23004_, _22799_, \oc8051_golden_model_1.PSW [7]);
  or (_23005_, _08917_, _07319_);
  and (_23006_, _23005_, _08875_);
  and (_23007_, _23006_, _23004_);
  nor (_23008_, _23007_, _09487_);
  and (_23009_, _23008_, _23002_);
  or (_23010_, _23009_, _22776_);
  nand (_23011_, _23010_, _07866_);
  nor (_23012_, _08917_, _07866_);
  nor (_23013_, _23012_, _03036_);
  and (_23015_, _23013_, _23011_);
  and (_23016_, _09108_, _03036_);
  or (_23017_, _23016_, _03127_);
  or (_23018_, _23017_, _23015_);
  nor (_23019_, _08864_, _02538_);
  and (_23020_, _22796_, _03127_);
  not (_23021_, _23020_);
  and (_23022_, _23021_, _23019_);
  nand (_23023_, _23022_, _23018_);
  nor (_23024_, _22799_, _07319_);
  nor (_23026_, _08917_, \oc8051_golden_model_1.PSW [7]);
  nor (_23027_, _23026_, _08865_);
  not (_23028_, _23027_);
  nor (_23029_, _23028_, _23024_);
  nor (_23030_, _23029_, _09503_);
  and (_23031_, _23030_, _23023_);
  or (_23032_, _23031_, _22774_);
  nand (_23033_, _23032_, _08860_);
  nor (_23034_, _08917_, _08860_);
  nor (_23035_, _23034_, _08029_);
  and (_23037_, _23035_, _23033_);
  or (_23038_, _23037_, _22773_);
  nand (_23039_, _23038_, _10250_);
  and (_23040_, _03817_, _03148_);
  nor (_23041_, _23040_, _02531_);
  nand (_23042_, _23041_, _23039_);
  nand (_23043_, _23042_, _03152_);
  and (_23044_, _22792_, _09709_);
  nor (_23045_, _09709_, _09108_);
  or (_23046_, _23045_, _03152_);
  or (_23048_, _23046_, _23044_);
  and (_23049_, _23048_, _08858_);
  and (_23050_, _23049_, _23043_);
  or (_23051_, _23050_, _22772_);
  nand (_23052_, _23051_, _08104_);
  nor (_23053_, _08917_, _08104_);
  nor (_23054_, _23053_, _08135_);
  and (_23055_, _23054_, _23052_);
  and (_23056_, _22771_, _08135_);
  or (_23057_, _23056_, _23055_);
  nand (_23059_, _23057_, _02898_);
  and (_23060_, _03817_, _02897_);
  nor (_23061_, _23060_, _02536_);
  nand (_23062_, _23061_, _23059_);
  nand (_23063_, _23062_, _02896_);
  and (_23064_, _09709_, _09109_);
  nor (_23065_, _22791_, _09709_);
  nor (_23066_, _23065_, _23064_);
  and (_23067_, _23066_, _02895_);
  nor (_23068_, _23067_, _09737_);
  nand (_23070_, _23068_, _23063_);
  nor (_23071_, _22771_, _09736_);
  nor (_23072_, _23071_, _03166_);
  nand (_23073_, _23072_, _23070_);
  and (_23074_, _08917_, _03166_);
  nor (_23075_, _23074_, _09744_);
  nand (_23076_, _23075_, _23073_);
  nor (_23077_, _22771_, _09743_);
  nor (_23078_, _23077_, _03004_);
  and (_23079_, _23078_, _23076_);
  or (_23081_, _23079_, _22769_);
  nor (_23082_, _02528_, _02500_);
  nand (_23083_, _23082_, _23081_);
  and (_23084_, _23066_, _02500_);
  nor (_23085_, _23084_, _09759_);
  nand (_23086_, _23085_, _23083_);
  nor (_23087_, _22771_, _09758_);
  nor (_23088_, _23087_, _03174_);
  nand (_23089_, _23088_, _23086_);
  and (_23090_, _08917_, _03174_);
  nor (_23092_, _23090_, _09766_);
  nand (_23093_, _23092_, _23089_);
  nor (_23094_, _22771_, _09765_);
  nor (_23095_, _23094_, _03006_);
  and (_23096_, _23095_, _23093_);
  or (_23097_, _23096_, _22768_);
  nor (_23098_, _09777_, _02526_);
  and (_23099_, _23098_, _23097_);
  and (_23100_, _22771_, _09777_);
  or (_23101_, _23100_, _23099_);
  or (_23103_, _23101_, _34702_);
  or (_23104_, _34698_, \oc8051_golden_model_1.PC [8]);
  and (_23105_, _23104_, _36029_);
  and (_35247_, _23105_, _23103_);
  nor (_23106_, _03671_, _09770_);
  nor (_23107_, _03671_, _06195_);
  nor (_23108_, _08849_, \oc8051_golden_model_1.PC [9]);
  nor (_23109_, _23108_, _08850_);
  nor (_23110_, _23109_, _08858_);
  nor (_23111_, _23109_, _08862_);
  and (_23112_, _09047_, _03036_);
  nor (_23113_, _23109_, _08873_);
  and (_23114_, _09047_, _03020_);
  nor (_23115_, _23109_, _09473_);
  and (_23116_, _09047_, _03021_);
  nor (_23117_, _23109_, _09448_);
  and (_23118_, _08913_, _02938_);
  nor (_23119_, _23109_, _09012_);
  and (_23120_, _08913_, _02954_);
  nor (_23121_, _23109_, _09207_);
  not (_23124_, _08913_);
  and (_23125_, _23124_, _03825_);
  nor (_23126_, _03825_, \oc8051_golden_model_1.PC [9]);
  and (_23127_, _23126_, _09206_);
  or (_23128_, _23127_, _23125_);
  and (_23129_, _23128_, _09204_);
  and (_23130_, _23129_, _09203_);
  or (_23131_, _23130_, _23121_);
  and (_23132_, _23131_, _02558_);
  nor (_23133_, _23109_, _09203_);
  nor (_23135_, _23133_, _02954_);
  not (_23136_, _23135_);
  nor (_23137_, _23136_, _23132_);
  nor (_23138_, _23137_, _23120_);
  nor (_23139_, _23138_, _07452_);
  and (_23140_, _23109_, _07452_);
  nor (_23141_, _23140_, _23139_);
  and (_23142_, _23141_, _22821_);
  and (_23143_, _09196_, _08913_);
  or (_23144_, _08915_, _08914_);
  not (_23145_, _23144_);
  nor (_23146_, _23145_, _08969_);
  and (_23147_, _23145_, _08969_);
  nor (_23148_, _23147_, _23146_);
  nor (_23149_, _23148_, _09196_);
  or (_23150_, _23149_, _23143_);
  nor (_23151_, _23150_, _05387_);
  nor (_23152_, _23151_, _23142_);
  nor (_23153_, _23152_, _03818_);
  not (_23154_, _23109_);
  and (_23157_, _23154_, _03818_);
  or (_23158_, _23157_, _02952_);
  nor (_23159_, _23158_, _23153_);
  nor (_23160_, _09113_, _09110_);
  and (_23161_, _23160_, _09051_);
  nor (_23162_, _23160_, _09051_);
  nor (_23163_, _23162_, _23161_);
  and (_23164_, _23163_, _09186_);
  nor (_23165_, _09186_, _09047_);
  nor (_23166_, _23165_, _23164_);
  and (_23168_, _23166_, _02952_);
  or (_23169_, _23168_, _23159_);
  nor (_23170_, _23169_, _21709_);
  nor (_23171_, _23109_, _09180_);
  nor (_23172_, _23171_, _02891_);
  not (_23173_, _23172_);
  nor (_23174_, _23173_, _23170_);
  and (_23175_, _08913_, _02891_);
  or (_23176_, _23175_, _05382_);
  nor (_23177_, _23176_, _23174_);
  nor (_23178_, _23177_, _02947_);
  and (_23179_, _08913_, _02947_);
  nor (_23180_, _23179_, _09240_);
  not (_23181_, _23180_);
  nor (_23182_, _23181_, _23178_);
  nor (_23183_, _23109_, _09239_);
  nor (_23184_, _23183_, _02950_);
  not (_23185_, _23184_);
  nor (_23186_, _23185_, _23182_);
  and (_23187_, _08913_, _02950_);
  nor (_23190_, _23187_, _09249_);
  not (_23191_, _23190_);
  nor (_23192_, _23191_, _23186_);
  nor (_23193_, _23109_, _09247_);
  nor (_23194_, _23193_, _02887_);
  not (_23195_, _23194_);
  nor (_23196_, _23195_, _23192_);
  and (_23197_, _08913_, _02887_);
  or (_23198_, _23197_, _09251_);
  nor (_23199_, _23198_, _23196_);
  nor (_23201_, _23199_, _02886_);
  and (_23202_, _08913_, _02886_);
  nor (_23203_, _23202_, _09299_);
  not (_23204_, _23203_);
  nor (_23205_, _23204_, _23201_);
  and (_23206_, _09297_, _09047_);
  nor (_23207_, _23163_, _09297_);
  or (_23208_, _23207_, _23206_);
  nor (_23209_, _23208_, _09263_);
  nor (_23210_, _23209_, _23205_);
  nor (_23211_, _23210_, _03038_);
  and (_23212_, _09169_, _09048_);
  not (_23213_, _23163_);
  nor (_23214_, _23213_, _09169_);
  nor (_23215_, _23214_, _23212_);
  nor (_23216_, _23215_, _09172_);
  or (_23217_, _23216_, _02966_);
  nor (_23218_, _23217_, _23211_);
  and (_23219_, _09334_, _09047_);
  nor (_23220_, _23163_, _09334_);
  nor (_23223_, _23220_, _23219_);
  nor (_23224_, _23223_, _03377_);
  nor (_23225_, _23224_, _23218_);
  nor (_23226_, _23225_, _03025_);
  and (_23227_, _09325_, _09047_);
  nor (_23228_, _23163_, _09325_);
  or (_23229_, _23228_, _23227_);
  and (_23230_, _23229_, _03025_);
  or (_23231_, _23230_, _23226_);
  and (_23232_, _23231_, _09306_);
  and (_23234_, _23109_, _09305_);
  or (_23235_, _23234_, _23232_);
  nor (_23236_, _23235_, _02880_);
  and (_23237_, _23124_, _02880_);
  nor (_23238_, _23237_, _22892_);
  not (_23239_, _23238_);
  or (_23240_, _23239_, _23236_);
  nor (_23241_, _20340_, _23124_);
  nor (_23242_, _23241_, _20047_);
  and (_23243_, _23242_, _23240_);
  or (_23244_, _23243_, _23119_);
  and (_23245_, _23244_, _09346_);
  nand (_23246_, _23124_, _02987_);
  nand (_23247_, _23246_, _09348_);
  or (_23248_, _23247_, _23245_);
  and (_23249_, _08913_, _02986_);
  nor (_23250_, _23249_, _13666_);
  and (_23251_, _23250_, _23248_);
  nor (_23252_, _23109_, _09005_);
  or (_23253_, _23252_, _23251_);
  and (_23256_, _23253_, _07596_);
  nor (_23257_, _08913_, _07596_);
  nor (_23258_, _23257_, _02585_);
  not (_23259_, _23258_);
  or (_23260_, _23259_, _23256_);
  and (_23261_, _23109_, _02585_);
  nor (_23262_, _23261_, _02874_);
  nand (_23263_, _23262_, _23260_);
  and (_23264_, _23124_, _02874_);
  nor (_23265_, _23264_, _22922_);
  nand (_23267_, _23265_, _23263_);
  and (_23268_, _09047_, _03023_);
  nor (_23269_, _23268_, _20391_);
  nand (_23270_, _23269_, _23267_);
  nor (_23271_, _09369_, _08913_);
  nor (_23272_, _23271_, _02576_);
  nand (_23273_, _23272_, _23270_);
  and (_23274_, _09047_, _02576_);
  nor (_23275_, _23274_, _09378_);
  nand (_23276_, _23275_, _23273_);
  nor (_23277_, _23109_, _09376_);
  nor (_23278_, _23277_, _02938_);
  and (_23279_, _23278_, _23276_);
  or (_23280_, _23279_, _23118_);
  nand (_23281_, _23280_, _22780_);
  nor (_23282_, _23148_, _09385_);
  nor (_23283_, _23282_, _05562_);
  nand (_23284_, _23283_, _23281_);
  nor (_23285_, _08913_, _05322_);
  nor (_23286_, _23285_, _03014_);
  nand (_23289_, _23286_, _23284_);
  and (_23290_, _09047_, _03014_);
  nor (_23291_, _23290_, _07782_);
  and (_23292_, _23291_, _23289_);
  and (_23293_, _23124_, _07782_);
  or (_23294_, _23293_, _23292_);
  nand (_23295_, _23294_, _09401_);
  nor (_23296_, _09427_, \oc8051_golden_model_1.DPH [1]);
  nor (_23297_, _23296_, _09428_);
  nor (_23298_, _23297_, _09401_);
  nor (_23300_, _23298_, _02937_);
  nand (_23301_, _23300_, _23295_);
  and (_23302_, _08913_, _02937_);
  nor (_23303_, _23302_, _02517_);
  nand (_23304_, _23303_, _23301_);
  nand (_23305_, _23304_, _09442_);
  and (_23306_, _08913_, _08190_);
  nor (_23307_, _23148_, _08190_);
  or (_23308_, _23307_, _23306_);
  and (_23309_, _23308_, _09000_);
  nor (_23310_, _23309_, _20808_);
  and (_23311_, _23310_, _23305_);
  or (_23312_, _23311_, _23117_);
  nand (_23313_, _23312_, _09450_);
  nor (_23314_, _08913_, _09450_);
  nor (_23315_, _23314_, _03021_);
  and (_23316_, _23315_, _23313_);
  or (_23317_, _23316_, _23116_);
  nand (_23318_, _23317_, _03131_);
  and (_23319_, _08913_, _03130_);
  nor (_23322_, _23319_, _02512_);
  nand (_23323_, _23322_, _23318_);
  nand (_23324_, _23323_, _09462_);
  and (_23325_, _23148_, _08190_);
  nor (_23326_, _08913_, _08190_);
  nor (_23327_, _23326_, _09462_);
  not (_23328_, _23327_);
  nor (_23329_, _23328_, _23325_);
  nor (_23330_, _23329_, _20466_);
  and (_23331_, _23330_, _23324_);
  or (_23333_, _23331_, _23115_);
  nand (_23334_, _23333_, _09475_);
  nor (_23335_, _08913_, _09475_);
  nor (_23336_, _23335_, _03020_);
  and (_23337_, _23336_, _23334_);
  or (_23338_, _23337_, _23114_);
  nand (_23339_, _23338_, _03140_);
  and (_23340_, _08913_, _03139_);
  nor (_23341_, _23340_, _02533_);
  nand (_23342_, _23341_, _23339_);
  nand (_23344_, _23342_, _08876_);
  and (_23345_, _08913_, \oc8051_golden_model_1.PSW [7]);
  nor (_23346_, _23148_, \oc8051_golden_model_1.PSW [7]);
  or (_23347_, _23346_, _23345_);
  and (_23348_, _23347_, _08875_);
  nor (_23349_, _23348_, _09487_);
  and (_23350_, _23349_, _23344_);
  or (_23351_, _23350_, _23113_);
  nand (_23352_, _23351_, _07866_);
  nor (_23353_, _08913_, _07866_);
  nor (_23355_, _23353_, _03036_);
  and (_23356_, _23355_, _23352_);
  or (_23357_, _23356_, _23112_);
  nand (_23358_, _23357_, _05786_);
  and (_23359_, _08913_, _03127_);
  nor (_23360_, _23359_, _02538_);
  nand (_23361_, _23360_, _23358_);
  nand (_23362_, _23361_, _08865_);
  and (_23363_, _08913_, _07319_);
  nor (_23364_, _23148_, _07319_);
  or (_23366_, _23364_, _23363_);
  and (_23367_, _23366_, _08864_);
  nor (_23368_, _23367_, _09503_);
  and (_23369_, _23368_, _23362_);
  or (_23370_, _23369_, _23111_);
  nand (_23371_, _23370_, _08860_);
  nor (_23372_, _08913_, _08860_);
  nor (_23373_, _23372_, _08029_);
  nand (_23374_, _23373_, _23371_);
  and (_23375_, _23109_, _08029_);
  nor (_23377_, _23375_, _03148_);
  nand (_23378_, _23377_, _23374_);
  nor (_23379_, _03035_, _02531_);
  not (_23380_, _23379_);
  and (_23381_, _04038_, _03148_);
  nor (_23382_, _23381_, _23380_);
  nand (_23383_, _23382_, _23378_);
  nor (_23384_, _09709_, _09047_);
  and (_23385_, _23163_, _09709_);
  or (_23386_, _23385_, _03152_);
  or (_23388_, _23386_, _23384_);
  and (_23389_, _23388_, _08858_);
  and (_23390_, _23389_, _23383_);
  or (_23391_, _23390_, _23110_);
  nand (_23392_, _23391_, _08104_);
  nor (_23393_, _08913_, _08104_);
  nor (_23394_, _23393_, _08135_);
  nand (_23395_, _23394_, _23392_);
  and (_23396_, _23109_, _08135_);
  nor (_23397_, _23396_, _02897_);
  nand (_23399_, _23397_, _23395_);
  and (_23400_, _04038_, _02897_);
  nor (_23401_, _02895_, _02536_);
  not (_23402_, _23401_);
  nor (_23403_, _23402_, _23400_);
  nand (_23404_, _23403_, _23399_);
  nor (_23405_, _23213_, _09709_);
  and (_23406_, _09709_, _09048_);
  nor (_23407_, _23406_, _23405_);
  and (_23408_, _23407_, _02895_);
  nor (_23410_, _23408_, _09737_);
  nand (_23411_, _23410_, _23404_);
  nor (_23412_, _23109_, _09736_);
  nor (_23413_, _23412_, _03166_);
  nand (_23414_, _23413_, _23411_);
  and (_23415_, _08913_, _03166_);
  nor (_23416_, _23415_, _09744_);
  nand (_23417_, _23416_, _23414_);
  nor (_23418_, _23109_, _09743_);
  nor (_23419_, _23418_, _03004_);
  and (_23421_, _23419_, _23417_);
  or (_23422_, _23421_, _23107_);
  nand (_23423_, _23422_, _23082_);
  and (_23424_, _23407_, _02500_);
  nor (_23425_, _23424_, _09759_);
  nand (_23426_, _23425_, _23423_);
  nor (_23427_, _23109_, _09758_);
  nor (_23428_, _23427_, _03174_);
  nand (_23429_, _23428_, _23426_);
  and (_23430_, _08913_, _03174_);
  nor (_23432_, _23430_, _09766_);
  nand (_23433_, _23432_, _23429_);
  nor (_23434_, _23109_, _09765_);
  nor (_23435_, _23434_, _03006_);
  and (_23436_, _23435_, _23433_);
  or (_23437_, _23436_, _23106_);
  and (_23438_, _23437_, _23098_);
  and (_23439_, _23109_, _09777_);
  or (_23440_, _23439_, _23438_);
  or (_23441_, _23440_, _34702_);
  or (_23443_, _34698_, \oc8051_golden_model_1.PC [9]);
  and (_23444_, _23443_, _36029_);
  and (_35249_, _23444_, _23441_);
  nor (_23445_, _08850_, \oc8051_golden_model_1.PC [10]);
  nor (_23446_, _23445_, _08843_);
  or (_23447_, _23446_, _09758_);
  not (_23448_, _23446_);
  nand (_23449_, _23448_, _08135_);
  nand (_23450_, _23448_, _08029_);
  nand (_23451_, _09040_, _03036_);
  nand (_23453_, _09040_, _03020_);
  nand (_23454_, _09040_, _03021_);
  nor (_23455_, _09000_, _02517_);
  or (_23456_, _08908_, _09809_);
  or (_23457_, _20340_, _08908_);
  or (_23458_, _23446_, _09239_);
  nor (_23459_, _23448_, _09234_);
  nor (_23460_, _09117_, _09114_);
  not (_23461_, _23460_);
  and (_23462_, _23461_, _09043_);
  nor (_23464_, _23461_, _09043_);
  nor (_23465_, _23464_, _23462_);
  and (_23466_, _23465_, _09186_);
  nor (_23467_, _09186_, _09040_);
  or (_23468_, _23467_, _23466_);
  and (_23469_, _23468_, _02952_);
  and (_23470_, _09196_, _08908_);
  nor (_23471_, _08972_, _08911_);
  nor (_23472_, _23471_, _08974_);
  and (_23473_, _23472_, _09198_);
  or (_23475_, _23473_, _05387_);
  or (_23476_, _23475_, _23470_);
  nor (_23477_, _23448_, _09208_);
  and (_23478_, _08908_, _03825_);
  and (_23479_, _03826_, \oc8051_golden_model_1.PC [10]);
  and (_23480_, _23479_, _09206_);
  or (_23481_, _23480_, _23478_);
  and (_23482_, _23481_, _09204_);
  or (_23483_, _23482_, _03824_);
  and (_23484_, _23483_, _09203_);
  or (_23486_, _23484_, _02954_);
  or (_23487_, _23486_, _23477_);
  or (_23488_, _08908_, _07433_);
  and (_23489_, _23488_, _09202_);
  and (_23490_, _23489_, _23487_);
  nand (_23491_, _23446_, _07452_);
  nand (_23492_, _23491_, _22821_);
  or (_23493_, _23492_, _23490_);
  and (_23494_, _23493_, _09228_);
  and (_23495_, _23494_, _23476_);
  or (_23497_, _23495_, _23469_);
  and (_23498_, _23497_, _09180_);
  or (_23499_, _23498_, _23459_);
  and (_23500_, _23499_, _02951_);
  and (_23501_, _08908_, _09918_);
  nor (_23502_, _23501_, _05382_);
  nand (_23503_, _23502_, _09239_);
  or (_23504_, _23503_, _23500_);
  and (_23505_, _23504_, _23458_);
  or (_23506_, _23505_, _02950_);
  or (_23508_, _08908_, _02959_);
  and (_23509_, _23508_, _09247_);
  and (_23510_, _23509_, _23506_);
  nor (_23511_, _23448_, _09247_);
  or (_23512_, _23511_, _23510_);
  and (_23513_, _23512_, _02888_);
  and (_23514_, _08908_, _02887_);
  or (_23515_, _23514_, _09251_);
  or (_23516_, _23515_, _23513_);
  and (_23517_, _23516_, _03947_);
  nand (_23519_, _08908_, _02886_);
  nand (_23520_, _23519_, _09263_);
  or (_23521_, _23520_, _23517_);
  or (_23522_, _23465_, _09297_);
  nand (_23523_, _09297_, _09040_);
  and (_23524_, _23523_, _23522_);
  or (_23525_, _23524_, _09263_);
  and (_23526_, _23525_, _23521_);
  or (_23527_, _23526_, _03038_);
  or (_23528_, _23465_, _09169_);
  nand (_23530_, _09169_, _09040_);
  and (_23531_, _23530_, _23528_);
  or (_23532_, _23531_, _09172_);
  and (_23533_, _23532_, _03377_);
  and (_23534_, _23533_, _23527_);
  nand (_23535_, _09334_, _09040_);
  or (_23536_, _23465_, _09334_);
  and (_23537_, _23536_, _02966_);
  and (_23538_, _23537_, _23535_);
  or (_23539_, _23538_, _23534_);
  and (_23541_, _23539_, _10029_);
  or (_23542_, _23465_, _09325_);
  nand (_23543_, _09325_, _09040_);
  and (_23544_, _23543_, _03025_);
  and (_23545_, _23544_, _23542_);
  or (_23546_, _23545_, _09305_);
  or (_23547_, _23546_, _23541_);
  nand (_23548_, _23448_, _09305_);
  and (_23549_, _23548_, _02881_);
  and (_23550_, _23549_, _23547_);
  or (_23552_, _23550_, _22892_);
  and (_23553_, _23552_, _23457_);
  nand (_23554_, _08908_, _02880_);
  nand (_23555_, _23554_, _09012_);
  or (_23556_, _23555_, _23553_);
  or (_23557_, _23446_, _09012_);
  and (_23558_, _23557_, _09346_);
  nand (_23559_, _23558_, _23556_);
  nand (_23560_, _23559_, _09348_);
  and (_23561_, _23560_, _23456_);
  nand (_23563_, _08908_, _02987_);
  nand (_23564_, _23563_, _09005_);
  or (_23565_, _23564_, _23561_);
  or (_23566_, _23446_, _09005_);
  and (_23567_, _23566_, _07596_);
  and (_23568_, _23567_, _23565_);
  and (_23569_, _08908_, _07597_);
  or (_23570_, _23569_, _02585_);
  or (_23571_, _23570_, _23568_);
  nand (_23572_, _23448_, _02585_);
  and (_23574_, _23572_, _02875_);
  and (_23575_, _23574_, _23571_);
  nand (_23576_, _08908_, _02874_);
  nand (_23577_, _23576_, _22921_);
  or (_23578_, _23577_, _23575_);
  nand (_23579_, _09040_, _03023_);
  and (_23580_, _23579_, _09369_);
  and (_23581_, _23580_, _23578_);
  and (_23582_, _20391_, _08908_);
  or (_23583_, _23582_, _02576_);
  or (_23585_, _23583_, _23581_);
  nand (_23586_, _09040_, _02576_);
  and (_23587_, _23586_, _09376_);
  and (_23588_, _23587_, _23585_);
  nor (_23589_, _23448_, _09376_);
  or (_23590_, _23589_, _23588_);
  and (_23591_, _23590_, _09801_);
  nand (_23592_, _08908_, _02938_);
  nand (_23593_, _23592_, _22780_);
  or (_23594_, _23593_, _23591_);
  or (_23596_, _23472_, _09385_);
  and (_23597_, _23596_, _05322_);
  and (_23598_, _23597_, _23594_);
  and (_23599_, _08908_, _05562_);
  or (_23600_, _23599_, _03014_);
  or (_23601_, _23600_, _23598_);
  nand (_23602_, _09040_, _03014_);
  and (_23603_, _23602_, _07783_);
  and (_23604_, _23603_, _23601_);
  and (_23605_, _08908_, _07782_);
  or (_23607_, _23605_, _09400_);
  or (_23608_, _23607_, _23604_);
  nor (_23609_, _09428_, \oc8051_golden_model_1.DPH [2]);
  nor (_23610_, _23609_, _09429_);
  nor (_23611_, _23610_, _09401_);
  nor (_23612_, _23611_, _02937_);
  and (_23613_, _23612_, _23608_);
  and (_23614_, _08908_, _02937_);
  or (_23615_, _23614_, _23613_);
  and (_23616_, _23615_, _23455_);
  or (_23618_, _23472_, _08190_);
  or (_23619_, _08908_, _08880_);
  and (_23620_, _23619_, _09000_);
  and (_23621_, _23620_, _23618_);
  or (_23622_, _23621_, _20808_);
  or (_23623_, _23622_, _23616_);
  or (_23624_, _23446_, _09448_);
  and (_23625_, _23624_, _09450_);
  and (_23626_, _23625_, _23623_);
  and (_23627_, _08908_, _09451_);
  or (_23629_, _23627_, _03021_);
  or (_23630_, _23629_, _23626_);
  and (_23631_, _23630_, _23454_);
  or (_23632_, _23631_, _03130_);
  or (_23633_, _08908_, _03131_);
  nor (_23634_, _08994_, _02512_);
  and (_23635_, _23634_, _23633_);
  and (_23636_, _23635_, _23632_);
  or (_23637_, _23472_, _08880_);
  or (_23638_, _08908_, _08190_);
  and (_23640_, _23638_, _08994_);
  and (_23641_, _23640_, _23637_);
  or (_23642_, _23641_, _20466_);
  or (_23643_, _23642_, _23636_);
  or (_23644_, _23446_, _09473_);
  and (_23645_, _23644_, _09475_);
  and (_23646_, _23645_, _23643_);
  and (_23647_, _08908_, _09476_);
  or (_23648_, _23647_, _03020_);
  or (_23649_, _23648_, _23646_);
  and (_23651_, _23649_, _23453_);
  or (_23652_, _23651_, _03139_);
  or (_23653_, _08908_, _03140_);
  and (_23654_, _23653_, _22998_);
  and (_23655_, _23654_, _23652_);
  or (_23656_, _23472_, \oc8051_golden_model_1.PSW [7]);
  or (_23657_, _08908_, _07319_);
  and (_23658_, _23657_, _08875_);
  and (_23659_, _23658_, _23656_);
  or (_23660_, _23659_, _09487_);
  or (_23662_, _23660_, _23655_);
  or (_23663_, _23446_, _08873_);
  and (_23664_, _23663_, _07866_);
  and (_23665_, _23664_, _23662_);
  and (_23666_, _08908_, _07867_);
  or (_23667_, _23666_, _03036_);
  or (_23668_, _23667_, _23665_);
  and (_23669_, _23668_, _23451_);
  or (_23670_, _23669_, _03127_);
  or (_23671_, _08908_, _05786_);
  and (_23673_, _23671_, _23019_);
  and (_23674_, _23673_, _23670_);
  or (_23675_, _23472_, _07319_);
  or (_23676_, _08908_, \oc8051_golden_model_1.PSW [7]);
  and (_23677_, _23676_, _08864_);
  and (_23678_, _23677_, _23675_);
  or (_23679_, _23678_, _09503_);
  or (_23680_, _23679_, _23674_);
  or (_23681_, _23446_, _08862_);
  and (_23682_, _23681_, _08860_);
  and (_23684_, _23682_, _23680_);
  and (_23685_, _08908_, _08861_);
  or (_23686_, _23685_, _08029_);
  or (_23687_, _23686_, _23684_);
  and (_23688_, _23687_, _23450_);
  or (_23689_, _23688_, _03148_);
  nand (_23690_, _04440_, _03148_);
  and (_23691_, _23690_, _23379_);
  and (_23692_, _23691_, _23689_);
  or (_23693_, _23465_, _09710_);
  or (_23695_, _09709_, _09038_);
  and (_23696_, _23695_, _03035_);
  and (_23697_, _23696_, _23693_);
  or (_23698_, _23697_, _09524_);
  or (_23699_, _23698_, _23692_);
  or (_23700_, _23446_, _08858_);
  and (_23701_, _23700_, _08104_);
  and (_23702_, _23701_, _23699_);
  and (_23703_, _08908_, _08105_);
  or (_23704_, _23703_, _08135_);
  or (_23706_, _23704_, _23702_);
  and (_23707_, _23706_, _23449_);
  or (_23708_, _23707_, _02897_);
  nand (_23709_, _04440_, _02897_);
  and (_23710_, _23709_, _23401_);
  and (_23711_, _23710_, _23708_);
  nand (_23712_, _09709_, _09040_);
  or (_23713_, _23465_, _09709_);
  and (_23714_, _23713_, _23712_);
  and (_23715_, _23714_, _02895_);
  or (_23717_, _23715_, _09737_);
  or (_23718_, _23717_, _23711_);
  or (_23719_, _23446_, _09736_);
  and (_23720_, _23719_, _23718_);
  or (_23721_, _23720_, _03166_);
  or (_23722_, _08908_, _03563_);
  and (_23723_, _23722_, _09743_);
  and (_23724_, _23723_, _23721_);
  nor (_23725_, _23448_, _09743_);
  or (_23726_, _23725_, _03004_);
  or (_23728_, _23726_, _23724_);
  nand (_23729_, _03260_, _03004_);
  and (_23730_, _23729_, _23082_);
  and (_23731_, _23730_, _23728_);
  and (_23732_, _23714_, _02500_);
  or (_23733_, _23732_, _09759_);
  or (_23734_, _23733_, _23731_);
  and (_23735_, _23734_, _23447_);
  or (_23736_, _23735_, _03174_);
  or (_23737_, _08908_, _03178_);
  and (_23739_, _23737_, _09765_);
  and (_23740_, _23739_, _23736_);
  nor (_23741_, _23448_, _09765_);
  or (_23742_, _23741_, _03006_);
  or (_23743_, _23742_, _23740_);
  nand (_23744_, _03260_, _03006_);
  and (_23745_, _23744_, _23098_);
  and (_23746_, _23745_, _23743_);
  and (_23747_, _23446_, _09777_);
  or (_23748_, _23747_, _23746_);
  or (_23750_, _23748_, _34702_);
  or (_23751_, _34698_, \oc8051_golden_model_1.PC [10]);
  and (_23752_, _23751_, _36029_);
  and (_35250_, _23752_, _23750_);
  nor (_23753_, _08843_, _08901_);
  and (_23754_, _08843_, _08901_);
  or (_23755_, _23754_, _23753_);
  nor (_23756_, _23755_, _08858_);
  nor (_23757_, _23755_, _08862_);
  nor (_23758_, _08904_, _08866_);
  or (_23760_, _23758_, _08864_);
  nor (_23761_, _23755_, _08873_);
  and (_23762_, _08904_, _08880_);
  or (_23763_, _08905_, _08906_);
  and (_23764_, _23763_, _08975_);
  nor (_23765_, _23763_, _08975_);
  nor (_23766_, _23765_, _23764_);
  and (_23767_, _23766_, _08190_);
  or (_23768_, _23767_, _23762_);
  and (_23769_, _23768_, _08994_);
  nor (_23771_, _23755_, _09448_);
  nor (_23772_, _08904_, _05322_);
  and (_23773_, _09032_, _02576_);
  nor (_23774_, _23755_, _09005_);
  not (_23775_, _09349_);
  not (_23776_, _23755_);
  nor (_23777_, _23776_, _09012_);
  and (_23778_, _09325_, _09032_);
  nor (_23779_, _23462_, _09041_);
  and (_23780_, _23779_, _09036_);
  nor (_23782_, _23779_, _09036_);
  nor (_23783_, _23782_, _23780_);
  nor (_23784_, _23783_, _09325_);
  or (_23785_, _23784_, _23778_);
  and (_23786_, _23785_, _03025_);
  and (_23787_, _09169_, _09033_);
  not (_23788_, _23783_);
  nor (_23789_, _23788_, _09169_);
  nor (_23790_, _23789_, _23787_);
  nor (_23791_, _23790_, _09172_);
  and (_23793_, _08904_, _02950_);
  nor (_23794_, _09177_, _08904_);
  nor (_23795_, _09186_, _09032_);
  and (_23796_, _23783_, _09186_);
  or (_23797_, _23796_, _03821_);
  or (_23798_, _23797_, _23795_);
  and (_23799_, _09196_, _08904_);
  and (_23800_, _23766_, _09198_);
  or (_23801_, _23800_, _05387_);
  nor (_23802_, _23801_, _23799_);
  not (_23804_, _09228_);
  nor (_23805_, _23755_, _09208_);
  not (_23806_, _23805_);
  nor (_23807_, _09213_, _08904_);
  and (_23808_, _02558_, _08901_);
  nor (_23809_, _07442_, _03825_);
  and (_23810_, _23809_, _23808_);
  and (_23811_, _23810_, _09206_);
  nor (_23812_, _23811_, _23807_);
  nor (_23813_, _23812_, _20635_);
  nor (_23815_, _23813_, _02954_);
  and (_23816_, _23815_, _23806_);
  and (_23817_, _08904_, _02954_);
  or (_23818_, _23817_, _23816_);
  and (_23819_, _23818_, _09202_);
  and (_23820_, _23755_, _07452_);
  or (_23821_, _23820_, _23819_);
  and (_23822_, _23821_, _02563_);
  not (_23823_, _08904_);
  nor (_23824_, _23823_, _02563_);
  nor (_23826_, _23824_, _10433_);
  not (_23827_, _23826_);
  nor (_23828_, _23827_, _23822_);
  or (_23829_, _23828_, _23804_);
  or (_23830_, _23829_, _23802_);
  and (_23831_, _23830_, _23798_);
  or (_23832_, _23831_, _21709_);
  or (_23833_, _23776_, _09234_);
  and (_23834_, _23833_, _09177_);
  and (_23835_, _23834_, _23832_);
  nor (_23837_, _23835_, _23794_);
  nor (_23838_, _23837_, _09240_);
  nor (_23839_, _23755_, _09239_);
  nor (_23840_, _23839_, _02950_);
  not (_23841_, _23840_);
  nor (_23842_, _23841_, _23838_);
  nor (_23843_, _23842_, _23793_);
  nor (_23844_, _23843_, _09249_);
  nor (_23845_, _23776_, _09247_);
  nor (_23846_, _23845_, _09254_);
  not (_23848_, _23846_);
  nor (_23849_, _23848_, _23844_);
  nor (_23850_, _09253_, _08904_);
  or (_23851_, _23850_, _09299_);
  or (_23852_, _23851_, _23849_);
  and (_23853_, _09297_, _09033_);
  nor (_23854_, _23788_, _09297_);
  or (_23855_, _23854_, _09263_);
  or (_23856_, _23855_, _23853_);
  and (_23857_, _23856_, _09172_);
  and (_23859_, _23857_, _23852_);
  nor (_23860_, _23859_, _23791_);
  and (_23861_, _23860_, _03377_);
  nor (_23862_, _23783_, _09334_);
  and (_23863_, _09334_, _09032_);
  or (_23864_, _23863_, _23862_);
  and (_23865_, _23864_, _02966_);
  or (_23866_, _23865_, _23861_);
  and (_23867_, _23866_, _10029_);
  nor (_23868_, _23867_, _23786_);
  nor (_23870_, _23868_, _09305_);
  and (_23871_, _23755_, _09305_);
  not (_23872_, _23871_);
  and (_23873_, _23872_, _09314_);
  not (_23874_, _23873_);
  nor (_23875_, _23874_, _23870_);
  nor (_23876_, _09314_, _08904_);
  nor (_23877_, _23876_, _20047_);
  not (_23878_, _23877_);
  nor (_23879_, _23878_, _23875_);
  nor (_23881_, _23879_, _23777_);
  nor (_23882_, _23881_, _23775_);
  nor (_23883_, _09349_, _23823_);
  nor (_23884_, _23883_, _13666_);
  not (_23885_, _23884_);
  nor (_23886_, _23885_, _23882_);
  nor (_23887_, _23886_, _23774_);
  nor (_23888_, _23887_, _07597_);
  nor (_23889_, _08904_, _07596_);
  nor (_23890_, _23889_, _02585_);
  not (_23892_, _23890_);
  nor (_23893_, _23892_, _23888_);
  and (_23894_, _23755_, _02585_);
  nor (_23895_, _23894_, _09362_);
  not (_23896_, _23895_);
  nor (_23897_, _23896_, _23893_);
  nor (_23898_, _09361_, _08904_);
  nor (_23899_, _23898_, _03023_);
  not (_23900_, _23899_);
  nor (_23901_, _23900_, _23897_);
  and (_23903_, _09032_, _03023_);
  nor (_23904_, _23903_, _20391_);
  not (_23905_, _23904_);
  or (_23906_, _23905_, _23901_);
  nor (_23907_, _09369_, _08904_);
  nor (_23908_, _23907_, _02576_);
  and (_23909_, _23908_, _23906_);
  or (_23910_, _23909_, _23773_);
  and (_23911_, _23910_, _09376_);
  nor (_23912_, _23776_, _09376_);
  nor (_23914_, _23912_, _09381_);
  not (_23915_, _23914_);
  or (_23916_, _23915_, _23911_);
  nor (_23917_, _09380_, _08904_);
  nor (_23918_, _23917_, _09384_);
  nand (_23919_, _23918_, _23916_);
  and (_23920_, _23766_, _09384_);
  nor (_23921_, _23920_, _05562_);
  and (_23922_, _23921_, _23919_);
  or (_23923_, _23922_, _23772_);
  nand (_23925_, _23923_, _03884_);
  and (_23926_, _09033_, _03014_);
  nor (_23927_, _23926_, _07782_);
  and (_23928_, _23927_, _23925_);
  and (_23929_, _08904_, _07782_);
  or (_23930_, _23929_, _23928_);
  nand (_23931_, _23930_, _09401_);
  nor (_23932_, _09429_, \oc8051_golden_model_1.DPH [3]);
  nor (_23933_, _23932_, _09430_);
  and (_23934_, _23933_, _09400_);
  nor (_23936_, _23934_, _09439_);
  nand (_23937_, _23936_, _23931_);
  nor (_23938_, _09438_, _08904_);
  nor (_23939_, _23938_, _09000_);
  nand (_23940_, _23939_, _23937_);
  and (_23941_, _08904_, _08190_);
  and (_23942_, _23766_, _08880_);
  or (_23943_, _23942_, _23941_);
  and (_23944_, _23943_, _09000_);
  nor (_23945_, _23944_, _20808_);
  and (_23947_, _23945_, _23940_);
  or (_23948_, _23947_, _23771_);
  nand (_23949_, _23948_, _09450_);
  nor (_23950_, _08904_, _09450_);
  nor (_23951_, _23950_, _03021_);
  nand (_23952_, _23951_, _23949_);
  not (_23953_, _09459_);
  and (_23954_, _09032_, _03021_);
  nor (_23955_, _23954_, _23953_);
  nand (_23956_, _23955_, _23952_);
  nor (_23958_, _09459_, _08904_);
  nor (_23959_, _23958_, _08994_);
  and (_23960_, _23959_, _23956_);
  or (_23961_, _23960_, _23769_);
  nand (_23962_, _23961_, _09473_);
  nor (_23963_, _23776_, _09473_);
  nor (_23964_, _23963_, _09476_);
  nand (_23965_, _23964_, _23962_);
  nor (_23966_, _08904_, _09475_);
  nor (_23967_, _23966_, _03020_);
  nand (_23969_, _23967_, _23965_);
  and (_23970_, _09032_, _03020_);
  nor (_23971_, _23970_, _10251_);
  and (_23972_, _23971_, _23969_);
  nor (_23973_, _08904_, _08877_);
  or (_23974_, _23973_, _08875_);
  or (_23975_, _23974_, _23972_);
  and (_23976_, _08904_, \oc8051_golden_model_1.PSW [7]);
  and (_23977_, _23766_, _07319_);
  or (_23978_, _23977_, _23976_);
  and (_23980_, _23978_, _08875_);
  nor (_23981_, _23980_, _09487_);
  and (_23982_, _23981_, _23975_);
  or (_23983_, _23982_, _23761_);
  nand (_23984_, _23983_, _07866_);
  nor (_23985_, _08904_, _07866_);
  nor (_23986_, _23985_, _03036_);
  nand (_23987_, _23986_, _23984_);
  not (_23988_, _08866_);
  and (_23989_, _09032_, _03036_);
  nor (_23991_, _23989_, _23988_);
  and (_23992_, _23991_, _23987_);
  or (_23993_, _23992_, _23760_);
  nor (_23994_, _23766_, _07319_);
  nor (_23995_, _08904_, \oc8051_golden_model_1.PSW [7]);
  nor (_23996_, _23995_, _08865_);
  not (_23997_, _23996_);
  nor (_23998_, _23997_, _23994_);
  nor (_23999_, _23998_, _09503_);
  and (_24000_, _23999_, _23993_);
  or (_24002_, _24000_, _23757_);
  nand (_24003_, _24002_, _08860_);
  nor (_24004_, _08904_, _08860_);
  nor (_24005_, _24004_, _08029_);
  nand (_24006_, _24005_, _24003_);
  and (_24007_, _23755_, _08029_);
  nor (_24008_, _24007_, _03148_);
  and (_24009_, _24008_, _24006_);
  and (_24010_, _04242_, _03148_);
  or (_24011_, _24010_, _24009_);
  nand (_24013_, _24011_, _05792_);
  and (_24014_, _23823_, _02531_);
  nor (_24015_, _24014_, _03035_);
  nand (_24016_, _24015_, _24013_);
  nor (_24017_, _09709_, _09032_);
  and (_24018_, _23783_, _09709_);
  or (_24019_, _24018_, _03152_);
  or (_24020_, _24019_, _24017_);
  and (_24021_, _24020_, _08858_);
  and (_24022_, _24021_, _24016_);
  or (_24024_, _24022_, _23756_);
  nand (_24025_, _24024_, _08104_);
  nor (_24026_, _08904_, _08104_);
  nor (_24027_, _24026_, _08135_);
  and (_24028_, _24027_, _24025_);
  and (_24029_, _23755_, _08135_);
  or (_24030_, _24029_, _02897_);
  nor (_24031_, _24030_, _24028_);
  and (_24032_, _04242_, _02897_);
  or (_24033_, _24032_, _24031_);
  nand (_24035_, _24033_, _09728_);
  and (_24036_, _23823_, _02536_);
  nor (_24037_, _24036_, _02895_);
  nand (_24038_, _24037_, _24035_);
  nor (_24039_, _23788_, _09709_);
  and (_24040_, _09709_, _09033_);
  nor (_24041_, _24040_, _24039_);
  and (_24042_, _24041_, _02895_);
  nor (_24043_, _24042_, _09737_);
  nand (_24044_, _24043_, _24038_);
  nor (_24046_, _23755_, _09736_);
  nor (_24047_, _24046_, _03166_);
  nand (_24048_, _24047_, _24044_);
  and (_24049_, _08904_, _03166_);
  nor (_24050_, _24049_, _09744_);
  nand (_24051_, _24050_, _24048_);
  nor (_24052_, _23755_, _09743_);
  nor (_24053_, _24052_, _03004_);
  and (_24054_, _24053_, _24051_);
  nor (_24055_, _06195_, _02799_);
  or (_24057_, _24055_, _02528_);
  or (_24058_, _24057_, _24054_);
  and (_24059_, _23823_, _02528_);
  nor (_24060_, _24059_, _02500_);
  nand (_24061_, _24060_, _24058_);
  and (_24062_, _24041_, _02500_);
  nor (_24063_, _24062_, _09759_);
  nand (_24064_, _24063_, _24061_);
  nor (_24065_, _23755_, _09758_);
  nor (_24066_, _24065_, _03174_);
  nand (_24068_, _24066_, _24064_);
  and (_24069_, _08904_, _03174_);
  nor (_24070_, _24069_, _09766_);
  nand (_24071_, _24070_, _24068_);
  nor (_24072_, _23755_, _09765_);
  nor (_24073_, _24072_, _03006_);
  nand (_24074_, _24073_, _24071_);
  nor (_24075_, _09770_, _02799_);
  nor (_24076_, _24075_, _02526_);
  and (_24077_, _24076_, _24074_);
  and (_24079_, _23823_, _02526_);
  nor (_24080_, _24079_, _24077_);
  and (_24081_, _24080_, _09778_);
  and (_24082_, _23755_, _09777_);
  or (_24083_, _24082_, _24081_);
  or (_24084_, _24083_, _34702_);
  or (_24085_, _34698_, \oc8051_golden_model_1.PC [11]);
  and (_24086_, _24085_, _36029_);
  and (_35251_, _24086_, _24084_);
  nor (_24087_, _08844_, \oc8051_golden_model_1.PC [12]);
  nor (_24089_, _24087_, _08845_);
  not (_24090_, _24089_);
  and (_24091_, _24090_, _08135_);
  nor (_24092_, _11423_, _08866_);
  nor (_24093_, _11423_, _08877_);
  nor (_24094_, _09459_, _11423_);
  nor (_24095_, _09438_, _11423_);
  and (_24096_, _09124_, _09121_);
  nor (_24097_, _24096_, _09125_);
  nor (_24098_, _24097_, _09169_);
  nor (_24100_, _09170_, _09027_);
  or (_24101_, _24100_, _09172_);
  nor (_24102_, _24101_, _24098_);
  and (_24103_, _11423_, _02950_);
  nor (_24104_, _24089_, _09234_);
  and (_24105_, _24089_, _07452_);
  or (_24106_, _24090_, _09207_);
  nand (_24107_, _09203_, _09204_);
  not (_24108_, \oc8051_golden_model_1.PC [12]);
  nor (_24109_, _03825_, _24108_);
  nand (_24111_, _24109_, _09206_);
  or (_24112_, _24111_, _24107_);
  and (_24113_, _24112_, _24106_);
  or (_24114_, _24113_, _03824_);
  or (_24115_, _24090_, _09203_);
  or (_24116_, _09213_, _11423_);
  and (_24117_, _24116_, _07433_);
  and (_24118_, _24117_, _24115_);
  and (_24119_, _24118_, _24114_);
  nand (_24120_, _11423_, _02954_);
  and (_24122_, _24120_, _09202_);
  not (_24123_, _24122_);
  nor (_24124_, _24123_, _24119_);
  nor (_24125_, _24124_, _24105_);
  nor (_24126_, _24125_, _09224_);
  nor (_24127_, _11423_, _02563_);
  nor (_24128_, _24127_, _10433_);
  not (_24129_, _24128_);
  nor (_24130_, _24129_, _24126_);
  and (_24131_, _09196_, _08899_);
  nor (_24133_, _08979_, _08977_);
  nor (_24134_, _24133_, _08980_);
  and (_24135_, _24134_, _09198_);
  or (_24136_, _24135_, _05387_);
  nor (_24137_, _24136_, _24131_);
  nor (_24138_, _24137_, _24130_);
  nor (_24139_, _24138_, _23804_);
  and (_24140_, _24097_, _09186_);
  not (_24141_, _24140_);
  and (_24142_, _09188_, _09027_);
  nor (_24144_, _24142_, _03821_);
  and (_24145_, _24144_, _24141_);
  nor (_24146_, _24145_, _24139_);
  nor (_24147_, _24146_, _21709_);
  nor (_24148_, _24147_, _24104_);
  nor (_24149_, _24148_, _09233_);
  nor (_24150_, _09177_, _08899_);
  nor (_24151_, _24150_, _09240_);
  not (_24152_, _24151_);
  nor (_24153_, _24152_, _24149_);
  nor (_24155_, _24090_, _09239_);
  nor (_24156_, _24155_, _02950_);
  not (_24157_, _24156_);
  nor (_24158_, _24157_, _24153_);
  nor (_24159_, _24158_, _24103_);
  nor (_24160_, _24159_, _09249_);
  nor (_24161_, _24089_, _09247_);
  nor (_24162_, _24161_, _09254_);
  not (_24163_, _24162_);
  nor (_24164_, _24163_, _24160_);
  nor (_24166_, _09253_, _11423_);
  nor (_24167_, _24166_, _09299_);
  not (_24168_, _24167_);
  or (_24169_, _24168_, _24164_);
  and (_24170_, _09297_, _09027_);
  not (_24171_, _24097_);
  nor (_24172_, _24171_, _09297_);
  or (_24173_, _24172_, _24170_);
  nor (_24174_, _24173_, _09263_);
  nor (_24175_, _24174_, _03038_);
  and (_24177_, _24175_, _24169_);
  or (_24178_, _24177_, _02966_);
  or (_24179_, _24178_, _24102_);
  nor (_24180_, _24171_, _09334_);
  and (_24181_, _09334_, _09027_);
  or (_24182_, _24181_, _03377_);
  or (_24183_, _24182_, _24180_);
  and (_24184_, _24183_, _10029_);
  nand (_24185_, _24184_, _24179_);
  and (_24186_, _09325_, _09027_);
  and (_24188_, _24097_, _21083_);
  or (_24189_, _24188_, _24186_);
  and (_24190_, _24189_, _03025_);
  nor (_24191_, _24190_, _09305_);
  and (_24192_, _24191_, _24185_);
  and (_24193_, _24090_, _09305_);
  or (_24194_, _24193_, _24192_);
  and (_24195_, _24194_, _09314_);
  nor (_24196_, _09314_, _08899_);
  or (_24197_, _24196_, _24195_);
  nand (_24199_, _24197_, _09012_);
  nor (_24200_, _24089_, _09012_);
  nor (_24201_, _24200_, _23775_);
  nand (_24202_, _24201_, _24199_);
  nor (_24203_, _09349_, _11423_);
  nor (_24204_, _24203_, _13666_);
  nand (_24205_, _24204_, _24202_);
  nor (_24206_, _24089_, _09005_);
  nor (_24207_, _24206_, _07597_);
  nand (_24208_, _24207_, _24205_);
  nor (_24210_, _11423_, _07596_);
  nor (_24211_, _24210_, _02585_);
  nand (_24212_, _24211_, _24208_);
  and (_24213_, _24090_, _02585_);
  nor (_24214_, _24213_, _09362_);
  nand (_24215_, _24214_, _24212_);
  nor (_24216_, _09361_, _11423_);
  nor (_24217_, _24216_, _03023_);
  nand (_24218_, _24217_, _24215_);
  nor (_24219_, _09027_, _08235_);
  nor (_24221_, _24219_, _20391_);
  nand (_24222_, _24221_, _24218_);
  nor (_24223_, _09369_, _11423_);
  nor (_24224_, _24223_, _02576_);
  nand (_24225_, _24224_, _24222_);
  nor (_24226_, _09027_, _02851_);
  nor (_24227_, _24226_, _09378_);
  nand (_24228_, _24227_, _24225_);
  nor (_24229_, _24090_, _09376_);
  nor (_24230_, _24229_, _09381_);
  nand (_24232_, _24230_, _24228_);
  nor (_24233_, _09380_, _08899_);
  nor (_24234_, _24233_, _09384_);
  and (_24235_, _24234_, _24232_);
  and (_24236_, _24134_, _09384_);
  nor (_24237_, _24236_, _24235_);
  or (_24238_, _24237_, _05562_);
  or (_24239_, _11423_, _05322_);
  and (_24240_, _24239_, _03884_);
  nand (_24241_, _24240_, _24238_);
  nor (_24243_, _09027_, _03884_);
  nor (_24244_, _24243_, _07782_);
  nand (_24245_, _24244_, _24241_);
  and (_24246_, _08899_, _07782_);
  nor (_24247_, _24246_, _09400_);
  nand (_24248_, _24247_, _24245_);
  nor (_24249_, _09430_, \oc8051_golden_model_1.DPH [4]);
  nor (_24250_, _24249_, _09431_);
  nor (_24251_, _24250_, _09401_);
  nor (_24252_, _24251_, _09439_);
  and (_24254_, _24252_, _24248_);
  or (_24255_, _24254_, _24095_);
  nand (_24256_, _24255_, _09442_);
  and (_24257_, _08899_, _08190_);
  and (_24258_, _24134_, _08880_);
  or (_24259_, _24258_, _24257_);
  and (_24260_, _24259_, _09000_);
  nor (_24261_, _24260_, _20808_);
  nand (_24262_, _24261_, _24256_);
  nor (_24263_, _24089_, _09448_);
  nor (_24265_, _24263_, _09451_);
  nand (_24266_, _24265_, _24262_);
  nor (_24267_, _11423_, _09450_);
  nor (_24268_, _24267_, _03021_);
  nand (_24269_, _24268_, _24266_);
  nor (_24270_, _09027_, _05279_);
  nor (_24271_, _24270_, _23953_);
  and (_24272_, _24271_, _24269_);
  or (_24273_, _24272_, _24094_);
  nand (_24274_, _24273_, _09462_);
  nor (_24276_, _24134_, _08880_);
  nor (_24277_, _08899_, _08190_);
  nor (_24278_, _24277_, _09462_);
  not (_24279_, _24278_);
  nor (_24280_, _24279_, _24276_);
  nor (_24281_, _24280_, _20466_);
  nand (_24282_, _24281_, _24274_);
  nor (_24283_, _24089_, _09473_);
  nor (_24284_, _24283_, _09476_);
  nand (_24285_, _24284_, _24282_);
  nor (_24287_, _11423_, _09475_);
  nor (_24288_, _24287_, _03020_);
  nand (_24289_, _24288_, _24285_);
  nor (_24290_, _09027_, _05274_);
  nor (_24291_, _24290_, _10251_);
  and (_24292_, _24291_, _24289_);
  or (_24293_, _24292_, _24093_);
  nand (_24294_, _24293_, _08876_);
  or (_24295_, _24134_, \oc8051_golden_model_1.PSW [7]);
  or (_24296_, _08899_, _07319_);
  and (_24298_, _24296_, _08875_);
  and (_24299_, _24298_, _24295_);
  nor (_24300_, _24299_, _09487_);
  nand (_24301_, _24300_, _24294_);
  nor (_24302_, _24089_, _08873_);
  nor (_24303_, _24302_, _07867_);
  nand (_24304_, _24303_, _24301_);
  nor (_24305_, _11423_, _07866_);
  nor (_24306_, _24305_, _03036_);
  nand (_24307_, _24306_, _24304_);
  nor (_24309_, _09027_, _05781_);
  nor (_24310_, _24309_, _23988_);
  and (_24311_, _24310_, _24307_);
  or (_24312_, _24311_, _24092_);
  nand (_24313_, _24312_, _08865_);
  nor (_24314_, _24134_, _07319_);
  nor (_24315_, _08899_, \oc8051_golden_model_1.PSW [7]);
  nor (_24316_, _24315_, _08865_);
  not (_24317_, _24316_);
  nor (_24318_, _24317_, _24314_);
  nor (_24321_, _24318_, _09503_);
  nand (_24322_, _24321_, _24313_);
  nor (_24323_, _24089_, _08862_);
  nor (_24324_, _24323_, _08861_);
  nand (_24325_, _24324_, _24322_);
  nor (_24326_, _11423_, _08860_);
  nor (_24327_, _24326_, _08029_);
  nand (_24328_, _24327_, _24325_);
  and (_24329_, _24090_, _08029_);
  nor (_24330_, _24329_, _03148_);
  and (_24333_, _24330_, _24328_);
  nor (_24334_, _05202_, _10250_);
  or (_24335_, _24334_, _02531_);
  or (_24336_, _24335_, _24333_);
  and (_24337_, _11423_, _02531_);
  nor (_24338_, _24337_, _03035_);
  nand (_24339_, _24338_, _24336_);
  and (_24340_, _24171_, _09709_);
  nor (_24341_, _09709_, _09027_);
  or (_24342_, _24341_, _03152_);
  or (_24345_, _24342_, _24340_);
  and (_24346_, _24345_, _08858_);
  nand (_24347_, _24346_, _24339_);
  nor (_24348_, _24089_, _08858_);
  nor (_24349_, _24348_, _08105_);
  nand (_24350_, _24349_, _24347_);
  nor (_24351_, _11423_, _08104_);
  nor (_24352_, _24351_, _08135_);
  and (_24353_, _24352_, _24350_);
  or (_24354_, _24353_, _24091_);
  nand (_24357_, _24354_, _02898_);
  and (_24358_, _05202_, _02897_);
  nor (_24359_, _24358_, _02536_);
  and (_24360_, _24359_, _24357_);
  and (_24361_, _08899_, _02536_);
  or (_24362_, _24361_, _02895_);
  nor (_24363_, _24362_, _24360_);
  and (_24364_, _09709_, _09027_);
  nor (_24365_, _24171_, _09709_);
  or (_24366_, _24365_, _24364_);
  nor (_24369_, _24366_, _02896_);
  or (_24370_, _24369_, _24363_);
  and (_24371_, _24370_, _09736_);
  nor (_24372_, _24089_, _09736_);
  or (_24373_, _24372_, _24371_);
  nand (_24374_, _24373_, _03563_);
  and (_24375_, _11423_, _03166_);
  nor (_24376_, _24375_, _09744_);
  nand (_24377_, _24376_, _24374_);
  nor (_24378_, _24090_, _09743_);
  nor (_24381_, _24378_, _03004_);
  nand (_24382_, _24381_, _24377_);
  and (_24383_, _03625_, _03004_);
  nor (_24384_, _24383_, _02528_);
  and (_24385_, _24384_, _24382_);
  and (_24386_, _08899_, _02528_);
  or (_24387_, _24386_, _02500_);
  or (_24388_, _24387_, _24385_);
  nor (_24389_, _24366_, _02501_);
  nor (_24390_, _24389_, _09759_);
  nand (_24393_, _24390_, _24388_);
  nor (_24394_, _24090_, _09758_);
  nor (_24395_, _24394_, _03174_);
  nand (_24396_, _24395_, _24393_);
  and (_24397_, _11423_, _03174_);
  nor (_24398_, _24397_, _09766_);
  nand (_24399_, _24398_, _24396_);
  nor (_24400_, _24090_, _09765_);
  nor (_24401_, _24400_, _03006_);
  nand (_24402_, _24401_, _24399_);
  and (_24404_, _03625_, _03006_);
  nor (_24405_, _24404_, _02526_);
  nand (_24406_, _24405_, _24402_);
  and (_24407_, _08899_, _02526_);
  nor (_24408_, _24407_, _09777_);
  and (_24409_, _24408_, _24406_);
  and (_24410_, _24090_, _09777_);
  nor (_24411_, _24410_, _24409_);
  or (_24412_, _24411_, _34702_);
  or (_24413_, _34698_, \oc8051_golden_model_1.PC [12]);
  and (_24415_, _24413_, _36029_);
  and (_35252_, _24415_, _24412_);
  and (_24416_, _08842_, _08889_);
  and (_24417_, _24416_, \oc8051_golden_model_1.PC [12]);
  nor (_24418_, _24417_, _08887_);
  and (_24419_, _24417_, _08887_);
  or (_24420_, _24419_, _24418_);
  nor (_24421_, _24420_, _08858_);
  nor (_24422_, _24420_, _08862_);
  nor (_24423_, _08894_, _08866_);
  or (_24425_, _24423_, _08864_);
  nor (_24426_, _24420_, _08873_);
  nor (_24427_, _08894_, _08877_);
  or (_24428_, _24427_, _08875_);
  and (_24429_, _08894_, _08190_);
  or (_24430_, _08895_, _08896_);
  not (_24431_, _24430_);
  nor (_24432_, _24431_, _08981_);
  and (_24433_, _24431_, _08981_);
  nor (_24434_, _24433_, _24432_);
  nor (_24436_, _24434_, _08190_);
  or (_24437_, _24436_, _24429_);
  and (_24438_, _24437_, _09000_);
  nor (_24439_, _08894_, _05322_);
  and (_24440_, _09022_, _02576_);
  nor (_24441_, _24420_, _09005_);
  not (_24442_, _24420_);
  nor (_24443_, _24442_, _09012_);
  and (_24444_, _09325_, _09022_);
  or (_24445_, _09025_, _09024_);
  not (_24447_, _24445_);
  nor (_24448_, _24447_, _09126_);
  and (_24449_, _24447_, _09126_);
  nor (_24450_, _24449_, _24448_);
  nor (_24451_, _24450_, _09325_);
  or (_24452_, _24451_, _24444_);
  and (_24453_, _24452_, _03025_);
  and (_24454_, _09169_, _09023_);
  not (_24455_, _24450_);
  nor (_24456_, _24455_, _09169_);
  nor (_24458_, _24456_, _24454_);
  nor (_24459_, _24458_, _09172_);
  and (_24460_, _08894_, _02950_);
  nor (_24461_, _09177_, _08894_);
  nor (_24462_, _09186_, _09022_);
  and (_24463_, _24450_, _09186_);
  or (_24464_, _24463_, _03821_);
  or (_24465_, _24464_, _24462_);
  and (_24466_, _09196_, _08894_);
  nor (_24467_, _24434_, _09196_);
  or (_24469_, _24467_, _05387_);
  nor (_24470_, _24469_, _24466_);
  or (_24471_, _24420_, _09208_);
  and (_24472_, _09213_, _08887_);
  and (_24473_, _24472_, _09207_);
  nand (_24474_, _24473_, _09203_);
  and (_24475_, _24474_, _24471_);
  or (_24476_, _24475_, _02954_);
  not (_24477_, _08894_);
  nand (_24478_, _09213_, _07433_);
  nand (_24480_, _24478_, _24477_);
  and (_24481_, _24480_, _24476_);
  and (_24482_, _24481_, _09202_);
  and (_24483_, _24420_, _07452_);
  or (_24484_, _24483_, _24482_);
  and (_24485_, _24484_, _02563_);
  nor (_24486_, _24477_, _02563_);
  nor (_24487_, _24486_, _10433_);
  not (_24488_, _24487_);
  nor (_24489_, _24488_, _24485_);
  or (_24491_, _24489_, _23804_);
  or (_24492_, _24491_, _24470_);
  and (_24493_, _24492_, _24465_);
  or (_24494_, _24493_, _21709_);
  or (_24495_, _24442_, _09234_);
  and (_24496_, _24495_, _09177_);
  and (_24497_, _24496_, _24494_);
  nor (_24498_, _24497_, _24461_);
  nor (_24499_, _24498_, _09240_);
  nor (_24500_, _24420_, _09239_);
  nor (_24502_, _24500_, _02950_);
  not (_24503_, _24502_);
  nor (_24504_, _24503_, _24499_);
  nor (_24505_, _24504_, _24460_);
  nor (_24506_, _24505_, _09249_);
  nor (_24507_, _24442_, _09247_);
  nor (_24508_, _24507_, _09254_);
  not (_24509_, _24508_);
  nor (_24510_, _24509_, _24506_);
  nor (_24511_, _09253_, _08894_);
  or (_24513_, _24511_, _09299_);
  or (_24514_, _24513_, _24510_);
  and (_24515_, _09297_, _09023_);
  nor (_24516_, _24455_, _09297_);
  or (_24517_, _24516_, _09263_);
  or (_24518_, _24517_, _24515_);
  and (_24519_, _24518_, _09172_);
  and (_24520_, _24519_, _24514_);
  nor (_24521_, _24520_, _24459_);
  and (_24522_, _24521_, _03377_);
  nor (_24524_, _24450_, _09334_);
  and (_24525_, _09334_, _09022_);
  or (_24526_, _24525_, _24524_);
  and (_24527_, _24526_, _02966_);
  or (_24528_, _24527_, _24522_);
  and (_24529_, _24528_, _10029_);
  nor (_24530_, _24529_, _24453_);
  nor (_24531_, _24530_, _09305_);
  and (_24532_, _24420_, _09305_);
  not (_24533_, _24532_);
  and (_24535_, _24533_, _09314_);
  not (_24536_, _24535_);
  nor (_24537_, _24536_, _24531_);
  nor (_24538_, _09314_, _08894_);
  nor (_24539_, _24538_, _20047_);
  not (_24540_, _24539_);
  nor (_24541_, _24540_, _24537_);
  nor (_24542_, _24541_, _24443_);
  nor (_24543_, _24542_, _23775_);
  nor (_24544_, _09349_, _24477_);
  nor (_24546_, _24544_, _13666_);
  not (_24547_, _24546_);
  nor (_24548_, _24547_, _24543_);
  nor (_24549_, _24548_, _24441_);
  nor (_24550_, _24549_, _07597_);
  nor (_24551_, _08894_, _07596_);
  nor (_24552_, _24551_, _02585_);
  not (_24553_, _24552_);
  nor (_24554_, _24553_, _24550_);
  and (_24555_, _24420_, _02585_);
  nor (_24557_, _24555_, _09362_);
  not (_24558_, _24557_);
  nor (_24559_, _24558_, _24554_);
  nor (_24560_, _09361_, _08894_);
  nor (_24561_, _24560_, _03023_);
  not (_24562_, _24561_);
  or (_24563_, _24562_, _24559_);
  and (_24564_, _09022_, _03023_);
  nor (_24565_, _24564_, _20391_);
  and (_24566_, _24565_, _24563_);
  nor (_24568_, _09369_, _08894_);
  nor (_24569_, _24568_, _02576_);
  not (_24570_, _24569_);
  nor (_24571_, _24570_, _24566_);
  or (_24572_, _24571_, _24440_);
  nand (_24573_, _24572_, _09376_);
  nor (_24574_, _24442_, _09376_);
  nor (_24575_, _24574_, _09381_);
  nand (_24576_, _24575_, _24573_);
  nor (_24577_, _09380_, _08894_);
  nor (_24579_, _24577_, _09384_);
  nand (_24580_, _24579_, _24576_);
  nor (_24581_, _24434_, _09385_);
  nor (_24582_, _24581_, _05562_);
  and (_24583_, _24582_, _24580_);
  or (_24584_, _24583_, _24439_);
  nand (_24585_, _24584_, _03884_);
  and (_24586_, _09023_, _03014_);
  nor (_24587_, _24586_, _07782_);
  and (_24588_, _24587_, _24585_);
  and (_24590_, _08894_, _07782_);
  or (_24591_, _24590_, _24588_);
  nand (_24592_, _24591_, _09401_);
  nor (_24593_, _09431_, \oc8051_golden_model_1.DPH [5]);
  nor (_24594_, _24593_, _09432_);
  and (_24595_, _24594_, _09400_);
  nor (_24596_, _24595_, _09439_);
  nand (_24597_, _24596_, _24592_);
  nor (_24598_, _09438_, _08894_);
  nor (_24599_, _24598_, _09000_);
  and (_24601_, _24599_, _24597_);
  or (_24602_, _24601_, _24438_);
  nand (_24603_, _24602_, _09448_);
  nor (_24604_, _24442_, _09448_);
  nor (_24605_, _24604_, _09451_);
  nand (_24606_, _24605_, _24603_);
  nor (_24607_, _08894_, _09450_);
  nor (_24608_, _24607_, _03021_);
  nand (_24609_, _24608_, _24606_);
  and (_24610_, _09022_, _03021_);
  nor (_24612_, _24610_, _23953_);
  nand (_24613_, _24612_, _24609_);
  nor (_24614_, _09459_, _08894_);
  nor (_24615_, _24614_, _08994_);
  nand (_24616_, _24615_, _24613_);
  nand (_24617_, _08894_, _08880_);
  or (_24618_, _24434_, _08880_);
  and (_24619_, _24618_, _24617_);
  or (_24620_, _24619_, _09462_);
  nand (_24621_, _24620_, _24616_);
  nand (_24623_, _24621_, _09473_);
  nor (_24624_, _24442_, _09473_);
  nor (_24625_, _24624_, _09476_);
  nand (_24626_, _24625_, _24623_);
  nor (_24627_, _08894_, _09475_);
  nor (_24628_, _24627_, _03020_);
  nand (_24629_, _24628_, _24626_);
  and (_24630_, _09022_, _03020_);
  nor (_24631_, _24630_, _10251_);
  and (_24632_, _24631_, _24629_);
  or (_24634_, _24632_, _24428_);
  and (_24635_, _24434_, _07319_);
  nor (_24636_, _08894_, _07319_);
  nor (_24637_, _24636_, _08876_);
  not (_24638_, _24637_);
  nor (_24639_, _24638_, _24635_);
  nor (_24640_, _24639_, _09487_);
  and (_24641_, _24640_, _24634_);
  or (_24642_, _24641_, _24426_);
  nand (_24643_, _24642_, _07866_);
  nor (_24645_, _08894_, _07866_);
  nor (_24646_, _24645_, _03036_);
  nand (_24647_, _24646_, _24643_);
  and (_24648_, _09022_, _03036_);
  nor (_24649_, _24648_, _23988_);
  and (_24650_, _24649_, _24647_);
  or (_24651_, _24650_, _24425_);
  and (_24652_, _24434_, \oc8051_golden_model_1.PSW [7]);
  nor (_24653_, _08894_, \oc8051_golden_model_1.PSW [7]);
  nor (_24654_, _24653_, _08865_);
  not (_24656_, _24654_);
  nor (_24657_, _24656_, _24652_);
  nor (_24658_, _24657_, _09503_);
  and (_24659_, _24658_, _24651_);
  or (_24660_, _24659_, _24422_);
  nand (_24661_, _24660_, _08860_);
  nor (_24662_, _08894_, _08860_);
  nor (_24663_, _24662_, _08029_);
  and (_24664_, _24663_, _24661_);
  and (_24665_, _24420_, _08029_);
  or (_24667_, _24665_, _03148_);
  nor (_24668_, _24667_, _24664_);
  and (_24669_, _04896_, _03148_);
  or (_24670_, _24669_, _24668_);
  nand (_24671_, _24670_, _05792_);
  and (_24672_, _24477_, _02531_);
  nor (_24673_, _24672_, _03035_);
  nand (_24674_, _24673_, _24671_);
  nor (_24675_, _09709_, _09022_);
  and (_24676_, _24450_, _09709_);
  or (_24678_, _24676_, _03152_);
  or (_24679_, _24678_, _24675_);
  and (_24680_, _24679_, _08858_);
  and (_24681_, _24680_, _24674_);
  or (_24682_, _24681_, _24421_);
  nand (_24683_, _24682_, _08104_);
  nor (_24684_, _08894_, _08104_);
  nor (_24685_, _24684_, _08135_);
  and (_24686_, _24685_, _24683_);
  and (_24687_, _24420_, _08135_);
  or (_24689_, _24687_, _02897_);
  nor (_24690_, _24689_, _24686_);
  and (_24691_, _04896_, _02897_);
  or (_24692_, _24691_, _24690_);
  nand (_24693_, _24692_, _09728_);
  and (_24694_, _24477_, _02536_);
  nor (_24695_, _24694_, _02895_);
  nand (_24696_, _24695_, _24693_);
  nor (_24697_, _24455_, _09709_);
  and (_24698_, _09709_, _09023_);
  nor (_24700_, _24698_, _24697_);
  and (_24701_, _24700_, _02895_);
  nor (_24702_, _24701_, _09737_);
  nand (_24703_, _24702_, _24696_);
  nor (_24704_, _24420_, _09736_);
  nor (_24705_, _24704_, _03166_);
  nand (_24706_, _24705_, _24703_);
  and (_24707_, _08894_, _03166_);
  nor (_24708_, _24707_, _09744_);
  nand (_24709_, _24708_, _24706_);
  nor (_24711_, _24420_, _09743_);
  nor (_24712_, _24711_, _03004_);
  nand (_24713_, _24712_, _24709_);
  nor (_24714_, _03215_, _06195_);
  nor (_24715_, _24714_, _02528_);
  nand (_24716_, _24715_, _24713_);
  and (_24717_, _24477_, _02528_);
  nor (_24718_, _24717_, _02500_);
  nand (_24719_, _24718_, _24716_);
  and (_24720_, _24700_, _02500_);
  nor (_24722_, _24720_, _09759_);
  nand (_24723_, _24722_, _24719_);
  nor (_24724_, _24420_, _09758_);
  nor (_24725_, _24724_, _03174_);
  nand (_24726_, _24725_, _24723_);
  and (_24727_, _08894_, _03174_);
  nor (_24728_, _24727_, _09766_);
  nand (_24729_, _24728_, _24726_);
  nor (_24730_, _24420_, _09765_);
  nor (_24731_, _24730_, _03006_);
  nand (_24733_, _24731_, _24729_);
  nor (_24734_, _03215_, _09770_);
  nor (_24735_, _24734_, _02526_);
  and (_24736_, _24735_, _24733_);
  and (_24737_, _24477_, _02526_);
  nor (_24738_, _24737_, _24736_);
  and (_24739_, _24738_, _09778_);
  and (_24740_, _24420_, _09777_);
  or (_24741_, _24740_, _24739_);
  or (_24742_, _24741_, _34702_);
  or (_24744_, _34698_, \oc8051_golden_model_1.PC [13]);
  and (_24745_, _24744_, _36029_);
  and (_35253_, _24745_, _24742_);
  nor (_24746_, _08846_, \oc8051_golden_model_1.PC [14]);
  nor (_24747_, _24746_, _08847_);
  not (_24748_, _24747_);
  and (_24749_, _24748_, _08135_);
  nor (_24750_, _11827_, _08866_);
  nor (_24751_, _11827_, _08877_);
  nor (_24752_, _09459_, _11827_);
  nor (_24755_, _09438_, _11827_);
  nor (_24756_, _09432_, \oc8051_golden_model_1.DPH [6]);
  nor (_24757_, _24756_, _09433_);
  nor (_24758_, _24757_, _09401_);
  and (_24759_, _08983_, _08886_);
  nor (_24760_, _24759_, _08985_);
  and (_24761_, _24760_, _09384_);
  or (_24762_, _24747_, _09012_);
  and (_24763_, _09169_, _09015_);
  and (_24764_, _09128_, _09020_);
  nor (_24766_, _24764_, _09129_);
  not (_24767_, _24766_);
  nor (_24768_, _24767_, _09169_);
  or (_24769_, _24768_, _24763_);
  or (_24770_, _24769_, _09172_);
  and (_24771_, _09297_, _09015_);
  nor (_24772_, _24767_, _09297_);
  or (_24773_, _24772_, _24771_);
  or (_24774_, _24773_, _09263_);
  or (_24775_, _24747_, _09234_);
  and (_24777_, _24747_, _09209_);
  and (_24778_, _24478_, _08882_);
  and (_24779_, _07433_, \oc8051_golden_model_1.PC [14]);
  and (_24780_, _24779_, _09213_);
  and (_24781_, _24780_, _09207_);
  and (_24782_, _24781_, _09203_);
  or (_24783_, _24782_, _24778_);
  and (_24784_, _24783_, _09202_);
  or (_24785_, _24784_, _24777_);
  and (_24786_, _24785_, _02563_);
  or (_24788_, _11827_, _02563_);
  nand (_24789_, _24788_, _05387_);
  or (_24790_, _24789_, _24786_);
  and (_24791_, _24760_, _09198_);
  and (_24792_, _09196_, _08882_);
  or (_24793_, _24792_, _05387_);
  or (_24794_, _24793_, _24791_);
  and (_24795_, _24794_, _24790_);
  or (_24796_, _24795_, _23804_);
  and (_24797_, _24766_, _09186_);
  and (_24799_, _09188_, _09015_);
  or (_24800_, _24799_, _03821_);
  or (_24801_, _24800_, _24797_);
  and (_24802_, _24801_, _24796_);
  or (_24803_, _24802_, _21709_);
  and (_24804_, _24803_, _24775_);
  or (_24805_, _24804_, _09233_);
  or (_24806_, _09177_, _08882_);
  and (_24807_, _24806_, _09239_);
  and (_24808_, _24807_, _24805_);
  nor (_24810_, _24748_, _09239_);
  or (_24811_, _24810_, _02950_);
  or (_24812_, _24811_, _24808_);
  nand (_24813_, _11827_, _02950_);
  and (_24814_, _24813_, _24812_);
  or (_24815_, _24814_, _09249_);
  or (_24816_, _24747_, _09247_);
  and (_24817_, _24816_, _09253_);
  and (_24818_, _24817_, _24815_);
  or (_24819_, _09253_, _11827_);
  nand (_24821_, _24819_, _09263_);
  or (_24822_, _24821_, _24818_);
  and (_24823_, _24822_, _24774_);
  or (_24824_, _24823_, _03038_);
  and (_24825_, _24824_, _24770_);
  or (_24826_, _24825_, _02966_);
  nor (_24827_, _24767_, _09334_);
  and (_24828_, _09334_, _09015_);
  or (_24829_, _24828_, _03377_);
  or (_24830_, _24829_, _24827_);
  and (_24832_, _24830_, _10029_);
  and (_24833_, _24832_, _24826_);
  or (_24834_, _24766_, _09325_);
  or (_24835_, _21083_, _09015_);
  and (_24836_, _24835_, _03025_);
  and (_24837_, _24836_, _24834_);
  or (_24838_, _24837_, _09305_);
  or (_24839_, _24838_, _24833_);
  nand (_24840_, _24748_, _09305_);
  and (_24841_, _24840_, _09314_);
  and (_24843_, _24841_, _24839_);
  nor (_24844_, _09314_, _11827_);
  or (_24845_, _24844_, _20047_);
  or (_24846_, _24845_, _24843_);
  and (_24847_, _24846_, _24762_);
  or (_24848_, _24847_, _23775_);
  or (_24849_, _09349_, _08882_);
  and (_24850_, _24849_, _09005_);
  and (_24851_, _24850_, _24848_);
  nor (_24852_, _24748_, _09005_);
  or (_24854_, _24852_, _07597_);
  nor (_24855_, _24854_, _24851_);
  nor (_24856_, _08882_, _07596_);
  nor (_24857_, _24856_, _24855_);
  nor (_24858_, _24857_, _02585_);
  and (_24859_, _24748_, _02585_);
  nor (_24860_, _24859_, _09362_);
  not (_24861_, _24860_);
  nor (_24862_, _24861_, _24858_);
  nor (_24863_, _09361_, _11827_);
  nor (_24865_, _24863_, _03023_);
  not (_24866_, _24865_);
  nor (_24867_, _24866_, _24862_);
  nor (_24868_, _09015_, _08235_);
  or (_24869_, _24868_, _20391_);
  or (_24870_, _24869_, _24867_);
  or (_24871_, _09369_, _11827_);
  and (_24872_, _24871_, _02851_);
  and (_24873_, _24872_, _24870_);
  nor (_24874_, _09015_, _02851_);
  nor (_24876_, _24874_, _09378_);
  not (_24877_, _24876_);
  nor (_24878_, _24877_, _24873_);
  nor (_24879_, _24748_, _09376_);
  or (_24880_, _24879_, _09381_);
  nor (_24881_, _24880_, _24878_);
  nor (_24882_, _09380_, _08882_);
  or (_24883_, _24882_, _09384_);
  nor (_24884_, _24883_, _24881_);
  nor (_24885_, _24884_, _24761_);
  and (_24887_, _24885_, _05322_);
  nor (_24888_, _08882_, _05322_);
  nor (_24889_, _24888_, _24887_);
  nand (_24890_, _24889_, _03884_);
  nand (_24891_, _09015_, _03014_);
  and (_24892_, _24891_, _24890_);
  or (_24893_, _24892_, _07782_);
  and (_24894_, _08882_, _07782_);
  nor (_24895_, _24894_, _09400_);
  and (_24896_, _24895_, _24893_);
  or (_24898_, _24896_, _09439_);
  nor (_24899_, _24898_, _24758_);
  or (_24900_, _24899_, _24755_);
  nand (_24901_, _24900_, _09442_);
  and (_24902_, _08882_, _08190_);
  and (_24903_, _24760_, _08880_);
  or (_24904_, _24903_, _24902_);
  and (_24905_, _24904_, _09000_);
  nor (_24906_, _24905_, _20808_);
  nand (_24907_, _24906_, _24901_);
  nor (_24909_, _24747_, _09448_);
  nor (_24910_, _24909_, _09451_);
  nand (_24911_, _24910_, _24907_);
  nor (_24912_, _11827_, _09450_);
  nor (_24913_, _24912_, _03021_);
  nand (_24914_, _24913_, _24911_);
  nor (_24915_, _09015_, _05279_);
  nor (_24916_, _24915_, _23953_);
  and (_24917_, _24916_, _24914_);
  or (_24918_, _24917_, _24752_);
  nand (_24920_, _24918_, _09462_);
  nor (_24921_, _24760_, _08880_);
  nor (_24922_, _08882_, _08190_);
  nor (_24923_, _24922_, _09462_);
  not (_24924_, _24923_);
  nor (_24925_, _24924_, _24921_);
  nor (_24926_, _24925_, _20466_);
  nand (_24927_, _24926_, _24920_);
  nor (_24928_, _24747_, _09473_);
  nor (_24929_, _24928_, _09476_);
  nand (_24931_, _24929_, _24927_);
  nor (_24932_, _11827_, _09475_);
  nor (_24933_, _24932_, _03020_);
  nand (_24934_, _24933_, _24931_);
  nor (_24935_, _09015_, _05274_);
  nor (_24936_, _24935_, _10251_);
  and (_24937_, _24936_, _24934_);
  or (_24938_, _24937_, _24751_);
  nand (_24939_, _24938_, _08876_);
  and (_24940_, _08882_, \oc8051_golden_model_1.PSW [7]);
  and (_24942_, _24760_, _07319_);
  or (_24943_, _24942_, _24940_);
  and (_24944_, _24943_, _08875_);
  nor (_24945_, _24944_, _09487_);
  nand (_24946_, _24945_, _24939_);
  nor (_24947_, _24747_, _08873_);
  nor (_24948_, _24947_, _07867_);
  nand (_24949_, _24948_, _24946_);
  nor (_24950_, _11827_, _07866_);
  nor (_24951_, _24950_, _03036_);
  nand (_24953_, _24951_, _24949_);
  nor (_24954_, _09015_, _05781_);
  nor (_24955_, _24954_, _23988_);
  and (_24956_, _24955_, _24953_);
  or (_24957_, _24956_, _24750_);
  nand (_24958_, _24957_, _08865_);
  nor (_24959_, _24760_, _07319_);
  nor (_24960_, _08882_, \oc8051_golden_model_1.PSW [7]);
  nor (_24961_, _24960_, _08865_);
  not (_24962_, _24961_);
  nor (_24964_, _24962_, _24959_);
  nor (_24965_, _24964_, _09503_);
  nand (_24966_, _24965_, _24958_);
  nor (_24967_, _24747_, _08862_);
  nor (_24968_, _24967_, _08861_);
  nand (_24969_, _24968_, _24966_);
  nor (_24970_, _11827_, _08860_);
  nor (_24971_, _24970_, _08029_);
  nand (_24972_, _24971_, _24969_);
  and (_24973_, _24748_, _08029_);
  nor (_24975_, _24973_, _03148_);
  and (_24976_, _24975_, _24972_);
  nor (_24977_, _04787_, _10250_);
  or (_24978_, _24977_, _02531_);
  or (_24979_, _24978_, _24976_);
  and (_24980_, _11827_, _02531_);
  nor (_24981_, _24980_, _03035_);
  nand (_24982_, _24981_, _24979_);
  and (_24983_, _24767_, _09709_);
  nor (_24984_, _09709_, _09015_);
  or (_24986_, _24984_, _03152_);
  or (_24987_, _24986_, _24983_);
  and (_24988_, _24987_, _08858_);
  nand (_24989_, _24988_, _24982_);
  nor (_24990_, _24747_, _08858_);
  nor (_24991_, _24990_, _08105_);
  nand (_24992_, _24991_, _24989_);
  nor (_24993_, _11827_, _08104_);
  nor (_24994_, _24993_, _08135_);
  and (_24995_, _24994_, _24992_);
  or (_24997_, _24995_, _24749_);
  nand (_24998_, _24997_, _02898_);
  and (_24999_, _04787_, _02897_);
  nor (_25000_, _24999_, _02536_);
  and (_25001_, _25000_, _24998_);
  and (_25002_, _08882_, _02536_);
  or (_25003_, _25002_, _02895_);
  nor (_25004_, _25003_, _25001_);
  and (_25005_, _09709_, _09015_);
  nor (_25006_, _24767_, _09709_);
  or (_25008_, _25006_, _25005_);
  nor (_25009_, _25008_, _02896_);
  or (_25010_, _25009_, _25004_);
  and (_25011_, _25010_, _09736_);
  nor (_25012_, _24747_, _09736_);
  or (_25013_, _25012_, _25011_);
  nand (_25014_, _25013_, _03563_);
  and (_25015_, _11827_, _03166_);
  nor (_25016_, _25015_, _09744_);
  nand (_25017_, _25016_, _25014_);
  nor (_25019_, _24748_, _09743_);
  nor (_25020_, _25019_, _03004_);
  nand (_25021_, _25020_, _25017_);
  and (_25022_, _03004_, _02932_);
  nor (_25023_, _25022_, _02528_);
  and (_25024_, _25023_, _25021_);
  and (_25025_, _08882_, _02528_);
  or (_25026_, _25025_, _02500_);
  or (_25027_, _25026_, _25024_);
  nor (_25028_, _25008_, _02501_);
  nor (_25030_, _25028_, _09759_);
  nand (_25031_, _25030_, _25027_);
  nor (_25032_, _24748_, _09758_);
  nor (_25033_, _25032_, _03174_);
  nand (_25034_, _25033_, _25031_);
  and (_25035_, _11827_, _03174_);
  nor (_25036_, _25035_, _09766_);
  nand (_25037_, _25036_, _25034_);
  nor (_25038_, _24748_, _09765_);
  nor (_25039_, _25038_, _03006_);
  nand (_25041_, _25039_, _25037_);
  and (_25042_, _03006_, _02932_);
  nor (_25043_, _25042_, _02526_);
  nand (_25044_, _25043_, _25041_);
  and (_25045_, _08882_, _02526_);
  nor (_25046_, _25045_, _09777_);
  and (_25047_, _25046_, _25044_);
  and (_25048_, _24748_, _09777_);
  nor (_25049_, _25048_, _25047_);
  or (_25050_, _25049_, _34702_);
  or (_25052_, _34698_, \oc8051_golden_model_1.PC [14]);
  and (_25053_, _25052_, _36029_);
  and (_35254_, _25053_, _25050_);
  not (_25054_, \oc8051_golden_model_1.PSW [0]);
  nor (_25055_, _34698_, _25054_);
  nor (_25056_, _06926_, _06925_);
  nor (_25057_, _25056_, _06833_);
  and (_25058_, _25056_, _06833_);
  nor (_25059_, _25058_, _25057_);
  nor (_25060_, _06850_, _06849_);
  nor (_25062_, _25060_, _13844_);
  and (_25063_, _25060_, _13844_);
  nor (_25064_, _25063_, _25062_);
  and (_25065_, _25064_, _25059_);
  nor (_25066_, _25064_, _25059_);
  nor (_25067_, _25066_, _25065_);
  nor (_25068_, _25067_, _05768_);
  and (_25069_, _25067_, _05768_);
  nor (_25070_, _25069_, _25068_);
  nor (_25071_, _08135_, _02897_);
  and (_25073_, _23401_, _25071_);
  or (_25074_, _25073_, _25070_);
  nor (_25075_, _03148_, _02531_);
  and (_25076_, _25075_, _03152_);
  or (_25077_, _25076_, _25070_);
  nor (_25078_, _13807_, _13344_);
  and (_25079_, _13807_, _13344_);
  or (_25080_, _25079_, _25078_);
  nor (_25081_, _25080_, _14115_);
  and (_25082_, _25080_, _14115_);
  nor (_25084_, _25082_, _25081_);
  and (_25085_, _25084_, _14416_);
  nor (_25086_, _25084_, _14416_);
  nor (_25087_, _25086_, _25085_);
  nor (_25088_, _25087_, _14712_);
  and (_25089_, _25087_, _14712_);
  or (_25090_, _25089_, _25088_);
  nor (_25091_, _25090_, _15035_);
  and (_25092_, _25090_, _15035_);
  or (_25093_, _25092_, _25091_);
  nor (_25095_, _25093_, _15104_);
  and (_25096_, _25093_, _15104_);
  or (_25097_, _25096_, _25095_);
  nor (_25098_, _25097_, _08025_);
  and (_25099_, _25097_, _08025_);
  or (_25100_, _25099_, _25098_);
  or (_25101_, _25100_, _03138_);
  and (_25102_, _08866_, _08865_);
  nor (_25103_, _13795_, _13514_);
  and (_25104_, _13795_, _13514_);
  or (_25106_, _25104_, _25103_);
  nor (_25107_, _14402_, _14100_);
  and (_25108_, _14402_, _14100_);
  nor (_25109_, _25108_, _25107_);
  nor (_25110_, _25109_, _25106_);
  and (_25111_, _25109_, _25106_);
  nor (_25112_, _25111_, _25110_);
  nor (_25113_, _15346_, _15022_);
  and (_25114_, _15346_, _15022_);
  nor (_25115_, _25114_, _25113_);
  not (_25117_, _14699_);
  and (_25118_, _25117_, _07876_);
  nor (_25119_, _25117_, _07876_);
  nor (_25120_, _25119_, _25118_);
  nor (_25121_, _25120_, _25115_);
  and (_25122_, _25120_, _25115_);
  nor (_25123_, _25122_, _25121_);
  not (_25124_, _25123_);
  nand (_25125_, _25124_, _25112_);
  or (_25126_, _25124_, _25112_);
  and (_25128_, _25126_, _03036_);
  and (_25129_, _25128_, _25125_);
  or (_25130_, _08157_, _08154_);
  nand (_25131_, _08157_, _08154_);
  and (_25132_, _25131_, _25130_);
  not (_25133_, _08148_);
  and (_25134_, _25133_, _08150_);
  nor (_25135_, _25133_, _08150_);
  nor (_25136_, _25135_, _25134_);
  and (_25137_, _25136_, _25132_);
  nor (_25139_, _25136_, _25132_);
  nor (_25140_, _25139_, _25137_);
  nor (_25141_, _08137_, _07819_);
  and (_25142_, _08137_, _07819_);
  nor (_25143_, _25142_, _25141_);
  nor (_25144_, _08140_, _08144_);
  and (_25145_, _08140_, _08144_);
  nor (_25146_, _25145_, _25144_);
  nor (_25147_, _25146_, _25143_);
  and (_25148_, _25146_, _25143_);
  or (_25150_, _25148_, _25147_);
  not (_25151_, _25150_);
  nor (_25152_, _25151_, _25140_);
  and (_25153_, _25151_, _25140_);
  or (_25154_, _25153_, _25152_);
  and (_25155_, _25154_, _07836_);
  nor (_25156_, _02942_, _04125_);
  not (_25157_, _13942_);
  and (_25158_, _25157_, _13655_);
  nor (_25159_, _25157_, _13655_);
  nor (_25161_, _25159_, _25158_);
  and (_25162_, _25161_, _14821_);
  nor (_25163_, _25161_, _14821_);
  or (_25164_, _25163_, _25162_);
  not (_25165_, _25164_);
  not (_25166_, _13374_);
  nor (_25167_, _14212_, _25166_);
  and (_25168_, _14212_, _25166_);
  nor (_25169_, _25168_, _25167_);
  not (_25170_, _25169_);
  not (_25172_, _14549_);
  and (_25173_, _25172_, _07510_);
  nor (_25174_, _25172_, _07510_);
  nor (_25175_, _25174_, _25173_);
  and (_25176_, _25175_, _15199_);
  nor (_25177_, _25175_, _15199_);
  nor (_25178_, _25177_, _25176_);
  nor (_25179_, _25178_, _25170_);
  and (_25180_, _25178_, _25170_);
  nor (_25181_, _25180_, _25179_);
  nand (_25183_, _25181_, _25165_);
  or (_25184_, _25181_, _25165_);
  and (_25185_, _25184_, _02880_);
  and (_25186_, _25185_, _25183_);
  or (_25187_, _06178_, _06030_);
  nand (_25188_, _25187_, _10802_);
  or (_25189_, _25187_, _10802_);
  nand (_25190_, _25189_, _25188_);
  nor (_25191_, _06182_, _06122_);
  nand (_25192_, _25191_, _05847_);
  or (_25194_, _25191_, _05847_);
  and (_25195_, _25194_, _25192_);
  nand (_25196_, _25195_, _25190_);
  or (_25197_, _25195_, _25190_);
  nand (_25198_, _25197_, _25196_);
  nor (_25199_, _25198_, _05490_);
  and (_25200_, _25198_, _05490_);
  or (_25201_, _25200_, _25199_);
  or (_25202_, _25201_, _02465_);
  and (_25203_, _25202_, _03413_);
  or (_25205_, _25201_, _07436_);
  nor (_25206_, _10608_, _06160_);
  and (_25207_, _10608_, _06160_);
  nor (_25208_, _25207_, _25206_);
  nor (_25209_, _06162_, _05262_);
  not (_25210_, _25209_);
  nor (_25211_, _09194_, _09791_);
  nor (_25212_, _25211_, _06159_);
  and (_25213_, _25211_, _06159_);
  nor (_25214_, _25213_, _25212_);
  and (_25216_, _25214_, _25210_);
  nor (_25217_, _25214_, _25210_);
  or (_25218_, _25217_, _25216_);
  nand (_25219_, _25218_, _25208_);
  or (_25220_, _25218_, _25208_);
  and (_25221_, _25220_, _25219_);
  or (_25222_, _25221_, _07440_);
  and (_25223_, _09213_, _09207_);
  and (_25224_, _25223_, _25054_);
  nor (_25225_, _25223_, _25070_);
  or (_25227_, _25225_, _25224_);
  nand (_25228_, _25227_, _09203_);
  and (_25229_, _25228_, _25222_);
  and (_25230_, _25229_, _25205_);
  or (_25231_, _25230_, _02954_);
  and (_25232_, _07640_, _07624_);
  nor (_25233_, _25232_, _07959_);
  nor (_25234_, _07651_, _07610_);
  and (_25235_, _07651_, _07610_);
  nor (_25236_, _25235_, _25234_);
  and (_25237_, _25236_, _25233_);
  nor (_25238_, _25236_, _25233_);
  nor (_25239_, _25238_, _25237_);
  nor (_25240_, _07681_, _05528_);
  and (_25241_, _07681_, _05528_);
  nor (_25242_, _25241_, _25240_);
  nor (_25243_, _07700_, _07670_);
  and (_25244_, _07700_, _07670_);
  nor (_25245_, _25244_, _25243_);
  nor (_25246_, _25245_, _25242_);
  and (_25249_, _25245_, _25242_);
  or (_25250_, _25249_, _25246_);
  and (_25251_, _25250_, _25239_);
  nor (_25252_, _25250_, _25239_);
  or (_25253_, _25252_, _25251_);
  or (_25254_, _25253_, _07433_);
  and (_25255_, _25254_, _09202_);
  nand (_25256_, _25255_, _25231_);
  nand (_25257_, _25256_, _22821_);
  or (_25258_, _25070_, _22821_);
  and (_25260_, _25258_, _05402_);
  and (_25261_, _25260_, _25257_);
  nor (_25262_, _25060_, \oc8051_golden_model_1.ACC [6]);
  and (_25263_, _25060_, \oc8051_golden_model_1.ACC [6]);
  nor (_25264_, _25263_, _25262_);
  nor (_25265_, _25264_, \oc8051_golden_model_1.ACC [7]);
  and (_25266_, _25264_, \oc8051_golden_model_1.ACC [7]);
  nor (_25267_, _25266_, _25265_);
  or (_25268_, _25267_, _25190_);
  nand (_25269_, _25267_, _25190_);
  and (_25271_, _25269_, _25268_);
  and (_25272_, _25271_, _03818_);
  or (_25273_, _25272_, _02952_);
  or (_25274_, _25273_, _25261_);
  not (_25275_, _15159_);
  nor (_25276_, _13616_, _25166_);
  and (_25277_, _13616_, _25166_);
  nor (_25278_, _25277_, _25276_);
  and (_25279_, _25278_, _13905_);
  nor (_25280_, _25278_, _13905_);
  nor (_25281_, _25280_, _25279_);
  and (_25282_, _25281_, _14840_);
  nor (_25283_, _25281_, _14840_);
  or (_25284_, _25283_, _25282_);
  nor (_25285_, _14514_, _14231_);
  and (_25286_, _14514_, _14231_);
  nor (_25287_, _25286_, _25285_);
  and (_25288_, _25287_, _25284_);
  nor (_25289_, _25287_, _25284_);
  nor (_25290_, _25289_, _25288_);
  nor (_25293_, _25290_, _25275_);
  and (_25294_, _25290_, _25275_);
  or (_25295_, _25294_, _25293_);
  and (_25296_, _25295_, _07457_);
  nor (_25297_, _25295_, _07457_);
  or (_25298_, _25297_, _25296_);
  nor (_25299_, _25298_, _03821_);
  nor (_25300_, _25299_, _07455_);
  and (_25301_, _25300_, _25274_);
  and (_25302_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_25304_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_25305_, _25304_, _25302_);
  and (_25306_, _25305_, _13622_);
  nor (_25307_, _25305_, _13622_);
  nor (_25308_, _25307_, _25306_);
  and (_25309_, _14520_, _14238_);
  and (_25310_, _14519_, _14239_);
  nor (_25311_, _25310_, _25309_);
  nor (_25312_, _25311_, _25308_);
  and (_25313_, _25311_, _25308_);
  nor (_25314_, _25313_, _25312_);
  and (_25315_, _25314_, _14847_);
  nor (_25316_, _25314_, _14847_);
  nor (_25317_, _25316_, _25315_);
  nor (_25318_, _15167_, _07480_);
  and (_25319_, _15167_, _07480_);
  nor (_25320_, _25319_, _25318_);
  not (_25321_, _25320_);
  nand (_25322_, _25321_, _25317_);
  or (_25323_, _25321_, _25317_);
  and (_25326_, _25323_, _25322_);
  and (_25327_, _25326_, _07455_);
  or (_25328_, _25327_, _09179_);
  or (_25329_, _25328_, _25301_);
  not (_25330_, _25070_);
  nand (_25331_, _25330_, _09179_);
  and (_25332_, _25331_, _02892_);
  and (_25333_, _25332_, _25329_);
  and (_25334_, _13630_, _13380_);
  nor (_25335_, _13630_, _13380_);
  or (_25337_, _25335_, _25334_);
  not (_25338_, _14243_);
  and (_25339_, _25338_, _13919_);
  nor (_25340_, _25338_, _13919_);
  nor (_25341_, _25340_, _25339_);
  and (_25342_, _25341_, _25337_);
  nor (_25343_, _25341_, _25337_);
  or (_25344_, _25343_, _25342_);
  nor (_25345_, _14851_, _14526_);
  and (_25346_, _14851_, _14526_);
  nor (_25348_, _25346_, _25345_);
  and (_25349_, _25348_, _15174_);
  nor (_25350_, _25348_, _15174_);
  nor (_25351_, _25350_, _25349_);
  nor (_25352_, _25351_, _25344_);
  and (_25353_, _25351_, _25344_);
  nor (_25354_, _25353_, _25352_);
  and (_25355_, _25354_, _07486_);
  nor (_25356_, _25354_, _07486_);
  or (_25357_, _25356_, _25355_);
  and (_25359_, _25357_, _02891_);
  or (_25360_, _25359_, _22787_);
  or (_25361_, _25360_, _25333_);
  and (_25362_, _13586_, _13352_);
  nor (_25363_, _13586_, _13352_);
  nor (_25364_, _25363_, _25362_);
  not (_25365_, _25364_);
  not (_25366_, _14194_);
  and (_25367_, _25366_, _13877_);
  nor (_25368_, _25366_, _13877_);
  nor (_25369_, _25368_, _25367_);
  and (_25370_, _25369_, _25365_);
  nor (_25371_, _25369_, _25365_);
  nor (_25372_, _25371_, _25370_);
  nor (_25373_, _14800_, _14493_);
  and (_25374_, _14800_, _14493_);
  nor (_25375_, _25374_, _25373_);
  and (_25376_, _25375_, _15122_);
  nor (_25377_, _25375_, _15122_);
  nor (_25378_, _25377_, _25376_);
  nor (_25381_, _25378_, _25372_);
  and (_25382_, _25378_, _25372_);
  nor (_25383_, _25382_, _25381_);
  nand (_25384_, _25383_, _07274_);
  or (_25385_, _25383_, _07274_);
  and (_25386_, _25385_, _25384_);
  or (_25387_, _25386_, _03327_);
  or (_25388_, _25070_, _02556_);
  and (_25389_, _25388_, _07430_);
  and (_25390_, _25389_, _25387_);
  and (_25392_, _25390_, _25361_);
  and (_25393_, _25221_, _07431_);
  or (_25394_, _25393_, _25392_);
  and (_25395_, _25394_, _03849_);
  or (_25396_, _25395_, _25203_);
  not (_25397_, _03414_);
  or (_25398_, _25201_, _25397_);
  and (_25399_, _25398_, _02959_);
  and (_25400_, _25399_, _25396_);
  and (_25401_, _25253_, _02950_);
  or (_25403_, _25401_, _09249_);
  or (_25404_, _25403_, _25400_);
  or (_25405_, _25070_, _09247_);
  and (_25406_, _25405_, _02888_);
  and (_25407_, _25406_, _25404_);
  nor (_25408_, _13650_, _13350_);
  and (_25409_, _13650_, _13350_);
  nor (_25410_, _25409_, _25408_);
  not (_25411_, _25410_);
  not (_25412_, _14262_);
  and (_25414_, _25412_, _13937_);
  nor (_25415_, _25412_, _13937_);
  nor (_25416_, _25415_, _25414_);
  and (_25417_, _25416_, _25411_);
  nor (_25418_, _25416_, _25411_);
  nor (_25419_, _25418_, _25417_);
  nor (_25420_, _14870_, _14544_);
  and (_25421_, _14870_, _14544_);
  nor (_25422_, _25421_, _25420_);
  not (_25423_, _15193_);
  and (_25425_, _25423_, _07505_);
  nor (_25426_, _25423_, _07505_);
  or (_25427_, _25426_, _25425_);
  or (_25428_, _25427_, _25422_);
  nand (_25429_, _25427_, _25422_);
  and (_25430_, _25429_, _25428_);
  nor (_25431_, _25430_, _25419_);
  and (_25432_, _25430_, _25419_);
  or (_25433_, _25432_, _25431_);
  nand (_25434_, _25433_, _02887_);
  and (_25436_, _09262_, _09172_);
  and (_25437_, _25436_, _09252_);
  and (_25438_, _09308_, _09258_);
  and (_25439_, _25438_, _25437_);
  nand (_25440_, _25439_, _25434_);
  or (_25441_, _25440_, _25407_);
  or (_25442_, _25439_, _25070_);
  and (_25443_, _25442_, _02881_);
  and (_25444_, _25443_, _25441_);
  or (_25445_, _25444_, _25186_);
  and (_25447_, _25445_, _25156_);
  or (_25448_, _25330_, _25156_);
  and (_25449_, _02982_, _10788_);
  nor (_25450_, _25449_, _02978_);
  nand (_25451_, _25450_, _25448_);
  or (_25452_, _25451_, _25447_);
  nor (_25453_, _25450_, _25070_);
  and (_25454_, _02981_, _02498_);
  nor (_25455_, _25454_, _25453_);
  and (_25456_, _25455_, _25452_);
  nor (_25458_, _09009_, _03867_);
  nand (_25459_, _25454_, _25070_);
  nand (_25460_, _25459_, _25458_);
  or (_25461_, _25460_, _25456_);
  or (_25462_, _25458_, _25070_);
  and (_25463_, _25462_, _06277_);
  and (_25464_, _25463_, _25461_);
  nor (_25465_, _02987_, _09347_);
  and (_25466_, _25465_, _08251_);
  nor (_25467_, _13661_, _06732_);
  nor (_25469_, _13662_, _13404_);
  nor (_25470_, _25469_, _25467_);
  nor (_25471_, _25470_, _13947_);
  and (_25472_, _25470_, _13947_);
  nor (_25473_, _25472_, _25471_);
  nor (_25474_, _25473_, _14269_);
  and (_25475_, _25473_, _14269_);
  or (_25476_, _25475_, _25474_);
  not (_25477_, _25476_);
  nor (_25478_, _25477_, _14554_);
  and (_25480_, _25477_, _14554_);
  nor (_25481_, _25480_, _25478_);
  nor (_25482_, _25481_, _14878_);
  and (_25483_, _25481_, _14878_);
  or (_25484_, _25483_, _25482_);
  not (_25485_, _25484_);
  nor (_25486_, _25485_, _15204_);
  and (_25487_, _25485_, _15204_);
  nor (_25488_, _25487_, _25486_);
  and (_25489_, _25488_, _07515_);
  nor (_25491_, _25488_, _07515_);
  or (_25492_, _25491_, _25489_);
  nand (_25493_, _25492_, _06271_);
  nand (_25494_, _25493_, _25466_);
  or (_25495_, _25494_, _25464_);
  or (_25496_, _25466_, _25070_);
  and (_25497_, _25496_, _09809_);
  and (_25498_, _25497_, _25495_);
  nand (_25499_, _25070_, _02986_);
  nand (_25500_, _25499_, _07426_);
  or (_25501_, _25500_, _25498_);
  not (_25502_, _14571_);
  not (_25503_, _07577_);
  and (_25504_, _13673_, _25503_);
  nor (_25505_, _25504_, _07578_);
  and (_25506_, _25505_, _13965_);
  nor (_25507_, _25505_, _13965_);
  or (_25508_, _25507_, _25506_);
  nor (_25509_, _25508_, _14283_);
  and (_25510_, _25508_, _14283_);
  nor (_25513_, _25510_, _25509_);
  and (_25514_, _25513_, _25502_);
  nor (_25515_, _25513_, _25502_);
  nor (_25516_, _25515_, _25514_);
  or (_25517_, _25516_, _14895_);
  nand (_25518_, _25516_, _14895_);
  and (_25519_, _25518_, _25517_);
  nor (_25520_, _25519_, _15221_);
  and (_25521_, _25519_, _15221_);
  nor (_25522_, _25521_, _25520_);
  not (_25524_, _25522_);
  or (_25525_, _25524_, _07591_);
  nand (_25526_, _07590_, _07427_);
  or (_25527_, _25526_, _25522_);
  and (_25528_, _25527_, _25525_);
  and (_25529_, _25528_, _25501_);
  or (_25530_, _25529_, _03441_);
  not (_25531_, _07407_);
  and (_25532_, _13682_, _25531_);
  or (_25533_, _25532_, _07408_);
  nor (_25535_, _25533_, _13983_);
  and (_25536_, _25533_, _13983_);
  nor (_25537_, _25536_, _25535_);
  and (_25538_, _25537_, _14207_);
  nor (_25539_, _25537_, _14207_);
  or (_25540_, _25539_, _25538_);
  and (_25541_, _14913_, _14588_);
  nor (_25542_, _14913_, _14588_);
  or (_25543_, _25542_, _25541_);
  and (_25544_, _25543_, _25540_);
  nor (_25546_, _25543_, _25540_);
  nor (_25547_, _25546_, _25544_);
  nor (_25548_, _25547_, _15141_);
  and (_25549_, _25547_, _15141_);
  nor (_25550_, _25549_, _25548_);
  and (_25551_, _25550_, _07417_);
  nor (_25552_, _25550_, _07417_);
  or (_25553_, _25552_, _25551_);
  or (_25554_, _25553_, _07344_);
  and (_25555_, _25554_, _02997_);
  and (_25557_, _25555_, _25530_);
  nand (_25558_, _13690_, _13344_);
  or (_25559_, _13690_, _13344_);
  and (_25560_, _25559_, _25558_);
  nor (_25561_, _25560_, _13884_);
  and (_25562_, _25560_, _13884_);
  nor (_25563_, _25562_, _25561_);
  nor (_25564_, _25563_, _14295_);
  and (_25565_, _25563_, _14295_);
  nor (_25566_, _25565_, _25564_);
  and (_25568_, _25566_, _14496_);
  nor (_25569_, _25566_, _14496_);
  or (_25570_, _25569_, _25568_);
  and (_25571_, _25570_, _14918_);
  nor (_25572_, _25570_, _14918_);
  nor (_25573_, _25572_, _25571_);
  nor (_25574_, _15124_, _07720_);
  and (_25575_, _15124_, _07720_);
  nor (_25576_, _25575_, _25574_);
  not (_25577_, _25576_);
  nand (_25579_, _25577_, _25573_);
  or (_25580_, _25577_, _25573_);
  and (_25581_, _25580_, _25579_);
  and (_25582_, _25581_, _02992_);
  or (_25583_, _25582_, _07276_);
  or (_25584_, _25583_, _25557_);
  nand (_25585_, _13595_, _13355_);
  or (_25586_, _13595_, _13355_);
  and (_25587_, _25586_, _25585_);
  and (_25588_, _25587_, _14000_);
  nor (_25590_, _25587_, _14000_);
  or (_25591_, _25590_, _25588_);
  nor (_25592_, _25591_, _14312_);
  and (_25593_, _25591_, _14312_);
  nor (_25594_, _25593_, _25592_);
  or (_25595_, _25594_, _14604_);
  nand (_25596_, _25594_, _14604_);
  and (_25597_, _25596_, _25595_);
  nor (_25598_, _25597_, _14816_);
  and (_25599_, _25597_, _14816_);
  or (_25601_, _25599_, _25598_);
  nor (_25602_, _25601_, _15238_);
  and (_25603_, _25601_, _15238_);
  nor (_25604_, _25603_, _25602_);
  not (_25605_, _25604_);
  nor (_25606_, _25605_, _07342_);
  and (_25607_, _25605_, _07342_);
  or (_25608_, _25607_, _25606_);
  or (_25609_, _25608_, _07277_);
  and (_25610_, _25609_, _25584_);
  or (_25612_, _25610_, _02585_);
  or (_25613_, _04635_, _04630_);
  nor (_25614_, _04701_, _04636_);
  and (_25615_, _25614_, _25613_);
  nor (_25616_, _25614_, _25613_);
  nor (_25617_, _25616_, _25615_);
  nor (_25618_, _04626_, _02933_);
  not (_25619_, _25618_);
  nor (_25620_, _04670_, _04663_);
  nor (_25621_, _25620_, _25619_);
  and (_25623_, _25620_, _25619_);
  nor (_25624_, _25623_, _25621_);
  or (_25625_, _25624_, _25617_);
  nand (_25626_, _25624_, _25617_);
  and (_25627_, _25626_, _25625_);
  or (_25628_, _25627_, _02586_);
  and (_25629_, _25628_, _02875_);
  and (_25630_, _25629_, _25612_);
  not (_25631_, _14320_);
  and (_25632_, _25631_, _14008_);
  nor (_25634_, _25631_, _14008_);
  nor (_25635_, _25634_, _25632_);
  nor (_25636_, _14929_, _14612_);
  and (_25637_, _14929_, _14612_);
  nor (_25638_, _25637_, _25636_);
  nor (_25639_, _25638_, _25635_);
  and (_25640_, _25638_, _25635_);
  nor (_25641_, _25640_, _25639_);
  and (_25642_, _13701_, _13423_);
  nor (_25643_, _13701_, _13423_);
  nor (_25645_, _25643_, _25642_);
  and (_25646_, _15247_, _07757_);
  nor (_25647_, _15247_, _07757_);
  nor (_25648_, _25647_, _25646_);
  not (_25649_, _25648_);
  and (_25650_, _25649_, _25645_);
  nor (_25651_, _25649_, _25645_);
  nor (_25652_, _25651_, _25650_);
  nand (_25653_, _25652_, _25641_);
  or (_25654_, _25652_, _25641_);
  and (_25656_, _25654_, _02874_);
  and (_25657_, _25656_, _25653_);
  or (_25658_, _25657_, _22922_);
  or (_25659_, _25658_, _25630_);
  nor (_25660_, _25070_, _22921_);
  nor (_25661_, _25660_, _06240_);
  and (_25662_, _25661_, _25659_);
  and (_25663_, _25386_, _06240_);
  nor (_25664_, _25663_, _25662_);
  nor (_25665_, _25664_, _06238_);
  and (_25667_, _25386_, _06238_);
  or (_25668_, _25667_, _02855_);
  or (_25669_, _25668_, _25665_);
  and (_25670_, _13709_, _13430_);
  nor (_25671_, _13709_, _13430_);
  nor (_25672_, _25671_, _25670_);
  not (_25673_, _25672_);
  not (_25674_, _14327_);
  and (_25675_, _25674_, _14015_);
  nor (_25676_, _25674_, _14015_);
  nor (_25677_, _25676_, _25675_);
  and (_25678_, _25677_, _25673_);
  nor (_25679_, _25677_, _25673_);
  nor (_25680_, _25679_, _25678_);
  not (_25681_, _14937_);
  and (_25682_, _25681_, _14619_);
  nor (_25683_, _25681_, _14619_);
  nor (_25684_, _25683_, _25682_);
  nand (_25685_, _25684_, _15255_);
  or (_25686_, _25684_, _15255_);
  and (_25689_, _25686_, _25685_);
  nor (_25690_, _25689_, _25680_);
  and (_25691_, _25689_, _25680_);
  or (_25692_, _25691_, _25690_);
  nor (_25693_, _25692_, _07764_);
  and (_25694_, _25692_, _07764_);
  or (_25695_, _25694_, _02856_);
  or (_25696_, _25695_, _25693_);
  and (_25697_, _25696_, _02851_);
  and (_25698_, _25697_, _25669_);
  and (_25700_, _13714_, _13435_);
  nor (_25701_, _13714_, _13435_);
  nor (_25702_, _25701_, _25700_);
  and (_25703_, _25702_, _14020_);
  nor (_25704_, _25702_, _14020_);
  or (_25705_, _25704_, _25703_);
  nand (_25706_, _25705_, _14332_);
  or (_25707_, _25705_, _14332_);
  and (_25708_, _25707_, _25706_);
  nor (_25709_, _15260_, _14942_);
  and (_25711_, _15260_, _14942_);
  nor (_25712_, _25711_, _25709_);
  not (_25713_, _14624_);
  and (_25714_, _25713_, _07769_);
  nor (_25715_, _25713_, _07769_);
  nor (_25716_, _25715_, _25714_);
  nor (_25717_, _25716_, _25712_);
  and (_25718_, _25716_, _25712_);
  nor (_25719_, _25718_, _25717_);
  or (_25720_, _25719_, _25708_);
  nand (_25722_, _25719_, _25708_);
  and (_25723_, _25722_, _02576_);
  and (_25724_, _25723_, _25720_);
  or (_25725_, _25724_, _06807_);
  or (_25726_, _25725_, _25698_);
  and (_25727_, _06864_, _15266_);
  nor (_25728_, _06864_, _15266_);
  nor (_25729_, _25728_, _25727_);
  nor (_25730_, _07004_, _06948_);
  and (_25731_, _07004_, _06948_);
  nor (_25733_, _25731_, _25730_);
  nor (_25734_, _25733_, _06894_);
  and (_25735_, _25733_, _06894_);
  nor (_25736_, _25735_, _25734_);
  nor (_25737_, _25736_, _25729_);
  and (_25738_, _25736_, _25729_);
  or (_25739_, _25738_, _25737_);
  nor (_25740_, _25739_, _07775_);
  and (_25741_, _25739_, _07775_);
  or (_25742_, _25741_, _25740_);
  and (_25744_, _25742_, _07069_);
  nor (_25745_, _25742_, _07069_);
  nor (_25746_, _25745_, _25744_);
  and (_25747_, _25746_, _07164_);
  nor (_25748_, _25746_, _07164_);
  or (_25749_, _25748_, _06813_);
  or (_25750_, _25749_, _25747_);
  and (_25751_, _25750_, _25726_);
  or (_25752_, _25751_, _02548_);
  or (_25753_, _25627_, _02584_);
  and (_25755_, _25753_, _09801_);
  and (_25756_, _25755_, _25752_);
  nand (_25757_, _25070_, _02938_);
  not (_25758_, _02516_);
  nor (_25759_, _02975_, _25758_);
  not (_25760_, _25759_);
  and (_25761_, _25760_, _22780_);
  nor (_25762_, _04144_, _10788_);
  nor (_25763_, _04110_, _02498_);
  nor (_25764_, _25763_, _25762_);
  not (_25766_, _25764_);
  and (_25767_, _25766_, _25761_);
  nand (_25768_, _25767_, _25757_);
  or (_25769_, _25768_, _25756_);
  and (_25770_, _02862_, _02516_);
  nor (_25771_, _25767_, _25070_);
  nor (_25772_, _25771_, _25770_);
  and (_25773_, _25772_, _25769_);
  and (_25774_, _25070_, _25770_);
  or (_25775_, _25774_, _03879_);
  or (_25777_, _25775_, _25773_);
  nand (_25778_, _25330_, _03879_);
  and (_25779_, _25778_, _03884_);
  and (_25780_, _25779_, _25777_);
  nor (_25781_, _14343_, _14031_);
  and (_25782_, _14343_, _14031_);
  nor (_25783_, _25782_, _25781_);
  nor (_25784_, _13725_, _13446_);
  and (_25785_, _13725_, _13446_);
  or (_25786_, _25785_, _25784_);
  nor (_25788_, _25786_, _25783_);
  and (_25789_, _25786_, _25783_);
  nor (_25790_, _25789_, _25788_);
  not (_25791_, _15275_);
  nor (_25792_, _14955_, _14635_);
  and (_25793_, _14955_, _14635_);
  nor (_25794_, _25793_, _25792_);
  nor (_25795_, _25794_, _25791_);
  and (_25796_, _25794_, _25791_);
  nor (_25797_, _25796_, _25795_);
  nor (_25799_, _25797_, _25790_);
  and (_25800_, _25797_, _25790_);
  or (_25801_, _25800_, _25799_);
  or (_25802_, _25801_, _07785_);
  nand (_25803_, _25801_, _07785_);
  and (_25804_, _25803_, _03014_);
  and (_25805_, _25804_, _25802_);
  or (_25806_, _25805_, _25780_);
  and (_25807_, _25806_, _07783_);
  nand (_25808_, _25627_, _07782_);
  nor (_25810_, _09400_, _09000_);
  and (_25811_, _25810_, _09438_);
  nand (_25812_, _25811_, _25808_);
  or (_25813_, _25812_, _25807_);
  or (_25814_, _25811_, _25070_);
  and (_25815_, _25814_, _07798_);
  and (_25816_, _25815_, _25813_);
  and (_25817_, _15119_, _07220_);
  nor (_25818_, _15119_, _07220_);
  nor (_25819_, _25818_, _25817_);
  and (_25821_, _13454_, _07241_);
  nor (_25822_, _25821_, _13958_);
  and (_25823_, _14179_, _07237_);
  nor (_25824_, _14179_, _07237_);
  nor (_25825_, _25824_, _25823_);
  nor (_25826_, _25825_, _25822_);
  and (_25827_, _25825_, _25822_);
  nor (_25828_, _25827_, _25826_);
  and (_25829_, _07230_, _07226_);
  nor (_25830_, _07230_, _07226_);
  nor (_25832_, _25830_, _25829_);
  nor (_25833_, _25832_, _25828_);
  and (_25834_, _25832_, _25828_);
  nor (_25835_, _25834_, _25833_);
  nor (_25836_, _25835_, _25819_);
  and (_25837_, _25835_, _25819_);
  or (_25838_, _25837_, _25836_);
  and (_25839_, _25838_, _07799_);
  or (_25840_, _25839_, _07802_);
  or (_25841_, _25840_, _25816_);
  not (_25843_, _08067_);
  and (_25844_, _25843_, _07808_);
  nor (_25845_, _25843_, _07808_);
  nor (_25846_, _25845_, _25844_);
  and (_25847_, _13340_, _08083_);
  nor (_25848_, _25847_, _13976_);
  nor (_25849_, _14198_, _08079_);
  and (_25850_, _14198_, _08079_);
  nor (_25851_, _25850_, _25849_);
  nor (_25852_, _25851_, _25848_);
  and (_25854_, _25851_, _25848_);
  nor (_25855_, _25854_, _25852_);
  nor (_25856_, _14797_, _08072_);
  and (_25857_, _14797_, _08072_);
  nor (_25858_, _25857_, _25856_);
  nor (_25859_, _25858_, _25855_);
  and (_25860_, _25858_, _25855_);
  nor (_25861_, _25860_, _25859_);
  nor (_25862_, _25861_, _25846_);
  and (_25863_, _25861_, _25846_);
  or (_25865_, _25863_, _25862_);
  or (_25866_, _25865_, _14491_);
  or (_25867_, _25865_, _20444_);
  and (_25868_, _25867_, _07814_);
  and (_25869_, _25868_, _25866_);
  and (_25870_, _25869_, _25841_);
  not (_25871_, _11769_);
  and (_25872_, _10739_, _10546_);
  nor (_25873_, _10739_, _10546_);
  or (_25874_, _25873_, _25872_);
  nor (_25875_, _11028_, _10831_);
  and (_25876_, _11028_, _10831_);
  nor (_25877_, _25876_, _25875_);
  and (_25878_, _25877_, _25874_);
  nor (_25879_, _25877_, _25874_);
  nor (_25880_, _25879_, _25878_);
  or (_25881_, _25880_, _11368_);
  nand (_25882_, _25880_, _11368_);
  and (_25883_, _25882_, _25881_);
  nor (_25884_, _25883_, _11436_);
  and (_25887_, _25883_, _11436_);
  or (_25888_, _25887_, _25884_);
  nand (_25889_, _25888_, _25871_);
  or (_25890_, _25888_, _25871_);
  and (_25891_, _25890_, _25889_);
  nor (_25892_, _25891_, _05771_);
  and (_25893_, _25891_, _05771_);
  or (_25894_, _25893_, _25892_);
  and (_25895_, _25894_, _03132_);
  or (_25896_, _25895_, _07812_);
  or (_25898_, _25896_, _25870_);
  and (_25899_, _08139_, _07820_);
  nor (_25900_, _25899_, _09322_);
  and (_25901_, _08142_, _08146_);
  nor (_25902_, _08142_, _08146_);
  or (_25903_, _25902_, _25901_);
  not (_25904_, _25903_);
  and (_25905_, _09319_, _08152_);
  nor (_25906_, _25905_, _09320_);
  not (_25907_, _25906_);
  and (_25909_, _09317_, _08156_);
  nor (_25910_, _25909_, _09318_);
  and (_25911_, _25910_, _25907_);
  nor (_25912_, _25910_, _25907_);
  nor (_25913_, _25912_, _25911_);
  nor (_25914_, _25913_, _25904_);
  and (_25915_, _25913_, _25904_);
  nor (_25916_, _25915_, _25914_);
  or (_25917_, _25916_, _25900_);
  nand (_25918_, _25916_, _25900_);
  and (_25920_, _25918_, _25917_);
  or (_25921_, _25920_, _07813_);
  and (_25922_, _25921_, _05279_);
  and (_25923_, _25922_, _25898_);
  nor (_25924_, _13753_, _13468_);
  and (_25925_, _13753_, _13468_);
  nor (_25926_, _25925_, _25924_);
  not (_25927_, _25926_);
  not (_25928_, _14191_);
  and (_25929_, _25928_, _14055_);
  nor (_25931_, _25928_, _14055_);
  nor (_25932_, _25931_, _25929_);
  and (_25933_, _25932_, _25927_);
  nor (_25934_, _25932_, _25927_);
  or (_25935_, _25934_, _25933_);
  nor (_25936_, _15113_, _14795_);
  and (_25937_, _15113_, _14795_);
  nor (_25938_, _25937_, _25936_);
  not (_25939_, _14489_);
  and (_25940_, _25939_, _07270_);
  nor (_25942_, _25939_, _07270_);
  nor (_25943_, _25942_, _25940_);
  nor (_25944_, _25943_, _25938_);
  and (_25945_, _25943_, _25938_);
  nor (_25946_, _25945_, _25944_);
  or (_25947_, _25946_, _25935_);
  nand (_25948_, _25946_, _25935_);
  and (_25949_, _25948_, _03021_);
  and (_25950_, _25949_, _25947_);
  or (_25951_, _25950_, _25923_);
  and (_25953_, _25951_, _03131_);
  nand (_25954_, _25070_, _03130_);
  or (_25955_, _25954_, _04712_);
  nand (_25956_, _25955_, _23634_);
  or (_25957_, _25956_, _25953_);
  and (_25958_, _13762_, _09471_);
  or (_25959_, _25070_, _23634_);
  and (_25960_, _25959_, _13581_);
  and (_25961_, _25960_, _25958_);
  and (_25962_, _25961_, _25957_);
  or (_25964_, _07242_, _07239_);
  nand (_25965_, _07242_, _07239_);
  and (_25966_, _25965_, _25964_);
  nor (_25967_, _07235_, _07234_);
  and (_25968_, _07235_, _07234_);
  nor (_25969_, _25968_, _25967_);
  not (_25970_, _25969_);
  and (_25971_, _25970_, _25966_);
  nor (_25972_, _25970_, _25966_);
  nor (_25973_, _25972_, _25971_);
  nor (_25975_, _07228_, _07224_);
  and (_25976_, _07228_, _07224_);
  nor (_25977_, _25976_, _25975_);
  and (_25978_, _07221_, _07219_);
  nor (_25979_, _25978_, _10204_);
  nor (_25980_, _25979_, _25977_);
  and (_25981_, _25979_, _25977_);
  nor (_25982_, _25981_, _25980_);
  or (_25983_, _25982_, _25973_);
  nand (_25984_, _25982_, _25973_);
  and (_25986_, _25984_, _25983_);
  and (_25987_, _25986_, _07827_);
  or (_25988_, _25987_, _03513_);
  or (_25989_, _25988_, _25962_);
  or (_25990_, _08084_, _08081_);
  nand (_25991_, _08084_, _08081_);
  and (_25992_, _25991_, _25990_);
  and (_25993_, _08076_, _08077_);
  nor (_25994_, _08076_, _08077_);
  nor (_25995_, _25994_, _25993_);
  and (_25997_, _25995_, _25992_);
  nor (_25998_, _25995_, _25992_);
  nor (_25999_, _25998_, _25997_);
  not (_26000_, _25999_);
  nor (_26001_, _08065_, _07266_);
  and (_26002_, _08065_, _07266_);
  nor (_26003_, _26002_, _26001_);
  nor (_26004_, _08068_, _08070_);
  and (_26005_, _08068_, _08070_);
  nor (_26006_, _26005_, _26004_);
  not (_26008_, _26006_);
  and (_26009_, _26008_, _26003_);
  nor (_26010_, _26008_, _26003_);
  nor (_26011_, _26010_, _26009_);
  nor (_26012_, _26011_, _26000_);
  and (_26013_, _26011_, _26000_);
  or (_26014_, _26013_, _07265_);
  or (_26015_, _26014_, _26012_);
  and (_26016_, _26015_, _25989_);
  or (_26017_, _26016_, _03141_);
  nor (_26019_, _10737_, _10545_);
  and (_26020_, _10737_, _10545_);
  nor (_26021_, _26020_, _26019_);
  not (_26022_, _26021_);
  not (_26023_, _11026_);
  and (_26024_, _26023_, _10829_);
  nor (_26025_, _26023_, _10829_);
  nor (_26026_, _26025_, _26024_);
  nor (_26027_, _26026_, _26022_);
  and (_26028_, _26026_, _26022_);
  nor (_26030_, _26028_, _26027_);
  not (_26031_, _11767_);
  nor (_26032_, _11434_, _11366_);
  and (_26033_, _11434_, _11366_);
  nor (_26034_, _26033_, _26032_);
  nor (_26035_, _26034_, _26031_);
  and (_26036_, _26034_, _26031_);
  nor (_26037_, _26036_, _26035_);
  not (_26038_, _26037_);
  nor (_26039_, _26038_, _26030_);
  and (_26041_, _26038_, _26030_);
  or (_26042_, _26041_, _26039_);
  and (_26043_, _26042_, _05769_);
  nor (_26044_, _26042_, _05769_);
  or (_26045_, _26044_, _26043_);
  or (_26046_, _26045_, _07838_);
  and (_26047_, _26046_, _07837_);
  and (_26048_, _26047_, _26017_);
  or (_26049_, _26048_, _25155_);
  and (_26050_, _26049_, _05274_);
  and (_26052_, _08877_, _08876_);
  nor (_26053_, _14079_, _13488_);
  and (_26054_, _14079_, _13488_);
  nor (_26055_, _26054_, _26053_);
  nor (_26056_, _15324_, _14683_);
  and (_26057_, _15324_, _14683_);
  nor (_26058_, _26057_, _26056_);
  and (_26059_, _26058_, _26055_);
  nor (_26060_, _26058_, _26055_);
  nor (_26061_, _26060_, _26059_);
  nor (_26063_, _14997_, _14382_);
  and (_26064_, _14997_, _14382_);
  nor (_26065_, _26064_, _26063_);
  nor (_26066_, _13779_, _07845_);
  and (_26067_, _13779_, _07845_);
  nor (_26068_, _26067_, _26066_);
  and (_26069_, _26068_, _26065_);
  nor (_26070_, _26068_, _26065_);
  nor (_26071_, _26070_, _26069_);
  not (_26072_, _26071_);
  nand (_26074_, _26072_, _26061_);
  or (_26075_, _26072_, _26061_);
  and (_26076_, _26075_, _03020_);
  nand (_26077_, _26076_, _26074_);
  nand (_26078_, _26077_, _26052_);
  or (_26079_, _26078_, _26050_);
  nand (_26080_, _03029_, _02537_);
  or (_26081_, _25070_, _26052_);
  and (_26082_, _26081_, _26080_);
  and (_26083_, _26082_, _26079_);
  nor (_26085_, _13453_, _07240_);
  and (_26086_, _13453_, _07240_);
  nor (_26087_, _26086_, _26085_);
  nor (_26088_, _07236_, _07232_);
  and (_26089_, _07236_, _07232_);
  nor (_26090_, _26089_, _26088_);
  and (_26091_, _26090_, _26087_);
  nor (_26092_, _26090_, _26087_);
  nor (_26093_, _26092_, _26091_);
  not (_26094_, _07225_);
  nor (_26096_, _07229_, _07222_);
  and (_26097_, _07229_, _07222_);
  nor (_26098_, _26097_, _26096_);
  nor (_26099_, _26098_, _26094_);
  and (_26100_, _26098_, _26094_);
  nor (_26101_, _26100_, _26099_);
  and (_26102_, _26101_, _26093_);
  nor (_26103_, _26101_, _26093_);
  or (_26104_, _26103_, _26102_);
  and (_26105_, _26104_, _07218_);
  nor (_26107_, _26104_, _07218_);
  or (_26108_, _26107_, _26105_);
  or (_26109_, _26108_, _02979_);
  and (_26110_, _26109_, _03360_);
  or (_26111_, _26110_, _26083_);
  not (_26112_, _03360_);
  or (_26113_, _26108_, _26112_);
  or (_26114_, _26113_, _02546_);
  and (_26115_, _26114_, _26111_);
  not (_26116_, _03715_);
  and (_26118_, _08870_, _26116_);
  and (_26119_, _26118_, _26115_);
  and (_26120_, _14648_, _02537_);
  not (_26121_, _26118_);
  and (_26122_, _26121_, _26108_);
  or (_26123_, _26122_, _26120_);
  or (_26124_, _26123_, _26119_);
  nor (_26125_, _13339_, _08082_);
  and (_26126_, _13339_, _08082_);
  nor (_26127_, _26126_, _26125_);
  not (_26129_, _26127_);
  and (_26130_, _08074_, _08078_);
  nor (_26131_, _08074_, _08078_);
  nor (_26132_, _26131_, _26130_);
  nor (_26133_, _26132_, _26129_);
  and (_26134_, _26132_, _26129_);
  nor (_26135_, _26134_, _26133_);
  not (_26136_, _08069_);
  nor (_26137_, _08071_, _08066_);
  and (_26138_, _08071_, _08066_);
  nor (_26140_, _26138_, _26137_);
  nor (_26141_, _26140_, _26136_);
  and (_26142_, _26140_, _26136_);
  nor (_26143_, _26142_, _26141_);
  not (_26144_, _26143_);
  nor (_26145_, _26144_, _26135_);
  and (_26146_, _26144_, _26135_);
  nor (_26147_, _26146_, _26145_);
  nand (_26148_, _26147_, _07807_);
  or (_26149_, _26147_, _07807_);
  and (_26151_, _26149_, _26148_);
  or (_26152_, _26151_, _08869_);
  and (_26153_, _26152_, _26124_);
  or (_26154_, _26153_, _03524_);
  not (_26155_, _03524_);
  or (_26156_, _26151_, _26155_);
  and (_26157_, _26156_, _03126_);
  and (_26158_, _26157_, _26154_);
  nor (_26159_, _10738_, _10421_);
  and (_26160_, _10738_, _10421_);
  nor (_26162_, _26160_, _26159_);
  and (_26163_, _26162_, _10830_);
  nor (_26164_, _26162_, _10830_);
  or (_26165_, _26164_, _26163_);
  nand (_26166_, _26165_, _11027_);
  or (_26167_, _26165_, _11027_);
  and (_26168_, _26167_, _26166_);
  nor (_26169_, _11435_, _11367_);
  and (_26170_, _11435_, _11367_);
  nor (_26171_, _26170_, _26169_);
  nor (_26173_, _26171_, _11768_);
  and (_26174_, _26171_, _11768_);
  nor (_26175_, _26174_, _26173_);
  and (_26176_, _26175_, _26168_);
  nor (_26177_, _26175_, _26168_);
  nor (_26178_, _26177_, _26176_);
  and (_26179_, _26178_, _05770_);
  nor (_26180_, _26178_, _05770_);
  or (_26181_, _26180_, _26179_);
  and (_26182_, _26181_, _03125_);
  or (_26184_, _26182_, _07865_);
  or (_26185_, _26184_, _26158_);
  nor (_26186_, _09316_, _08155_);
  and (_26187_, _09316_, _08155_);
  nor (_26188_, _26187_, _26186_);
  not (_26189_, _26188_);
  not (_26190_, _08149_);
  and (_26191_, _26190_, _08151_);
  nor (_26192_, _26190_, _08151_);
  nor (_26193_, _26192_, _26191_);
  nor (_26195_, _26193_, _26189_);
  and (_26196_, _26193_, _26189_);
  nor (_26197_, _26196_, _26195_);
  and (_26198_, _26197_, _08145_);
  nor (_26199_, _26197_, _08145_);
  or (_26200_, _26199_, _26198_);
  and (_26201_, _26200_, _08141_);
  nor (_26202_, _26200_, _08141_);
  or (_26203_, _26202_, _26201_);
  and (_26204_, _26203_, _08138_);
  nor (_26206_, _26203_, _08138_);
  or (_26207_, _26206_, _26204_);
  and (_26208_, _26207_, _07818_);
  nor (_26209_, _26207_, _07818_);
  or (_26210_, _26209_, _26208_);
  or (_26211_, _26210_, _07868_);
  and (_26212_, _26211_, _05781_);
  and (_26213_, _26212_, _26185_);
  or (_26214_, _26213_, _25129_);
  and (_26215_, _26214_, _25102_);
  or (_26217_, _25330_, _25102_);
  nand (_26218_, _26217_, _07889_);
  or (_26219_, _26218_, _26215_);
  nor (_26220_, _07577_, _07575_);
  nor (_26221_, _13800_, _25503_);
  nor (_26222_, _26221_, _26220_);
  nor (_26223_, _26222_, _14105_);
  and (_26224_, _26222_, _14105_);
  nor (_26225_, _26224_, _26223_);
  nor (_26226_, _26225_, _14185_);
  and (_26227_, _26225_, _14185_);
  or (_26228_, _26227_, _26226_);
  nor (_26229_, _26228_, _14705_);
  and (_26230_, _26228_, _14705_);
  or (_26231_, _26230_, _26229_);
  nor (_26232_, _26231_, _14787_);
  and (_26233_, _26231_, _14787_);
  or (_26234_, _26233_, _26232_);
  and (_26235_, _26234_, _15352_);
  nor (_26236_, _26234_, _15352_);
  or (_26239_, _26236_, _26235_);
  nand (_26240_, _26239_, _07913_);
  or (_26241_, _26239_, _07913_);
  and (_26242_, _26241_, _26240_);
  or (_26243_, _26242_, _07889_);
  and (_26244_, _26243_, _07922_);
  and (_26245_, _26244_, _26219_);
  not (_26246_, _14411_);
  nor (_26247_, _07407_, _07405_);
  nor (_26248_, _13577_, _25531_);
  nor (_26250_, _26248_, _26247_);
  nor (_26251_, _26250_, _14110_);
  and (_26252_, _26250_, _14110_);
  nor (_26253_, _26252_, _26251_);
  and (_26254_, _26253_, _26246_);
  nor (_26255_, _26253_, _26246_);
  nor (_26256_, _26255_, _26254_);
  and (_26257_, _26256_, _14482_);
  nor (_26258_, _26256_, _14482_);
  nor (_26259_, _26258_, _26257_);
  nor (_26261_, _26259_, _15029_);
  and (_26262_, _26259_, _15029_);
  or (_26263_, _26262_, _26261_);
  nor (_26264_, _26263_, _15357_);
  and (_26265_, _26263_, _15357_);
  or (_26266_, _26265_, _26264_);
  and (_26267_, _26266_, _07946_);
  nor (_26268_, _26266_, _07946_);
  or (_26269_, _26268_, _26267_);
  and (_26270_, _26269_, _07917_);
  or (_26272_, _26270_, _03137_);
  or (_26273_, _26272_, _26245_);
  and (_26274_, _26273_, _25101_);
  or (_26275_, _26274_, _07950_);
  not (_26276_, _08055_);
  nor (_26277_, _13812_, _13355_);
  and (_26278_, _13812_, _13355_);
  or (_26279_, _26278_, _26277_);
  nor (_26280_, _26279_, _14120_);
  and (_26281_, _26279_, _14120_);
  nor (_26283_, _26281_, _26280_);
  nor (_26284_, _26283_, _14421_);
  and (_26285_, _26283_, _14421_);
  or (_26286_, _26285_, _26284_);
  nor (_26287_, _26286_, _14718_);
  and (_26288_, _26286_, _14718_);
  or (_26289_, _26288_, _26287_);
  nor (_26290_, _26289_, _15040_);
  and (_26291_, _26289_, _15040_);
  or (_26292_, _26291_, _26290_);
  nor (_26294_, _26292_, _15365_);
  and (_26295_, _26292_, _15365_);
  or (_26296_, _26295_, _26294_);
  nor (_26297_, _26296_, _26276_);
  and (_26298_, _26296_, _26276_);
  or (_26299_, _26298_, _08031_);
  or (_26300_, _26299_, _26297_);
  and (_26301_, _26300_, _08030_);
  and (_26302_, _26301_, _26275_);
  nor (_26303_, _13589_, _13588_);
  nor (_26305_, _13911_, \oc8051_golden_model_1.ACC [3]);
  and (_26306_, _13911_, \oc8051_golden_model_1.ACC [3]);
  nor (_26307_, _26306_, _26305_);
  and (_26308_, _26307_, _25264_);
  nor (_26309_, _26307_, _25264_);
  nor (_26310_, _26309_, _26308_);
  not (_26311_, _26310_);
  nand (_26312_, _26311_, _26303_);
  or (_26313_, _26311_, _26303_);
  and (_26314_, _26313_, _26312_);
  nand (_26316_, _26314_, _08029_);
  nand (_26317_, _26316_, _25076_);
  or (_26318_, _26317_, _26302_);
  and (_26319_, _26318_, _25077_);
  or (_26320_, _26319_, _07258_);
  not (_26321_, _14726_);
  and (_26322_, _13495_, _07241_);
  nor (_26323_, _13495_, _07241_);
  nor (_26324_, _26323_, _26322_);
  and (_26325_, _26324_, _14127_);
  nor (_26327_, _26324_, _14127_);
  nor (_26328_, _26327_, _26325_);
  and (_26329_, _26328_, _14182_);
  nor (_26330_, _26328_, _14182_);
  or (_26331_, _26330_, _26329_);
  and (_26332_, _26331_, _26321_);
  nor (_26333_, _26331_, _26321_);
  nor (_26334_, _26333_, _26332_);
  and (_26335_, _26334_, _14784_);
  nor (_26336_, _26334_, _14784_);
  nor (_26337_, _26336_, _26335_);
  nor (_26338_, _26337_, _15374_);
  and (_26339_, _26337_, _15374_);
  or (_26340_, _26339_, _26338_);
  or (_26341_, _26340_, _07257_);
  nand (_26342_, _26340_, _07257_);
  and (_26343_, _26342_, _26341_);
  nor (_26344_, _26343_, _07259_);
  nor (_26345_, _26344_, _13341_);
  and (_26346_, _26345_, _26320_);
  not (_26349_, _13339_);
  and (_26350_, _26349_, _08083_);
  nor (_26351_, _26349_, _08083_);
  nor (_26352_, _26351_, _26350_);
  and (_26353_, _26352_, _14132_);
  nor (_26354_, _26352_, _14132_);
  nor (_26355_, _26354_, _26353_);
  and (_26356_, _26355_, _14432_);
  nor (_26357_, _26355_, _14432_);
  nor (_26358_, _26357_, _26356_);
  and (_26360_, _26358_, _14731_);
  nor (_26361_, _26358_, _14731_);
  nor (_26362_, _26361_, _26360_);
  nor (_26363_, _26362_, _15052_);
  and (_26364_, _26362_, _15052_);
  nor (_26365_, _26364_, _26363_);
  nor (_26366_, _26365_, _15379_);
  and (_26367_, _26365_, _15379_);
  or (_26368_, _26367_, _26366_);
  not (_26369_, _26368_);
  nor (_26371_, _26369_, _08099_);
  and (_26372_, _26369_, _08099_);
  or (_26373_, _26372_, _26371_);
  and (_26374_, _26373_, _13341_);
  or (_26375_, _26374_, _13541_);
  or (_26376_, _26375_, _26346_);
  not (_26377_, _13541_);
  or (_26378_, _26373_, _26377_);
  and (_26379_, _26378_, _02901_);
  and (_26380_, _26379_, _26376_);
  not (_26382_, _14137_);
  nor (_26383_, _13830_, _07734_);
  and (_26384_, _13830_, _07734_);
  or (_26385_, _26384_, _26383_);
  and (_26386_, _26385_, _26382_);
  nor (_26387_, _26385_, _26382_);
  nor (_26388_, _26387_, _26386_);
  and (_26389_, _26388_, _14438_);
  nor (_26390_, _26388_, _14438_);
  nor (_26391_, _26390_, _26389_);
  nor (_26393_, _26391_, _14737_);
  and (_26394_, _26391_, _14737_);
  or (_26395_, _26394_, _26393_);
  nor (_26396_, _26395_, _15058_);
  and (_26397_, _26395_, _15058_);
  or (_26398_, _26397_, _26396_);
  nor (_26399_, _26398_, _15385_);
  and (_26400_, _26398_, _15385_);
  nor (_26401_, _26400_, _26399_);
  or (_26402_, _26401_, _08131_);
  nand (_26404_, _26401_, _08131_);
  and (_26405_, _26404_, _02899_);
  and (_26406_, _26405_, _26402_);
  or (_26407_, _26406_, _26380_);
  and (_26408_, _26407_, _08106_);
  nor (_26409_, _13835_, _09317_);
  nor (_26410_, _26409_, _25909_);
  nor (_26411_, _26410_, _14140_);
  and (_26412_, _26410_, _14140_);
  or (_26413_, _26412_, _26411_);
  nor (_26415_, _26413_, _14444_);
  and (_26416_, _26413_, _14444_);
  nor (_26417_, _26416_, _26415_);
  and (_26418_, _26417_, _14740_);
  nor (_26419_, _26417_, _14740_);
  nor (_26420_, _26419_, _26418_);
  nor (_26421_, _26420_, _15063_);
  and (_26422_, _26420_, _15063_);
  or (_26423_, _26422_, _26421_);
  nor (_26424_, _26423_, _15390_);
  and (_26426_, _26423_, _15390_);
  or (_26427_, _26426_, _26424_);
  nand (_26428_, _26427_, _08172_);
  or (_26429_, _26427_, _08172_);
  and (_26430_, _26429_, _08103_);
  nand (_26431_, _26430_, _26428_);
  nand (_26432_, _26431_, _25073_);
  or (_26433_, _26432_, _26408_);
  nand (_26434_, _26433_, _25074_);
  nand (_26435_, _26434_, _11584_);
  nor (_26437_, _25070_, _11584_);
  nor (_26438_, _26437_, _03570_);
  and (_26439_, _26438_, _26435_);
  and (_26440_, _25070_, _03570_);
  or (_26441_, _26440_, _03909_);
  or (_26442_, _26441_, _26439_);
  nand (_26443_, _25330_, _03909_);
  and (_26444_, _26443_, _03563_);
  and (_26445_, _26444_, _26442_);
  and (_26446_, _25298_, _03166_);
  or (_26448_, _26446_, _08179_);
  or (_26449_, _26448_, _26445_);
  not (_26450_, _08185_);
  and (_26451_, _13911_, _26450_);
  and (_26452_, _26451_, \oc8051_golden_model_1.ACC [3]);
  nor (_26453_, _26451_, \oc8051_golden_model_1.ACC [3]);
  nor (_26454_, _26453_, _26452_);
  and (_26455_, _26454_, _14755_);
  nor (_26456_, _26454_, _14755_);
  nor (_26457_, _26456_, _26455_);
  and (_26459_, _15074_, _06833_);
  nor (_26460_, _15074_, _06833_);
  nor (_26461_, _26460_, _26459_);
  nor (_26462_, _26461_, _26457_);
  and (_26463_, _26461_, _26457_);
  or (_26464_, _26463_, _26462_);
  nor (_26465_, _26464_, _08191_);
  and (_26466_, _26464_, _08191_);
  nor (_26467_, _26466_, _26465_);
  nand (_26468_, _26467_, _08179_);
  and (_26470_, _26468_, _09787_);
  and (_26471_, _26470_, _26449_);
  and (_26472_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_26473_, _26472_, _07476_);
  or (_26474_, _26473_, _26310_);
  nand (_26475_, _26473_, _26310_);
  and (_26476_, _26475_, _26474_);
  nand (_26477_, _26476_, _08184_);
  nand (_26478_, _26477_, _03916_);
  or (_26479_, _26478_, _26471_);
  or (_26481_, _25070_, _03916_);
  and (_26482_, _26481_, _02501_);
  and (_26483_, _26482_, _26479_);
  and (_26484_, _25433_, _02500_);
  or (_26485_, _26484_, _09759_);
  or (_26486_, _26485_, _26483_);
  or (_26487_, _25070_, _09758_);
  and (_26488_, _26487_, _03178_);
  and (_26489_, _26488_, _26486_);
  not (_26490_, _14466_);
  nor (_26492_, _14767_, _26490_);
  and (_26493_, _14767_, _26490_);
  nor (_26494_, _26493_, _26492_);
  nor (_26495_, _26494_, _15414_);
  and (_26496_, _26494_, _15414_);
  nor (_26497_, _26496_, _26495_);
  not (_26498_, _26497_);
  nor (_26499_, _13854_, _13374_);
  and (_26500_, _13854_, _13374_);
  nor (_26501_, _26500_, _26499_);
  nor (_26503_, _26501_, _14164_);
  and (_26504_, _26501_, _14164_);
  nor (_26505_, _26504_, _26503_);
  and (_26506_, _26505_, _15088_);
  nor (_26507_, _26505_, _15088_);
  or (_26508_, _26507_, _26506_);
  and (_26509_, _26508_, _08204_);
  nor (_26510_, _26508_, _08204_);
  or (_26511_, _26510_, _26509_);
  nand (_26512_, _26511_, _26498_);
  or (_26514_, _26511_, _26498_);
  and (_26515_, _26514_, _03174_);
  and (_26516_, _26515_, _26512_);
  or (_26517_, _26516_, _26489_);
  and (_26518_, _26517_, _08202_);
  not (_26519_, _08209_);
  and (_26520_, _13911_, _26519_);
  and (_26521_, _26520_, _02701_);
  nor (_26522_, _26520_, _02701_);
  nor (_26523_, _26522_, _26521_);
  nor (_26525_, _26523_, _14773_);
  and (_26526_, _26523_, _14773_);
  or (_26527_, _26526_, _26525_);
  or (_26528_, _26527_, _15093_);
  nand (_26529_, _26527_, _15093_);
  and (_26530_, _26529_, _26528_);
  or (_26531_, _26530_, _15420_);
  nand (_26532_, _26530_, _15420_);
  and (_26533_, _26532_, _26531_);
  nor (_26534_, _26533_, _08216_);
  and (_26536_, _26533_, _08216_);
  or (_26537_, _26536_, _26534_);
  nand (_26538_, _26537_, _08201_);
  nor (_26539_, _09777_, _08208_);
  and (_26540_, _26539_, _19937_);
  nand (_26541_, _26540_, _26538_);
  or (_26542_, _26541_, _26518_);
  or (_26543_, _26540_, _25070_);
  and (_26544_, _26543_, _34698_);
  and (_26545_, _26544_, _26542_);
  or (_26547_, _26545_, _25055_);
  and (_35256_, _26547_, _36029_);
  nand (_26548_, _04709_, _03705_);
  or (_26549_, _04709_, \oc8051_golden_model_1.PSW [1]);
  and (_26550_, _26549_, _03014_);
  and (_26551_, _26550_, _26548_);
  nand (_26552_, _10720_, _04709_);
  and (_26553_, _26549_, _02576_);
  and (_26554_, _26553_, _26552_);
  and (_26555_, _10622_, _04709_);
  not (_26557_, _26555_);
  and (_26558_, _26557_, _26549_);
  or (_26559_, _26558_, _03821_);
  nand (_26560_, _04709_, _02618_);
  and (_26561_, _26560_, _26549_);
  and (_26562_, _26561_, _03825_);
  not (_26563_, \oc8051_golden_model_1.PSW [1]);
  nor (_26564_, _03825_, _26563_);
  or (_26565_, _26564_, _02952_);
  or (_26566_, _26565_, _26562_);
  and (_26568_, _26566_, _02892_);
  and (_26569_, _26568_, _26559_);
  and (_26570_, _10617_, _05329_);
  nor (_26571_, _05329_, _26563_);
  or (_26572_, _26571_, _02947_);
  or (_26573_, _26572_, _26570_);
  and (_26574_, _26573_, _09918_);
  or (_26575_, _26574_, _26569_);
  or (_26576_, _09802_, _04005_);
  and (_26577_, _26576_, _26549_);
  or (_26579_, _26577_, _03327_);
  and (_26580_, _26579_, _26575_);
  or (_26581_, _26580_, _02950_);
  or (_26582_, _26561_, _02959_);
  and (_26583_, _26582_, _02888_);
  and (_26584_, _26583_, _26581_);
  and (_26585_, _10620_, _05329_);
  or (_26586_, _26585_, _26571_);
  and (_26587_, _26586_, _02887_);
  or (_26588_, _26587_, _02880_);
  or (_26590_, _26588_, _26584_);
  and (_26591_, _26570_, _10616_);
  or (_26592_, _26571_, _02881_);
  or (_26593_, _26592_, _26591_);
  and (_26594_, _26593_, _26590_);
  and (_26595_, _26594_, _02875_);
  not (_26596_, _05329_);
  nor (_26597_, _10661_, _26596_);
  or (_26598_, _26571_, _26597_);
  and (_26599_, _26598_, _02874_);
  or (_26601_, _26599_, _06793_);
  or (_26602_, _26601_, _26595_);
  or (_26603_, _26577_, _06241_);
  and (_26604_, _26603_, _26602_);
  or (_26605_, _26604_, _02855_);
  or (_26606_, _06173_, _09802_);
  and (_26607_, _26606_, _26549_);
  or (_26608_, _26607_, _02856_);
  and (_26609_, _26608_, _02851_);
  and (_26610_, _26609_, _26605_);
  or (_26612_, _26610_, _26554_);
  and (_26613_, _26612_, _03884_);
  or (_26614_, _26613_, _26551_);
  and (_26615_, _26614_, _05279_);
  or (_26616_, _10612_, _09802_);
  and (_26617_, _26549_, _03021_);
  and (_26618_, _26617_, _26616_);
  or (_26619_, _26618_, _26615_);
  and (_26620_, _26619_, _03131_);
  or (_26621_, _10739_, _09802_);
  and (_26623_, _26549_, _03130_);
  and (_26624_, _26623_, _26621_);
  or (_26625_, _26624_, _26620_);
  and (_26626_, _26625_, _05274_);
  or (_26627_, _10611_, _09802_);
  and (_26628_, _26549_, _03020_);
  and (_26629_, _26628_, _26627_);
  or (_26630_, _26629_, _26626_);
  and (_26631_, _26630_, _03140_);
  nor (_26632_, _04709_, _26563_);
  or (_26634_, _26632_, _12724_);
  and (_26635_, _26561_, _03139_);
  and (_26636_, _26635_, _26634_);
  or (_26637_, _26636_, _26631_);
  and (_26638_, _26637_, _03128_);
  or (_26639_, _26548_, _12724_);
  and (_26640_, _26549_, _03036_);
  and (_26641_, _26640_, _26639_);
  or (_26642_, _26560_, _12724_);
  and (_26643_, _26549_, _03127_);
  and (_26645_, _26643_, _26642_);
  or (_26646_, _26645_, _03166_);
  or (_26647_, _26646_, _26641_);
  or (_26648_, _26647_, _26638_);
  or (_26649_, _26558_, _03563_);
  and (_26650_, _26649_, _02501_);
  and (_26651_, _26650_, _26648_);
  and (_26652_, _26586_, _02500_);
  or (_26653_, _26652_, _03174_);
  or (_26654_, _26653_, _26651_);
  or (_26656_, _26632_, _03178_);
  or (_26657_, _26656_, _26555_);
  and (_26658_, _26657_, _26654_);
  or (_26659_, _26658_, _34702_);
  or (_26660_, _34698_, \oc8051_golden_model_1.PSW [1]);
  and (_26661_, _26660_, _36029_);
  and (_35257_, _26661_, _26659_);
  and (_26662_, _07520_, \oc8051_golden_model_1.ACC [7]);
  nor (_26663_, _07520_, \oc8051_golden_model_1.ACC [7]);
  nor (_26664_, _26663_, _09794_);
  nor (_26666_, _26664_, _26662_);
  nand (_26667_, _26666_, _07913_);
  nand (_26668_, _26662_, _07910_);
  and (_26669_, _26668_, _26667_);
  and (_26670_, _26669_, _13517_);
  not (_26671_, \oc8051_golden_model_1.PSW [2]);
  nor (_26672_, _04709_, _26671_);
  not (_26673_, _26672_);
  and (_26674_, _26673_, _05142_);
  and (_26675_, _04709_, _05727_);
  nor (_26677_, _26675_, _26672_);
  or (_26678_, _26677_, _05274_);
  or (_26679_, _26678_, _26674_);
  nor (_26680_, _09802_, _04440_);
  nor (_26681_, _26680_, _26672_);
  and (_26682_, _26681_, _06793_);
  nor (_26683_, _05329_, _26671_);
  and (_26684_, _10838_, _05329_);
  or (_26685_, _26684_, _26683_);
  and (_26686_, _26685_, _02887_);
  nor (_26688_, _26681_, _03327_);
  and (_26689_, _10853_, _05329_);
  or (_26690_, _26689_, _26683_);
  or (_26691_, _26690_, _02892_);
  nor (_26692_, _10849_, _09802_);
  or (_26693_, _26692_, _26672_);
  and (_26694_, _26693_, _02952_);
  nor (_26695_, _03825_, _26671_);
  and (_26696_, _04709_, \oc8051_golden_model_1.ACC [2]);
  nor (_26697_, _26696_, _26672_);
  nor (_26699_, _26697_, _03826_);
  or (_26700_, _26699_, _26695_);
  and (_26701_, _26700_, _03821_);
  or (_26702_, _26701_, _02891_);
  or (_26703_, _26702_, _26694_);
  and (_26704_, _26703_, _26691_);
  and (_26705_, _26704_, _03327_);
  or (_26706_, _26705_, _26688_);
  or (_26707_, _26706_, _02950_);
  nand (_26708_, _26697_, _02950_);
  and (_26710_, _26708_, _02888_);
  and (_26711_, _26710_, _26707_);
  or (_26712_, _26711_, _26686_);
  and (_26713_, _26712_, _02881_);
  not (_26714_, _26683_);
  nand (_26715_, _26714_, _09820_);
  and (_26716_, _26690_, _02880_);
  and (_26717_, _26716_, _26715_);
  or (_26718_, _26717_, _26713_);
  and (_26719_, _26718_, _06277_);
  or (_26721_, _12677_, _12563_);
  or (_26722_, _26721_, _12795_);
  or (_26723_, _26722_, _12914_);
  or (_26724_, _26723_, _13031_);
  or (_26725_, _26724_, _13148_);
  or (_26726_, _26725_, _06789_);
  or (_26727_, _26726_, _13265_);
  and (_26728_, _26727_, _06271_);
  or (_26729_, _26728_, _07427_);
  or (_26730_, _26729_, _26719_);
  nor (_26732_, _26662_, _26663_);
  and (_26733_, _26732_, _10061_);
  nor (_26734_, _26732_, _10061_);
  nor (_26735_, _26734_, _26733_);
  nand (_26736_, _26735_, _07590_);
  or (_26737_, _26735_, _07590_);
  and (_26738_, _26737_, _26736_);
  or (_26739_, _26738_, _07426_);
  and (_26740_, _26739_, _26730_);
  and (_26741_, _26740_, _07344_);
  and (_26743_, _07345_, _05802_);
  not (_26744_, _26743_);
  and (_26745_, _26744_, _10076_);
  nor (_26746_, _26744_, _10076_);
  nor (_26747_, _26746_, _26745_);
  or (_26748_, _26747_, _07414_);
  nand (_26749_, _26747_, _07414_);
  and (_26750_, _26749_, _03441_);
  and (_26751_, _26750_, _26748_);
  or (_26752_, _26751_, _26741_);
  nand (_26754_, _26752_, _02997_);
  nor (_26755_, _10097_, _07971_);
  or (_26756_, _26755_, _07972_);
  nor (_26757_, _07962_, \oc8051_golden_model_1.ACC [7]);
  nor (_26758_, _07961_, _10218_);
  nor (_26759_, _26758_, _26757_);
  nor (_26760_, _26759_, _07967_);
  nor (_26761_, _10101_, _07963_);
  or (_26762_, _26761_, _26760_);
  and (_26763_, _26762_, _26756_);
  nor (_26765_, _26762_, _26756_);
  or (_26766_, _26765_, _02997_);
  or (_26767_, _26766_, _26763_);
  and (_26768_, _26767_, _07277_);
  and (_26769_, _26768_, _26754_);
  not (_26770_, _07283_);
  and (_26771_, _07339_, _26770_);
  not (_26772_, _26771_);
  nor (_26773_, _26772_, _10118_);
  and (_26774_, _26772_, _10118_);
  or (_26776_, _26774_, _26773_);
  and (_26777_, _26776_, _07276_);
  or (_26778_, _26777_, _02874_);
  or (_26779_, _26778_, _26769_);
  or (_26780_, _10886_, _26596_);
  and (_26781_, _26780_, _26714_);
  or (_26782_, _26781_, _02875_);
  and (_26783_, _26782_, _06241_);
  and (_26784_, _26783_, _26779_);
  or (_26785_, _26784_, _26682_);
  and (_26786_, _26785_, _02856_);
  or (_26787_, _06029_, _09802_);
  nor (_26788_, _26672_, _02856_);
  and (_26789_, _26788_, _26787_);
  or (_26790_, _26789_, _02576_);
  or (_26791_, _26790_, _26786_);
  or (_26792_, _10943_, _09802_);
  and (_26793_, _26792_, _26673_);
  or (_26794_, _26793_, _02851_);
  and (_26795_, _26794_, _06813_);
  and (_26798_, _26795_, _26791_);
  nor (_26799_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  nand (_26800_, _26799_, _06831_);
  and (_26801_, _26800_, _06807_);
  or (_26802_, _26801_, _26798_);
  and (_26803_, _26802_, _03884_);
  and (_26804_, _26677_, _03014_);
  or (_26805_, _26804_, _03021_);
  or (_26806_, _26805_, _26803_);
  nand (_26807_, _10835_, _04709_);
  and (_26809_, _26807_, _26673_);
  or (_26810_, _26809_, _05279_);
  and (_26811_, _26810_, _03131_);
  and (_26812_, _26811_, _26806_);
  nand (_26813_, _10831_, _04709_);
  nor (_26814_, _26672_, _03131_);
  and (_26815_, _26814_, _26813_);
  or (_26816_, _26815_, _03020_);
  or (_26817_, _26816_, _26812_);
  and (_26818_, _26817_, _26679_);
  or (_26820_, _26818_, _03139_);
  or (_26821_, _26697_, _03140_);
  or (_26822_, _26821_, _26674_);
  and (_26823_, _26822_, _05781_);
  and (_26824_, _26823_, _26820_);
  or (_26825_, _10833_, _09802_);
  and (_26826_, _26825_, _26673_);
  and (_26827_, _26826_, _03036_);
  or (_26828_, _26827_, _03127_);
  or (_26829_, _26828_, _26824_);
  or (_26831_, _10830_, _09802_);
  and (_26832_, _26831_, _26673_);
  or (_26833_, _26832_, _05786_);
  and (_26834_, _26833_, _13518_);
  and (_26835_, _26834_, _26829_);
  nor (_26836_, _26835_, _26670_);
  nor (_26837_, _26836_, _07886_);
  and (_26838_, _26669_, _07886_);
  or (_26839_, _26838_, _07917_);
  or (_26840_, _26839_, _26837_);
  nor (_26842_, _07345_, _10211_);
  or (_26843_, _07345_, _05802_);
  nand (_26844_, _26843_, _05768_);
  and (_26845_, _26844_, _10181_);
  nor (_26846_, _26845_, _26842_);
  nand (_26847_, _26846_, _07946_);
  nand (_26848_, _26842_, _07943_);
  and (_26849_, _26848_, _26847_);
  or (_26850_, _26849_, _07922_);
  and (_26851_, _26850_, _03138_);
  and (_26853_, _26851_, _26840_);
  and (_26854_, _26759_, _10188_);
  nor (_26855_, _26854_, _26758_);
  nand (_26856_, _26855_, _08025_);
  nand (_26857_, _26758_, _08022_);
  and (_26858_, _26857_, _03137_);
  and (_26859_, _26858_, _26856_);
  or (_26860_, _26859_, _26853_);
  and (_26861_, _26860_, _08031_);
  or (_26862_, _07282_, \oc8051_golden_model_1.ACC [7]);
  and (_26864_, _07282_, \oc8051_golden_model_1.ACC [7]);
  or (_26865_, _26864_, _10194_);
  and (_26866_, _26865_, _26862_);
  nand (_26867_, _26866_, _08055_);
  or (_26868_, _26866_, _08055_);
  and (_26869_, _26868_, _26867_);
  or (_26870_, _26869_, _08031_);
  nand (_26871_, _26870_, _07259_);
  or (_26872_, _26871_, _26861_);
  nor (_26873_, _07254_, _07218_);
  not (_26875_, _10204_);
  nor (_26876_, _26875_, _07253_);
  or (_26877_, _26876_, _07259_);
  or (_26878_, _26877_, _26873_);
  and (_26879_, _26878_, _08064_);
  nand (_26880_, _26879_, _26872_);
  and (_26881_, _08096_, _10211_);
  or (_26882_, _26881_, _10212_);
  nand (_26883_, _26882_, _07217_);
  and (_26884_, _26883_, _08104_);
  and (_26886_, _26884_, _26880_);
  or (_26887_, _08128_, _07598_);
  and (_26888_, _26887_, _10220_);
  not (_26889_, _25141_);
  or (_26890_, _26889_, _08168_);
  and (_26891_, _26890_, _08103_);
  and (_26892_, _26891_, _09788_);
  or (_26893_, _26892_, _03166_);
  or (_26894_, _26893_, _26888_);
  or (_26895_, _26894_, _26886_);
  or (_26897_, _26693_, _03563_);
  and (_26898_, _26897_, _02501_);
  and (_26899_, _26898_, _26895_);
  and (_26900_, _26685_, _02500_);
  or (_26901_, _26900_, _03174_);
  or (_26902_, _26901_, _26899_);
  and (_26903_, _11008_, _04709_);
  or (_26904_, _26672_, _03178_);
  or (_26905_, _26904_, _26903_);
  and (_26906_, _26905_, _26902_);
  or (_26908_, _26906_, _34702_);
  or (_26909_, _34698_, \oc8051_golden_model_1.PSW [2]);
  and (_26910_, _26909_, _36029_);
  and (_35258_, _26910_, _26908_);
  not (_26911_, \oc8051_golden_model_1.PSW [3]);
  nor (_26912_, _04709_, _26911_);
  nor (_26913_, _26912_, _04996_);
  not (_26914_, _26913_);
  and (_26915_, _04709_, _05664_);
  nor (_26916_, _26915_, _26912_);
  nor (_26918_, _26916_, _05274_);
  and (_26919_, _26918_, _26914_);
  nor (_26920_, _09802_, _04242_);
  nor (_26921_, _26920_, _26912_);
  and (_26922_, _26921_, _06793_);
  nor (_26923_, _05329_, _26911_);
  and (_26924_, _11035_, _05329_);
  nor (_26925_, _26924_, _26923_);
  nor (_26926_, _26925_, _02888_);
  and (_26927_, _04709_, \oc8051_golden_model_1.ACC [3]);
  nor (_26929_, _26927_, _26912_);
  nor (_26930_, _26929_, _03826_);
  nor (_26931_, _03825_, _26911_);
  or (_26932_, _26931_, _26930_);
  and (_26933_, _26932_, _03821_);
  nor (_26934_, _11040_, _09802_);
  nor (_26935_, _26934_, _26912_);
  nor (_26936_, _26935_, _03821_);
  or (_26937_, _26936_, _26933_);
  and (_26938_, _26937_, _02892_);
  and (_26940_, _11037_, _05329_);
  nor (_26941_, _26940_, _26923_);
  nor (_26942_, _26941_, _02892_);
  or (_26943_, _26942_, _02947_);
  or (_26944_, _26943_, _26938_);
  nand (_26945_, _26921_, _02947_);
  and (_26946_, _26945_, _26944_);
  and (_26947_, _26946_, _02959_);
  nor (_26948_, _26929_, _02959_);
  or (_26949_, _26948_, _26947_);
  and (_26952_, _26949_, _02888_);
  nor (_26953_, _26952_, _26926_);
  nor (_26954_, _26953_, _02880_);
  and (_26955_, _11067_, _05329_);
  nor (_26956_, _26955_, _26923_);
  nor (_26957_, _26956_, _02881_);
  nor (_26958_, _26957_, _26954_);
  nor (_26959_, _26958_, _02874_);
  nor (_26960_, _11083_, _26596_);
  nor (_26961_, _26960_, _26923_);
  nor (_26963_, _26961_, _02875_);
  nor (_26964_, _26963_, _06793_);
  not (_26965_, _26964_);
  nor (_26966_, _26965_, _26959_);
  nor (_26967_, _26966_, _26922_);
  nor (_26968_, _26967_, _02855_);
  and (_26969_, _06176_, _04709_);
  or (_26970_, _26912_, _02856_);
  nor (_26971_, _26970_, _26969_);
  nor (_26972_, _26971_, _26968_);
  and (_26974_, _26972_, _02851_);
  nor (_26975_, _11143_, _09802_);
  nor (_26976_, _26975_, _26912_);
  nor (_26977_, _26976_, _02851_);
  or (_26978_, _26977_, _26974_);
  and (_26979_, _26978_, _03884_);
  nor (_26980_, _26916_, _03884_);
  or (_26981_, _26980_, _26979_);
  and (_26982_, _26981_, _05279_);
  and (_26983_, _11032_, _04709_);
  nor (_26985_, _26983_, _26912_);
  nor (_26986_, _26985_, _05279_);
  or (_26987_, _26986_, _26982_);
  and (_26988_, _26987_, _03131_);
  and (_26989_, _11028_, _04709_);
  nor (_26990_, _26989_, _26912_);
  nor (_26991_, _26990_, _03131_);
  or (_26992_, _26991_, _26988_);
  and (_26993_, _26992_, _05274_);
  nor (_26994_, _26993_, _26919_);
  nor (_26996_, _26994_, _03139_);
  nor (_26997_, _26929_, _03140_);
  and (_26998_, _26997_, _26914_);
  or (_26999_, _26998_, _26996_);
  and (_27000_, _26999_, _05781_);
  nor (_27001_, _11030_, _09802_);
  nor (_27002_, _27001_, _26912_);
  nor (_27003_, _27002_, _05781_);
  or (_27004_, _27003_, _27000_);
  and (_27005_, _27004_, _05786_);
  nor (_27007_, _11027_, _09802_);
  nor (_27008_, _27007_, _26912_);
  nor (_27009_, _27008_, _05786_);
  or (_27010_, _27009_, _27005_);
  and (_27011_, _27010_, _03563_);
  nor (_27012_, _26935_, _03563_);
  or (_27013_, _27012_, _27011_);
  and (_27014_, _27013_, _02501_);
  nor (_27015_, _26925_, _02501_);
  or (_27016_, _27015_, _27014_);
  and (_27018_, _27016_, _03178_);
  and (_27019_, _11213_, _04709_);
  nor (_27020_, _27019_, _26912_);
  nor (_27021_, _27020_, _03178_);
  or (_27022_, _27021_, _27018_);
  or (_27023_, _27022_, _34702_);
  or (_27024_, _34698_, \oc8051_golden_model_1.PSW [3]);
  and (_27025_, _27024_, _36029_);
  and (_35259_, _27025_, _27023_);
  not (_27026_, \oc8051_golden_model_1.PSW [4]);
  nor (_27028_, _04709_, _27026_);
  nor (_27029_, _05202_, _09802_);
  nor (_27030_, _27029_, _27028_);
  and (_27031_, _27030_, _06793_);
  nor (_27032_, _05329_, _27026_);
  and (_27033_, _11243_, _05329_);
  nor (_27034_, _27033_, _27032_);
  nor (_27035_, _27034_, _02888_);
  and (_27036_, _04709_, \oc8051_golden_model_1.ACC [4]);
  nor (_27037_, _27036_, _27028_);
  nor (_27039_, _27037_, _03826_);
  nor (_27040_, _03825_, _27026_);
  or (_27041_, _27040_, _27039_);
  and (_27042_, _27041_, _03821_);
  nor (_27043_, _11259_, _09802_);
  nor (_27044_, _27043_, _27028_);
  nor (_27045_, _27044_, _03821_);
  or (_27046_, _27045_, _27042_);
  and (_27047_, _27046_, _02892_);
  and (_27048_, _11245_, _05329_);
  nor (_27050_, _27048_, _27032_);
  nor (_27051_, _27050_, _02892_);
  or (_27052_, _27051_, _02947_);
  or (_27053_, _27052_, _27047_);
  nand (_27054_, _27030_, _02947_);
  and (_27055_, _27054_, _27053_);
  and (_27056_, _27055_, _02959_);
  nor (_27057_, _27037_, _02959_);
  or (_27058_, _27057_, _27056_);
  and (_27059_, _27058_, _02888_);
  nor (_27061_, _27059_, _27035_);
  nor (_27062_, _27061_, _02880_);
  and (_27063_, _11277_, _05329_);
  nor (_27064_, _27063_, _27032_);
  nor (_27065_, _27064_, _02881_);
  nor (_27066_, _27065_, _27062_);
  nor (_27067_, _27066_, _02874_);
  nor (_27068_, _11241_, _26596_);
  nor (_27069_, _27068_, _27032_);
  nor (_27070_, _27069_, _02875_);
  nor (_27072_, _27070_, _06793_);
  not (_27073_, _27072_);
  nor (_27074_, _27073_, _27067_);
  nor (_27075_, _27074_, _27031_);
  nor (_27076_, _27075_, _02855_);
  and (_27077_, _06181_, _04709_);
  or (_27078_, _27028_, _02856_);
  nor (_27079_, _27078_, _27077_);
  nor (_27080_, _27079_, _27076_);
  and (_27081_, _27080_, _02851_);
  nor (_27082_, _11348_, _09802_);
  nor (_27083_, _27082_, _27028_);
  nor (_27084_, _27083_, _02851_);
  or (_27085_, _27084_, _27081_);
  and (_27086_, _27085_, _03884_);
  and (_27087_, _05697_, _04709_);
  nor (_27088_, _27087_, _27028_);
  nor (_27089_, _27088_, _03884_);
  or (_27090_, _27089_, _27086_);
  and (_27091_, _27090_, _05279_);
  and (_27094_, _11362_, _04709_);
  nor (_27095_, _27094_, _27028_);
  nor (_27096_, _27095_, _05279_);
  or (_27097_, _27096_, _27091_);
  and (_27098_, _27097_, _03131_);
  and (_27099_, _11368_, _04709_);
  nor (_27100_, _27099_, _27028_);
  nor (_27101_, _27100_, _03131_);
  or (_27102_, _27101_, _27098_);
  and (_27103_, _27102_, _05274_);
  nor (_27105_, _27028_, _05251_);
  not (_27106_, _27105_);
  nor (_27107_, _27088_, _05274_);
  and (_27108_, _27107_, _27106_);
  nor (_27109_, _27108_, _27103_);
  nor (_27110_, _27109_, _03139_);
  nor (_27111_, _27037_, _03140_);
  and (_27112_, _27111_, _27106_);
  or (_27113_, _27112_, _27110_);
  and (_27114_, _27113_, _05781_);
  nor (_27116_, _11361_, _09802_);
  nor (_27117_, _27116_, _27028_);
  nor (_27118_, _27117_, _05781_);
  or (_27119_, _27118_, _27114_);
  and (_27120_, _27119_, _05786_);
  nor (_27121_, _11367_, _09802_);
  nor (_27122_, _27121_, _27028_);
  nor (_27123_, _27122_, _05786_);
  or (_27124_, _27123_, _27120_);
  and (_27125_, _27124_, _03563_);
  nor (_27127_, _27044_, _03563_);
  or (_27128_, _27127_, _27125_);
  and (_27129_, _27128_, _02501_);
  nor (_27130_, _27034_, _02501_);
  or (_27131_, _27130_, _27129_);
  and (_27132_, _27131_, _03178_);
  and (_27133_, _11417_, _04709_);
  nor (_27134_, _27133_, _27028_);
  nor (_27135_, _27134_, _03178_);
  or (_27136_, _27135_, _27132_);
  or (_27138_, _27136_, _34702_);
  or (_27139_, _34698_, \oc8051_golden_model_1.PSW [4]);
  and (_27140_, _27139_, _36029_);
  and (_35260_, _27140_, _27138_);
  not (_27141_, \oc8051_golden_model_1.PSW [5]);
  nor (_27142_, _04709_, _27141_);
  nor (_27143_, _27142_, _04944_);
  not (_27144_, _27143_);
  and (_27145_, _05701_, _04709_);
  nor (_27146_, _27145_, _27142_);
  nor (_27148_, _27146_, _05274_);
  and (_27149_, _27148_, _27144_);
  nor (_27150_, _04896_, _09802_);
  nor (_27151_, _27150_, _27142_);
  and (_27152_, _27151_, _06793_);
  and (_27153_, _04709_, \oc8051_golden_model_1.ACC [5]);
  nor (_27154_, _27153_, _27142_);
  nor (_27155_, _27154_, _03826_);
  nor (_27156_, _03825_, _27141_);
  or (_27157_, _27156_, _27155_);
  and (_27159_, _27157_, _03821_);
  nor (_27160_, _11445_, _09802_);
  nor (_27161_, _27160_, _27142_);
  nor (_27162_, _27161_, _03821_);
  or (_27163_, _27162_, _27159_);
  and (_27164_, _27163_, _02892_);
  nor (_27165_, _05329_, _27141_);
  and (_27166_, _11459_, _05329_);
  nor (_27167_, _27166_, _27165_);
  nor (_27168_, _27167_, _02892_);
  or (_27170_, _27168_, _02947_);
  or (_27171_, _27170_, _27164_);
  nand (_27172_, _27151_, _02947_);
  and (_27173_, _27172_, _27171_);
  and (_27174_, _27173_, _02959_);
  nor (_27175_, _27154_, _02959_);
  or (_27176_, _27175_, _27174_);
  and (_27177_, _27176_, _02888_);
  and (_27178_, _11442_, _05329_);
  nor (_27179_, _27178_, _27165_);
  nor (_27181_, _27179_, _02888_);
  or (_27182_, _27181_, _02880_);
  or (_27183_, _27182_, _27177_);
  nor (_27184_, _27165_, _11474_);
  nor (_27185_, _27184_, _27167_);
  or (_27186_, _27185_, _02881_);
  and (_27187_, _27186_, _02875_);
  and (_27188_, _27187_, _27183_);
  nor (_27189_, _11440_, _26596_);
  nor (_27190_, _27189_, _27165_);
  nor (_27191_, _27190_, _02875_);
  nor (_27192_, _27191_, _06793_);
  not (_27193_, _27192_);
  nor (_27194_, _27193_, _27188_);
  nor (_27195_, _27194_, _27152_);
  nor (_27196_, _27195_, _02855_);
  and (_27197_, _06180_, _04709_);
  or (_27198_, _27142_, _02856_);
  nor (_27199_, _27198_, _27197_);
  nor (_27200_, _27199_, _27196_);
  and (_27203_, _27200_, _02851_);
  nor (_27204_, _11546_, _09802_);
  nor (_27205_, _27204_, _27142_);
  nor (_27206_, _27205_, _02851_);
  or (_27207_, _27206_, _27203_);
  and (_27208_, _27207_, _03884_);
  nor (_27209_, _27146_, _03884_);
  or (_27210_, _27209_, _27208_);
  and (_27211_, _27210_, _05279_);
  and (_27212_, _11562_, _04709_);
  nor (_27214_, _27212_, _27142_);
  nor (_27215_, _27214_, _05279_);
  or (_27216_, _27215_, _27211_);
  and (_27217_, _27216_, _03131_);
  and (_27218_, _11436_, _04709_);
  nor (_27219_, _27218_, _27142_);
  nor (_27220_, _27219_, _03131_);
  or (_27221_, _27220_, _27217_);
  and (_27222_, _27221_, _05274_);
  nor (_27223_, _27222_, _27149_);
  nor (_27225_, _27223_, _03139_);
  nor (_27226_, _27154_, _03140_);
  and (_27227_, _27226_, _27144_);
  or (_27228_, _27227_, _27225_);
  and (_27229_, _27228_, _05781_);
  nor (_27230_, _11560_, _09802_);
  nor (_27231_, _27230_, _27142_);
  nor (_27232_, _27231_, _05781_);
  or (_27233_, _27232_, _27229_);
  and (_27234_, _27233_, _05786_);
  nor (_27236_, _11435_, _09802_);
  nor (_27237_, _27236_, _27142_);
  nor (_27238_, _27237_, _05786_);
  or (_27239_, _27238_, _27234_);
  and (_27240_, _27239_, _03563_);
  nor (_27241_, _27161_, _03563_);
  or (_27242_, _27241_, _27240_);
  and (_27243_, _27242_, _02501_);
  nor (_27244_, _27179_, _02501_);
  or (_27245_, _27244_, _27243_);
  and (_27247_, _27245_, _03178_);
  and (_27248_, _11619_, _04709_);
  nor (_27249_, _27248_, _27142_);
  nor (_27250_, _27249_, _03178_);
  or (_27251_, _27250_, _27247_);
  or (_27252_, _27251_, _34702_);
  or (_27253_, _34698_, \oc8051_golden_model_1.PSW [5]);
  and (_27254_, _27253_, _36029_);
  and (_35261_, _27254_, _27252_);
  not (_27255_, _07538_);
  and (_27257_, _07904_, _27255_);
  nor (_27258_, _27257_, _07881_);
  nor (_27259_, _04709_, _14235_);
  nor (_27260_, _27259_, _04838_);
  not (_27261_, _27260_);
  and (_27262_, _11758_, _04709_);
  nor (_27263_, _27262_, _27259_);
  nor (_27264_, _27263_, _05274_);
  and (_27265_, _27264_, _27261_);
  nor (_27266_, _04787_, _09802_);
  nor (_27268_, _27266_, _27259_);
  and (_27269_, _27268_, _06793_);
  nor (_27270_, _05329_, _14235_);
  and (_27271_, _11653_, _05329_);
  or (_27272_, _27271_, _27270_);
  or (_27273_, _27270_, _11682_);
  and (_27274_, _27273_, _27272_);
  or (_27275_, _27274_, _02881_);
  nor (_27276_, _11636_, _09802_);
  nor (_27277_, _27276_, _27259_);
  nand (_27279_, _27277_, _02952_);
  and (_27280_, _04709_, \oc8051_golden_model_1.ACC [6]);
  nor (_27281_, _27280_, _27259_);
  nor (_27282_, _27281_, _03826_);
  nor (_27283_, _03825_, _14235_);
  or (_27284_, _27283_, _02952_);
  or (_27285_, _27284_, _27282_);
  and (_27286_, _27285_, _02892_);
  and (_27287_, _27286_, _27279_);
  and (_27288_, _27272_, _02891_);
  or (_27290_, _27288_, _02947_);
  or (_27291_, _27290_, _27287_);
  nand (_27292_, _27268_, _02947_);
  and (_27293_, _27292_, _27291_);
  or (_27294_, _27293_, _02950_);
  nand (_27295_, _27281_, _02950_);
  and (_27296_, _27295_, _02888_);
  and (_27297_, _27296_, _27294_);
  and (_27298_, _11675_, _05329_);
  nor (_27299_, _27298_, _27270_);
  nor (_27301_, _27299_, _02888_);
  or (_27302_, _27301_, _02880_);
  or (_27303_, _27302_, _27297_);
  and (_27304_, _27303_, _27275_);
  and (_27305_, _27304_, _07426_);
  or (_27306_, _07538_, _03441_);
  or (_27307_, _27306_, _07580_);
  and (_27308_, _27307_, _13666_);
  or (_27309_, _27308_, _27305_);
  or (_27310_, _07365_, _07344_);
  or (_27312_, _27310_, _07410_);
  and (_27313_, _27312_, _27309_);
  nor (_27314_, _27313_, _07597_);
  nor (_27315_, _07958_, _02997_);
  and (_27316_, _27315_, _10095_);
  nor (_27317_, _07279_, _07277_);
  and (_27318_, _27317_, _07333_);
  nor (_27319_, _27318_, _02874_);
  not (_27320_, _27319_);
  nor (_27321_, _27320_, _27316_);
  not (_27323_, _27321_);
  nor (_27324_, _27323_, _27314_);
  nor (_27325_, _11650_, _26596_);
  nor (_27326_, _27325_, _27270_);
  nor (_27327_, _27326_, _02875_);
  nor (_27328_, _27327_, _06793_);
  not (_27329_, _27328_);
  nor (_27330_, _27329_, _27324_);
  nor (_27331_, _27330_, _27269_);
  nor (_27332_, _27331_, _02855_);
  and (_27334_, _05847_, _04709_);
  or (_27335_, _27259_, _02856_);
  nor (_27336_, _27335_, _27334_);
  nor (_27337_, _27336_, _27332_);
  and (_27338_, _27337_, _02851_);
  nor (_27339_, _11751_, _09802_);
  nor (_27340_, _27339_, _27259_);
  nor (_27341_, _27340_, _02851_);
  or (_27342_, _27341_, _27338_);
  and (_27343_, _27342_, _03884_);
  nor (_27345_, _27263_, _03884_);
  or (_27346_, _27345_, _27343_);
  and (_27347_, _27346_, _05279_);
  and (_27348_, _11646_, _04709_);
  nor (_27349_, _27348_, _27259_);
  nor (_27350_, _27349_, _05279_);
  or (_27351_, _27350_, _27347_);
  and (_27352_, _27351_, _03131_);
  and (_27353_, _11769_, _04709_);
  nor (_27354_, _27353_, _27259_);
  nor (_27356_, _27354_, _03131_);
  or (_27357_, _27356_, _27352_);
  and (_27358_, _27357_, _05274_);
  nor (_27359_, _27358_, _27265_);
  nor (_27360_, _27359_, _03139_);
  nor (_27361_, _27281_, _03140_);
  and (_27362_, _27361_, _27261_);
  or (_27363_, _27362_, _27360_);
  and (_27364_, _27363_, _05781_);
  nor (_27365_, _11644_, _09802_);
  nor (_27367_, _27365_, _27259_);
  nor (_27368_, _27367_, _05781_);
  or (_27369_, _27368_, _27364_);
  nor (_27370_, _27369_, _03127_);
  not (_27371_, _07881_);
  nor (_27372_, _11768_, _09802_);
  nor (_27373_, _27259_, _05786_);
  not (_27374_, _27373_);
  nor (_27375_, _27374_, _27372_);
  nor (_27376_, _27375_, _27371_);
  not (_27378_, _27376_);
  nor (_27379_, _27378_, _27370_);
  nor (_27380_, _27379_, _27258_);
  nor (_27381_, _27380_, _07878_);
  not (_27382_, _27257_);
  and (_27383_, _27382_, _07878_);
  nor (_27384_, _27383_, _27381_);
  nor (_27385_, _27384_, _03535_);
  and (_27386_, _27382_, _03535_);
  nor (_27387_, _27386_, _27385_);
  nor (_27389_, _27387_, _07887_);
  nor (_27390_, _27257_, _13516_);
  or (_27391_, _27390_, _07886_);
  nor (_27392_, _27391_, _27389_);
  and (_27393_, _27257_, _07886_);
  or (_27394_, _27393_, _07917_);
  or (_27395_, _27394_, _27392_);
  not (_27396_, _07365_);
  and (_27397_, _07937_, _27396_);
  or (_27398_, _27397_, _07922_);
  and (_27400_, _27398_, _03138_);
  and (_27401_, _27400_, _27395_);
  nor (_27402_, _07958_, _03138_);
  and (_27403_, _27402_, _08016_);
  nor (_27404_, _27403_, _07950_);
  not (_27405_, _27404_);
  nor (_27406_, _27405_, _27401_);
  not (_27407_, _07279_);
  and (_27408_, _08046_, _27407_);
  or (_27409_, _27408_, _08031_);
  and (_27410_, _27409_, _07259_);
  not (_27411_, _27410_);
  nor (_27412_, _27411_, _27406_);
  nor (_27413_, _07259_, _07248_);
  or (_27414_, _27413_, _07217_);
  or (_27415_, _27414_, _27412_);
  nand (_27416_, _08090_, _07217_);
  and (_27417_, _27416_, _02901_);
  and (_27418_, _27417_, _27415_);
  nor (_27419_, _08122_, _02901_);
  or (_27422_, _27419_, _08103_);
  nor (_27423_, _27422_, _27418_);
  and (_27424_, _08163_, _08103_);
  or (_27425_, _27424_, _27423_);
  and (_27426_, _27425_, _03563_);
  nor (_27427_, _27277_, _03563_);
  or (_27428_, _27427_, _27426_);
  and (_27429_, _27428_, _02501_);
  nor (_27430_, _27299_, _02501_);
  or (_27431_, _27430_, _27429_);
  and (_27433_, _27431_, _03178_);
  and (_27434_, _11821_, _04709_);
  nor (_27435_, _27434_, _27259_);
  nor (_27436_, _27435_, _03178_);
  or (_27437_, _27436_, _27433_);
  or (_27438_, _27437_, _34702_);
  or (_27439_, _34698_, \oc8051_golden_model_1.PSW [6]);
  and (_27440_, _27439_, _36029_);
  and (_35262_, _27440_, _27438_);
  and (_35264_, \oc8051_golden_model_1.PCON [0], _36029_);
  and (_35265_, \oc8051_golden_model_1.PCON [1], _36029_);
  and (_35266_, \oc8051_golden_model_1.PCON [2], _36029_);
  and (_35267_, \oc8051_golden_model_1.PCON [3], _36029_);
  and (_35268_, \oc8051_golden_model_1.PCON [4], _36029_);
  and (_35269_, \oc8051_golden_model_1.PCON [5], _36029_);
  and (_35270_, \oc8051_golden_model_1.PCON [6], _36029_);
  and (_35271_, \oc8051_golden_model_1.SBUF [0], _36029_);
  and (_35272_, \oc8051_golden_model_1.SBUF [1], _36029_);
  and (_35273_, \oc8051_golden_model_1.SBUF [2], _36029_);
  and (_35275_, \oc8051_golden_model_1.SBUF [3], _36029_);
  and (_35276_, \oc8051_golden_model_1.SBUF [4], _36029_);
  and (_35277_, \oc8051_golden_model_1.SBUF [5], _36029_);
  and (_35278_, \oc8051_golden_model_1.SBUF [6], _36029_);
  and (_35279_, \oc8051_golden_model_1.SCON [0], _36029_);
  and (_35280_, \oc8051_golden_model_1.SCON [1], _36029_);
  and (_35281_, \oc8051_golden_model_1.SCON [2], _36029_);
  and (_35282_, \oc8051_golden_model_1.SCON [3], _36029_);
  and (_35283_, \oc8051_golden_model_1.SCON [4], _36029_);
  and (_35284_, \oc8051_golden_model_1.SCON [5], _36029_);
  and (_35286_, \oc8051_golden_model_1.SCON [6], _36029_);
  nor (_27444_, _04650_, _02877_);
  and (_27445_, _05044_, _04650_);
  nor (_27446_, _27445_, _27444_);
  and (_27447_, _27446_, _15506_);
  and (_27448_, _10546_, _04650_);
  nor (_27449_, _27448_, _27444_);
  nor (_27450_, _27449_, _03131_);
  not (_27451_, _27444_);
  and (_27452_, _06174_, _04650_);
  nor (_27453_, _27452_, _02856_);
  and (_27455_, _27453_, _27451_);
  not (_27456_, _27455_);
  and (_27457_, _04650_, \oc8051_golden_model_1.ACC [0]);
  nor (_27458_, _27457_, _27444_);
  nor (_27459_, _27458_, _03826_);
  nor (_27460_, _03825_, _02877_);
  or (_27461_, _27460_, _27459_);
  and (_27462_, _27461_, _03821_);
  nor (_27463_, _27446_, _03821_);
  or (_27464_, _27463_, _27462_);
  and (_27466_, _27464_, _03327_);
  or (_27467_, _27466_, _03410_);
  and (_27468_, _27467_, _02959_);
  nor (_27469_, _27458_, _02959_);
  or (_27470_, _27469_, _27468_);
  and (_27471_, _27470_, _03947_);
  nor (_27472_, _06793_, _03860_);
  not (_27473_, _27472_);
  nor (_27474_, _27473_, _27471_);
  and (_27475_, _04650_, _03817_);
  nor (_27477_, _27475_, _06241_);
  and (_27478_, _27477_, _27451_);
  nor (_27479_, _27478_, _27474_);
  nor (_27480_, _27479_, _02855_);
  nor (_27481_, _27480_, _02576_);
  and (_27482_, _27481_, _27456_);
  nor (_27483_, _10530_, _10307_);
  nor (_27484_, _27483_, _27444_);
  nor (_27485_, _27484_, _02851_);
  or (_27486_, _27485_, _27482_);
  and (_27488_, _27486_, _03884_);
  and (_27489_, _04650_, _05566_);
  nor (_27490_, _27489_, _27444_);
  nor (_27491_, _27490_, _03884_);
  or (_27492_, _27491_, _27488_);
  and (_27493_, _27492_, _05279_);
  and (_27494_, _10425_, _04650_);
  nor (_27495_, _27494_, _27444_);
  nor (_27496_, _27495_, _05279_);
  or (_27497_, _27496_, _27493_);
  and (_27499_, _27497_, _03131_);
  nor (_27500_, _27499_, _27450_);
  nor (_27501_, _27500_, _03020_);
  or (_27502_, _27490_, _05274_);
  nor (_27503_, _27502_, _27445_);
  nor (_27504_, _27503_, _27501_);
  nor (_27505_, _27504_, _03139_);
  and (_27506_, _10545_, _04650_);
  or (_27507_, _27506_, _27444_);
  and (_27508_, _27507_, _03139_);
  or (_27510_, _27508_, _27505_);
  and (_27511_, _27510_, _05781_);
  nor (_27512_, _10423_, _10307_);
  nor (_27513_, _27512_, _27444_);
  nor (_27514_, _27513_, _05781_);
  or (_27515_, _27514_, _27511_);
  and (_27516_, _27515_, _05786_);
  nor (_27517_, _10421_, _10307_);
  nor (_27518_, _27517_, _27444_);
  nor (_27519_, _27518_, _05786_);
  nor (_27521_, _27519_, _15506_);
  not (_27522_, _27521_);
  nor (_27523_, _27522_, _27516_);
  nor (_27524_, _27523_, _27447_);
  and (_27525_, _27524_, _34698_);
  nor (_27526_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27527_, _27526_, _00000_);
  or (_35287_, _27527_, _27525_);
  nor (_27528_, _04650_, _03937_);
  and (_27529_, _10622_, _04650_);
  nor (_27531_, _27529_, _27528_);
  nor (_27532_, _27531_, _03178_);
  not (_27533_, _25075_);
  not (_27534_, _03128_);
  and (_27535_, _02533_, _03937_);
  and (_27536_, _10739_, _04650_);
  or (_27537_, _27536_, _27528_);
  and (_27538_, _27537_, _03130_);
  and (_27539_, _02517_, _03937_);
  nor (_27540_, _10720_, _10307_);
  or (_27542_, _27540_, _27528_);
  and (_27543_, _27542_, _02576_);
  nor (_27544_, _04650_, \oc8051_golden_model_1.SP [1]);
  and (_27545_, _04650_, _02618_);
  nor (_27546_, _27545_, _27544_);
  nor (_27547_, _27546_, _03826_);
  nor (_27548_, _09213_, \oc8051_golden_model_1.SP [1]);
  and (_27549_, _02558_, \oc8051_golden_model_1.SP [1]);
  nor (_27550_, _27549_, _27548_);
  nor (_27551_, _27550_, _27547_);
  and (_27553_, _27551_, _03821_);
  nor (_27554_, _27544_, _27529_);
  and (_27555_, _27554_, _02952_);
  or (_27556_, _27555_, _27553_);
  and (_27557_, _27556_, _02556_);
  nor (_27558_, _02556_, \oc8051_golden_model_1.SP [1]);
  or (_27559_, _27558_, _02947_);
  or (_27560_, _27559_, _27557_);
  nand (_27561_, _03941_, _02947_);
  and (_27562_, _27561_, _27560_);
  and (_27564_, _27562_, _02959_);
  and (_27565_, _27546_, _02950_);
  or (_27566_, _27565_, _27564_);
  and (_27567_, _27566_, _03947_);
  or (_27568_, _27567_, _10292_);
  nor (_27569_, _27568_, _03946_);
  nor (_27570_, _04126_, _03937_);
  or (_27571_, _27570_, _06793_);
  nor (_27572_, _27571_, _27569_);
  or (_27573_, _10307_, _04005_);
  nor (_27575_, _27544_, _06241_);
  and (_27576_, _27575_, _27573_);
  nor (_27577_, _27576_, _02855_);
  not (_27578_, _27577_);
  nor (_27579_, _27578_, _27572_);
  not (_27580_, _27528_);
  and (_27581_, _06173_, _04650_);
  nor (_27582_, _27581_, _02856_);
  and (_27583_, _27582_, _27580_);
  nor (_27584_, _27583_, _02576_);
  not (_27586_, _27584_);
  nor (_27587_, _27586_, _27579_);
  nor (_27588_, _27587_, _27543_);
  nor (_27589_, _27588_, _03014_);
  and (_27590_, _04650_, _03705_);
  not (_27591_, _27590_);
  nor (_27592_, _27544_, _03884_);
  and (_27593_, _27592_, _27591_);
  or (_27594_, _27593_, _27589_);
  and (_27595_, _27594_, _04123_);
  or (_27597_, _27595_, _27539_);
  and (_27598_, _27597_, _05279_);
  nor (_27599_, _10612_, _10307_);
  or (_27600_, _27599_, _05279_);
  nor (_27601_, _27600_, _27544_);
  nor (_27602_, _27601_, _27598_);
  nor (_27603_, _27602_, _03130_);
  nor (_27604_, _27603_, _27538_);
  nor (_27605_, _27604_, _03020_);
  and (_27606_, _10611_, _04650_);
  or (_27608_, _27606_, _27528_);
  and (_27609_, _27608_, _03020_);
  nor (_27610_, _27609_, _27605_);
  nor (_27611_, _27610_, _10251_);
  and (_27612_, _27580_, _05095_);
  nor (_27613_, _27612_, _03140_);
  and (_27614_, _27613_, _27546_);
  or (_27615_, _27614_, _27611_);
  nor (_27616_, _27615_, _27535_);
  or (_27617_, _27616_, _27534_);
  and (_27619_, _27590_, _05095_);
  or (_27620_, _27619_, _05781_);
  nor (_27621_, _27620_, _27544_);
  nand (_27622_, _27545_, _05095_);
  nor (_27623_, _27544_, _05786_);
  and (_27624_, _27623_, _27622_);
  nor (_27625_, _27624_, _27621_);
  and (_27626_, _27625_, _27617_);
  nor (_27627_, _27626_, _27533_);
  nor (_27628_, _25075_, \oc8051_golden_model_1.SP [1]);
  nor (_27630_, _27628_, _02897_);
  not (_27631_, _27630_);
  nor (_27632_, _27631_, _27627_);
  nor (_27633_, _03739_, _03166_);
  not (_27634_, _27633_);
  nor (_27635_, _27634_, _27632_);
  and (_27636_, _27554_, _03166_);
  nor (_27637_, _27636_, _04159_);
  not (_27638_, _27637_);
  nor (_27639_, _27638_, _27635_);
  nor (_27641_, _03916_, _03937_);
  nor (_27642_, _27641_, _03174_);
  not (_27643_, _27642_);
  nor (_27644_, _27643_, _27639_);
  nor (_27645_, _27644_, _27532_);
  nor (_27646_, _27645_, _34702_);
  nor (_27647_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27648_, _27647_, _00000_);
  or (_35288_, _27648_, _27646_);
  and (_27649_, _04543_, _02531_);
  and (_27650_, _04543_, _02533_);
  nor (_27651_, _27650_, _03036_);
  nor (_27652_, _04650_, _03326_);
  and (_27653_, _10831_, _04650_);
  nor (_27654_, _27653_, _27652_);
  nor (_27655_, _27654_, _03131_);
  nor (_27656_, _10307_, _04440_);
  nor (_27657_, _27652_, _06241_);
  not (_27658_, _27657_);
  nor (_27659_, _27658_, _27656_);
  nor (_27662_, _12174_, _02561_);
  nor (_27663_, _10849_, _10307_);
  nor (_27664_, _27663_, _27652_);
  and (_27665_, _27664_, _02952_);
  and (_27666_, _04650_, \oc8051_golden_model_1.ACC [2]);
  nor (_27667_, _27666_, _27652_);
  or (_27668_, _27667_, _03826_);
  nand (_27669_, _09213_, \oc8051_golden_model_1.SP [2]);
  nor (_27670_, _12174_, _02558_);
  nor (_27671_, _27670_, _02952_);
  and (_27673_, _27671_, _27669_);
  and (_27674_, _27673_, _27668_);
  nor (_27675_, _27674_, _05382_);
  not (_27676_, _27675_);
  nor (_27677_, _27676_, _27665_);
  nor (_27678_, _12174_, _02556_);
  or (_27679_, _27678_, _02947_);
  nor (_27680_, _27679_, _27677_);
  and (_27681_, _05420_, _02947_);
  nor (_27682_, _27681_, _27680_);
  and (_27684_, _27682_, _02959_);
  nor (_27685_, _27667_, _02959_);
  or (_27686_, _27685_, _27684_);
  and (_27687_, _27686_, _03947_);
  or (_27688_, _27687_, _04369_);
  and (_27689_, _27688_, _02561_);
  or (_27690_, _27689_, _27662_);
  and (_27691_, _27690_, _05325_);
  and (_27692_, _04543_, _02578_);
  nor (_27693_, _27692_, _06793_);
  not (_27695_, _27693_);
  nor (_27696_, _27695_, _27691_);
  nor (_27697_, _27696_, _27659_);
  nor (_27698_, _27697_, _02855_);
  and (_27699_, _06177_, _04650_);
  or (_27700_, _27652_, _02856_);
  nor (_27701_, _27700_, _27699_);
  nor (_27702_, _27701_, _27698_);
  and (_27703_, _27702_, _02851_);
  nor (_27704_, _10943_, _10307_);
  nor (_27706_, _27704_, _27652_);
  nor (_27707_, _27706_, _02851_);
  or (_27708_, _27707_, _27703_);
  and (_27709_, _27708_, _03884_);
  and (_27710_, _04650_, _05727_);
  nor (_27711_, _27710_, _27652_);
  nor (_27712_, _27711_, _03884_);
  or (_27713_, _27712_, _02517_);
  or (_27714_, _27713_, _27709_);
  nand (_27715_, _12174_, _02517_);
  and (_27717_, _27715_, _27714_);
  and (_27718_, _27717_, _05279_);
  and (_27719_, _10835_, _04650_);
  nor (_27720_, _27719_, _27652_);
  nor (_27721_, _27720_, _05279_);
  or (_27722_, _27721_, _27718_);
  and (_27723_, _27722_, _03131_);
  nor (_27724_, _27723_, _27655_);
  nor (_27725_, _27724_, _03020_);
  nor (_27726_, _27652_, _05143_);
  not (_27728_, _27726_);
  nor (_27729_, _27711_, _05274_);
  and (_27730_, _27729_, _27728_);
  nor (_27731_, _27730_, _27725_);
  nor (_27732_, _27731_, _10251_);
  nor (_27733_, _27667_, _03140_);
  and (_27734_, _27733_, _27728_);
  nor (_27735_, _27734_, _27732_);
  and (_27736_, _27735_, _27651_);
  nor (_27737_, _10833_, _10307_);
  nor (_27739_, _27737_, _27652_);
  and (_27740_, _27739_, _03036_);
  nor (_27741_, _27740_, _27736_);
  and (_27742_, _27741_, _05786_);
  nor (_27743_, _10830_, _10307_);
  nor (_27744_, _27743_, _27652_);
  nor (_27745_, _27744_, _05786_);
  or (_27746_, _27745_, _27742_);
  and (_27747_, _27746_, _10250_);
  and (_27748_, _12174_, _03148_);
  or (_27750_, _27748_, _27747_);
  and (_27751_, _27750_, _05792_);
  or (_27752_, _27751_, _27649_);
  and (_27753_, _27752_, _02898_);
  and (_27754_, _12174_, _02897_);
  or (_27755_, _27754_, _03166_);
  nor (_27756_, _27755_, _27753_);
  and (_27757_, _27664_, _03166_);
  nor (_27758_, _27757_, _04159_);
  not (_27759_, _27758_);
  nor (_27761_, _27759_, _27756_);
  nor (_27762_, _12174_, _03916_);
  nor (_27763_, _27762_, _03174_);
  not (_27764_, _27763_);
  nor (_27765_, _27764_, _27761_);
  and (_27766_, _11008_, _04650_);
  nor (_27767_, _27766_, _27652_);
  and (_27768_, _27767_, _03174_);
  nor (_27769_, _27768_, _27765_);
  and (_27770_, _27769_, _34698_);
  nor (_27772_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27773_, _27772_, _00000_);
  or (_35290_, _27773_, _27770_);
  nor (_27774_, _04546_, _03916_);
  nor (_27775_, _04650_, _02946_);
  nor (_27776_, _27775_, _04996_);
  not (_27777_, _27776_);
  and (_27778_, _04650_, _05664_);
  nor (_27779_, _27778_, _27775_);
  nor (_27780_, _27779_, _05274_);
  and (_27782_, _27780_, _27777_);
  nor (_27783_, _04546_, _04126_);
  nor (_27784_, _11040_, _10307_);
  nor (_27785_, _27784_, _27775_);
  and (_27786_, _27785_, _02952_);
  and (_27787_, _04650_, \oc8051_golden_model_1.ACC [3]);
  nor (_27788_, _27787_, _27775_);
  or (_27789_, _27788_, _03826_);
  nand (_27790_, _09213_, \oc8051_golden_model_1.SP [3]);
  nor (_27791_, _11986_, _02558_);
  nor (_27793_, _27791_, _02952_);
  and (_27794_, _27793_, _27790_);
  and (_27795_, _27794_, _27789_);
  nor (_27796_, _27795_, _05382_);
  not (_27797_, _27796_);
  nor (_27798_, _27797_, _27786_);
  nor (_27799_, _11986_, _02556_);
  or (_27800_, _27799_, _02947_);
  nor (_27801_, _27800_, _27798_);
  and (_27802_, _05409_, _02947_);
  nor (_27804_, _27802_, _27801_);
  and (_27805_, _27804_, _02959_);
  nor (_27806_, _27788_, _02959_);
  or (_27807_, _27806_, _27805_);
  and (_27808_, _27807_, _03947_);
  or (_27809_, _27808_, _10292_);
  nor (_27810_, _27809_, _04291_);
  nor (_27811_, _27810_, _27783_);
  nor (_27812_, _27811_, _06793_);
  nor (_27813_, _10307_, _04242_);
  nor (_27815_, _27775_, _06241_);
  not (_27816_, _27815_);
  nor (_27817_, _27816_, _27813_);
  nor (_27818_, _27817_, _27812_);
  nor (_27819_, _27818_, _02855_);
  and (_27820_, _06176_, _04650_);
  nor (_27821_, _27775_, _02856_);
  not (_27822_, _27821_);
  nor (_27823_, _27822_, _27820_);
  nor (_27824_, _27823_, _27819_);
  nor (_27826_, _27824_, _02576_);
  nor (_27827_, _11143_, _10307_);
  nor (_27828_, _27827_, _27775_);
  and (_27829_, _27828_, _02576_);
  nor (_27830_, _27829_, _27826_);
  and (_27831_, _27830_, _03884_);
  nor (_27832_, _27779_, _03884_);
  or (_27833_, _27832_, _27831_);
  and (_27834_, _27833_, _04123_);
  and (_27835_, _04546_, _02517_);
  or (_27837_, _27835_, _27834_);
  and (_27838_, _27837_, _05279_);
  and (_27839_, _11032_, _04650_);
  nor (_27840_, _27839_, _27775_);
  nor (_27841_, _27840_, _05279_);
  or (_27842_, _27841_, _27838_);
  and (_27843_, _27842_, _03131_);
  and (_27844_, _11028_, _04650_);
  nor (_27845_, _27844_, _27775_);
  nor (_27846_, _27845_, _03131_);
  or (_27848_, _27846_, _27843_);
  and (_27849_, _27848_, _05274_);
  nor (_27850_, _27849_, _27782_);
  nor (_27851_, _27850_, _10251_);
  and (_27852_, _04546_, _02533_);
  or (_27853_, _27776_, _03140_);
  nor (_27854_, _27853_, _27788_);
  nor (_27855_, _27854_, _27852_);
  and (_27856_, _27855_, _05781_);
  not (_27857_, _27856_);
  nor (_27859_, _27857_, _27851_);
  nor (_27860_, _11030_, _10307_);
  or (_27861_, _27775_, _05781_);
  nor (_27862_, _27861_, _27860_);
  nor (_27863_, _27862_, _27859_);
  and (_27864_, _27863_, _05786_);
  nor (_27865_, _11027_, _10307_);
  nor (_27866_, _27865_, _27775_);
  nor (_27867_, _27866_, _05786_);
  or (_27868_, _27867_, _27864_);
  and (_27870_, _27868_, _10250_);
  nor (_27871_, _05406_, _02946_);
  nor (_27872_, _27871_, _05407_);
  nor (_27873_, _27872_, _10250_);
  or (_27874_, _27873_, _02531_);
  nor (_27875_, _27874_, _27870_);
  and (_27876_, _11986_, _02531_);
  nor (_27877_, _27876_, _27875_);
  and (_27878_, _27877_, _02898_);
  nor (_27879_, _27872_, _02898_);
  or (_27881_, _27879_, _27878_);
  and (_27882_, _27881_, _03563_);
  nor (_27883_, _27785_, _03563_);
  nor (_27884_, _27883_, _04159_);
  not (_27885_, _27884_);
  nor (_27886_, _27885_, _27882_);
  nor (_27887_, _27886_, _27774_);
  nor (_27888_, _27887_, _03174_);
  and (_27889_, _11213_, _04650_);
  nor (_27890_, _27889_, _27775_);
  and (_27892_, _27890_, _03174_);
  nor (_27893_, _27892_, _27888_);
  or (_27894_, _27893_, _34702_);
  or (_27895_, _34698_, \oc8051_golden_model_1.SP [3]);
  and (_27896_, _27895_, _36029_);
  and (_35291_, _27896_, _27894_);
  nor (_27897_, _04248_, \oc8051_golden_model_1.SP [4]);
  nor (_27898_, _27897_, _10243_);
  nor (_27899_, _27898_, _03916_);
  nor (_27900_, _04650_, _10278_);
  and (_27902_, _11368_, _04650_);
  nor (_27903_, _27902_, _27900_);
  nor (_27904_, _27903_, _03131_);
  nor (_27905_, _05202_, _10307_);
  or (_27906_, _27900_, _02855_);
  or (_27907_, _27906_, _27905_);
  and (_27908_, _27907_, _20391_);
  nor (_27909_, _11259_, _10307_);
  nor (_27910_, _27909_, _27900_);
  and (_27911_, _27910_, _02952_);
  and (_27913_, _04650_, \oc8051_golden_model_1.ACC [4]);
  nor (_27914_, _27913_, _27900_);
  or (_27915_, _27914_, _03826_);
  nand (_27916_, _09213_, \oc8051_golden_model_1.SP [4]);
  not (_27917_, _27898_);
  nor (_27918_, _27917_, _02558_);
  nor (_27919_, _27918_, _02952_);
  and (_27920_, _27919_, _27916_);
  and (_27921_, _27920_, _27915_);
  nor (_27922_, _27921_, _05382_);
  not (_27924_, _27922_);
  nor (_27925_, _27924_, _27911_);
  nor (_27926_, _27917_, _02556_);
  or (_27927_, _27926_, _02947_);
  nor (_27928_, _27927_, _27925_);
  and (_27929_, _10279_, _02877_);
  nor (_27930_, _05408_, _10278_);
  nor (_27931_, _27930_, _27929_);
  and (_27932_, _27931_, _02947_);
  nor (_27933_, _27932_, _27928_);
  and (_27934_, _27933_, _02959_);
  nor (_27935_, _27914_, _02959_);
  or (_27936_, _27935_, _27934_);
  and (_27937_, _27936_, _03947_);
  nor (_27938_, _04249_, _10278_);
  and (_27939_, _04249_, _10278_);
  nor (_27940_, _27939_, _27938_);
  and (_27941_, _27940_, _02886_);
  nor (_27942_, _27941_, _10292_);
  not (_27943_, _27942_);
  nor (_27945_, _27943_, _27937_);
  nor (_27946_, _27898_, _04126_);
  or (_27947_, _27946_, _06793_);
  nor (_27948_, _27947_, _27945_);
  nor (_27949_, _27948_, _27908_);
  and (_27950_, _06181_, _04650_);
  nor (_27951_, _27900_, _02856_);
  not (_27952_, _27951_);
  nor (_27953_, _27952_, _27950_);
  or (_27954_, _27953_, _02576_);
  nor (_27956_, _27954_, _27949_);
  nor (_27957_, _11348_, _10307_);
  nor (_27958_, _27957_, _27900_);
  nor (_27959_, _27958_, _02851_);
  or (_27960_, _27959_, _03014_);
  or (_27961_, _27960_, _27956_);
  and (_27962_, _05697_, _04650_);
  nor (_27963_, _27962_, _27900_);
  nand (_27964_, _27963_, _03014_);
  and (_27965_, _27964_, _27961_);
  nor (_27967_, _27965_, _02517_);
  and (_27968_, _27917_, _02517_);
  nor (_27969_, _27968_, _27967_);
  and (_27970_, _27969_, _05279_);
  and (_27971_, _11362_, _04650_);
  nor (_27972_, _27971_, _27900_);
  nor (_27973_, _27972_, _05279_);
  or (_27974_, _27973_, _27970_);
  and (_27975_, _27974_, _03131_);
  nor (_27976_, _27975_, _27904_);
  nor (_27978_, _27976_, _03020_);
  nor (_27979_, _27900_, _05251_);
  not (_27980_, _27979_);
  nor (_27981_, _27963_, _05274_);
  and (_27982_, _27981_, _27980_);
  nor (_27983_, _27982_, _27978_);
  nor (_27984_, _27983_, _10251_);
  nor (_27985_, _27914_, _03140_);
  and (_27986_, _27985_, _27980_);
  and (_27987_, _27898_, _02533_);
  nor (_27989_, _27987_, _27986_);
  and (_27990_, _27989_, _05781_);
  not (_27991_, _27990_);
  nor (_27992_, _27991_, _27984_);
  nor (_27993_, _11361_, _10307_);
  or (_27994_, _27900_, _05781_);
  nor (_27995_, _27994_, _27993_);
  nor (_27996_, _27995_, _27992_);
  and (_27997_, _27996_, _05786_);
  nor (_27998_, _11367_, _10307_);
  nor (_28000_, _27998_, _27900_);
  nor (_28001_, _28000_, _05786_);
  or (_28002_, _28001_, _27997_);
  and (_28003_, _28002_, _10250_);
  nor (_28004_, _05407_, _10278_);
  nor (_28005_, _28004_, _10279_);
  nor (_28006_, _28005_, _10250_);
  or (_28007_, _28006_, _02531_);
  nor (_28008_, _28007_, _28003_);
  and (_28009_, _27917_, _02531_);
  nor (_28011_, _28009_, _28008_);
  and (_28012_, _28011_, _02898_);
  nor (_28013_, _28005_, _02898_);
  or (_28014_, _28013_, _28012_);
  and (_28015_, _28014_, _03563_);
  nor (_28016_, _27910_, _03563_);
  nor (_28017_, _28016_, _04159_);
  not (_28018_, _28017_);
  nor (_28019_, _28018_, _28015_);
  nor (_28020_, _28019_, _27899_);
  and (_28022_, _28020_, _03178_);
  and (_28023_, _11417_, _04650_);
  nor (_28024_, _28023_, _27900_);
  nor (_28025_, _28024_, _03178_);
  or (_28026_, _28025_, _28022_);
  or (_28027_, _28026_, _34702_);
  or (_28028_, _34698_, \oc8051_golden_model_1.SP [4]);
  and (_28029_, _28028_, _36029_);
  and (_35292_, _28029_, _28027_);
  nor (_28030_, _10243_, \oc8051_golden_model_1.SP [5]);
  nor (_28032_, _28030_, _10244_);
  nor (_28033_, _28032_, _03916_);
  nor (_28034_, _04650_, _10277_);
  nor (_28035_, _28034_, _04944_);
  not (_28036_, _28035_);
  and (_28037_, _05701_, _04650_);
  nor (_28038_, _28037_, _28034_);
  nor (_28039_, _28038_, _05274_);
  and (_28040_, _28039_, _28036_);
  nor (_28041_, _11546_, _10307_);
  or (_28043_, _28034_, _02851_);
  nor (_28044_, _28043_, _28041_);
  nor (_28045_, _28032_, _04126_);
  nor (_28046_, _11445_, _10307_);
  nor (_28047_, _28046_, _28034_);
  and (_28048_, _28047_, _02952_);
  and (_28049_, _04650_, \oc8051_golden_model_1.ACC [5]);
  nor (_28050_, _28049_, _28034_);
  or (_28051_, _28050_, _03826_);
  nand (_28052_, _09213_, \oc8051_golden_model_1.SP [5]);
  and (_28054_, _28032_, _03824_);
  nor (_28055_, _28054_, _02952_);
  and (_28056_, _28055_, _28052_);
  and (_28057_, _28056_, _28051_);
  nor (_28058_, _28057_, _05382_);
  not (_28059_, _28058_);
  nor (_28060_, _28059_, _28048_);
  or (_28061_, _28032_, _02947_);
  and (_28062_, _28061_, _22787_);
  nor (_28063_, _28062_, _28060_);
  and (_28065_, _10280_, _02877_);
  nor (_28066_, _27929_, _10277_);
  nor (_28067_, _28066_, _28065_);
  and (_28068_, _28067_, _02947_);
  nor (_28069_, _28068_, _28063_);
  and (_28070_, _28069_, _02959_);
  nor (_28071_, _28050_, _02959_);
  or (_28072_, _28071_, _28070_);
  and (_28073_, _28072_, _03947_);
  and (_28074_, _10244_, \oc8051_golden_model_1.SP [0]);
  nor (_28076_, _27938_, \oc8051_golden_model_1.SP [5]);
  nor (_28077_, _28076_, _28074_);
  and (_28078_, _28077_, _02886_);
  nor (_28079_, _28078_, _10292_);
  not (_28080_, _28079_);
  nor (_28081_, _28080_, _28073_);
  nor (_28082_, _28081_, _28045_);
  nor (_28083_, _28082_, _06793_);
  nor (_28084_, _04896_, _10307_);
  nor (_28085_, _28034_, _06241_);
  not (_28087_, _28085_);
  nor (_28088_, _28087_, _28084_);
  nor (_28089_, _28088_, _28083_);
  nor (_28090_, _28089_, _02855_);
  and (_28091_, _06180_, _04650_);
  nor (_28092_, _28034_, _02856_);
  not (_28093_, _28092_);
  nor (_28094_, _28093_, _28091_);
  nor (_28095_, _28094_, _28090_);
  nor (_28096_, _28095_, _02576_);
  nor (_28098_, _28096_, _28044_);
  and (_28099_, _28098_, _03884_);
  nor (_28100_, _28038_, _03884_);
  or (_28101_, _28100_, _28099_);
  and (_28102_, _28101_, _04123_);
  and (_28103_, _28032_, _02517_);
  or (_28104_, _28103_, _28102_);
  and (_28105_, _28104_, _05279_);
  and (_28106_, _11562_, _04650_);
  nor (_28107_, _28106_, _28034_);
  nor (_28109_, _28107_, _05279_);
  or (_28110_, _28109_, _28105_);
  and (_28111_, _28110_, _03131_);
  and (_28112_, _11436_, _04650_);
  nor (_28113_, _28112_, _28034_);
  nor (_28114_, _28113_, _03131_);
  or (_28115_, _28114_, _28111_);
  and (_28116_, _28115_, _05274_);
  nor (_28117_, _28116_, _28040_);
  nor (_28118_, _28117_, _10251_);
  nor (_28120_, _28050_, _03140_);
  and (_28121_, _28120_, _28036_);
  and (_28122_, _28032_, _02533_);
  nor (_28123_, _28122_, _28121_);
  and (_28124_, _28123_, _05781_);
  not (_28125_, _28124_);
  nor (_28126_, _28125_, _28118_);
  nor (_28127_, _11560_, _10307_);
  or (_28128_, _28034_, _05781_);
  nor (_28129_, _28128_, _28127_);
  nor (_28131_, _28129_, _28126_);
  and (_28132_, _28131_, _05786_);
  nor (_28133_, _11435_, _10307_);
  nor (_28134_, _28133_, _28034_);
  nor (_28135_, _28134_, _05786_);
  or (_28136_, _28135_, _28132_);
  and (_28137_, _28136_, _10250_);
  nor (_28138_, _10279_, _10277_);
  nor (_28139_, _28138_, _10280_);
  nor (_28140_, _28139_, _10250_);
  or (_28142_, _28140_, _02531_);
  nor (_28143_, _28142_, _28137_);
  nor (_28144_, _28032_, _05792_);
  nor (_28145_, _28144_, _28143_);
  and (_28146_, _28145_, _02898_);
  nor (_28147_, _28139_, _02898_);
  or (_28148_, _28147_, _28146_);
  and (_28149_, _28148_, _03563_);
  nor (_28150_, _28047_, _03563_);
  nor (_28151_, _28150_, _04159_);
  not (_28153_, _28151_);
  nor (_28154_, _28153_, _28149_);
  nor (_28155_, _28154_, _28033_);
  nor (_28156_, _28155_, _03174_);
  and (_28157_, _11619_, _04650_);
  nor (_28158_, _28157_, _28034_);
  and (_28159_, _28158_, _03174_);
  nor (_28160_, _28159_, _28156_);
  or (_28161_, _28160_, _34702_);
  or (_28162_, _34698_, \oc8051_golden_model_1.SP [5]);
  and (_28164_, _28162_, _36029_);
  and (_35293_, _28164_, _28161_);
  nor (_28165_, _04650_, _10276_);
  and (_28166_, _11769_, _04650_);
  nor (_28167_, _28166_, _28165_);
  nor (_28168_, _28167_, _03131_);
  nor (_28169_, _04787_, _10307_);
  nor (_28170_, _28165_, _06241_);
  not (_28171_, _28170_);
  nor (_28172_, _28171_, _28169_);
  nor (_28174_, _11636_, _10307_);
  nor (_28175_, _28174_, _28165_);
  and (_28176_, _28175_, _02952_);
  and (_28177_, _04650_, \oc8051_golden_model_1.ACC [6]);
  nor (_28178_, _28177_, _28165_);
  or (_28179_, _28178_, _03826_);
  nand (_28180_, _09213_, \oc8051_golden_model_1.SP [6]);
  nor (_28181_, _10244_, \oc8051_golden_model_1.SP [6]);
  nor (_28182_, _28181_, _10245_);
  not (_28183_, _28182_);
  nor (_28185_, _28183_, _02558_);
  nor (_28186_, _28185_, _02952_);
  and (_28187_, _28186_, _28180_);
  and (_28188_, _28187_, _28179_);
  nor (_28189_, _28188_, _05382_);
  not (_28190_, _28189_);
  nor (_28191_, _28190_, _28176_);
  nor (_28192_, _28183_, _02556_);
  or (_28193_, _28192_, _02947_);
  nor (_28194_, _28193_, _28191_);
  nor (_28196_, _28065_, _10276_);
  nor (_28197_, _28196_, _10282_);
  and (_28198_, _28197_, _02947_);
  nor (_28199_, _28198_, _28194_);
  and (_28200_, _28199_, _02959_);
  nor (_28201_, _28178_, _02959_);
  or (_28202_, _28201_, _28200_);
  and (_28203_, _28202_, _03947_);
  nor (_28204_, _28074_, \oc8051_golden_model_1.SP [6]);
  nor (_28205_, _28204_, _10293_);
  and (_28207_, _28205_, _02886_);
  nor (_28208_, _28207_, _28203_);
  nor (_28209_, _28208_, _10292_);
  nor (_28210_, _28183_, _04126_);
  nor (_28211_, _28210_, _06793_);
  not (_28212_, _28211_);
  nor (_28213_, _28212_, _28209_);
  nor (_28214_, _28213_, _28172_);
  nor (_28215_, _28214_, _02855_);
  and (_28216_, _05847_, _04650_);
  nor (_28218_, _28216_, _28165_);
  and (_28219_, _28218_, _02855_);
  nor (_28220_, _28219_, _28215_);
  and (_28221_, _28220_, _02851_);
  nor (_28222_, _11751_, _10307_);
  nor (_28223_, _28222_, _28165_);
  nor (_28224_, _28223_, _02851_);
  or (_28225_, _28224_, _28221_);
  and (_28226_, _28225_, _03884_);
  and (_28227_, _11758_, _04650_);
  nor (_28229_, _28227_, _28165_);
  nor (_28230_, _28229_, _03884_);
  or (_28231_, _28230_, _02517_);
  or (_28232_, _28231_, _28226_);
  nand (_28233_, _28183_, _02517_);
  and (_28234_, _28233_, _28232_);
  and (_28235_, _28234_, _05279_);
  and (_28236_, _11646_, _04650_);
  nor (_28237_, _28236_, _28165_);
  nor (_28238_, _28237_, _05279_);
  or (_28240_, _28238_, _28235_);
  and (_28241_, _28240_, _03131_);
  nor (_28242_, _28241_, _28168_);
  nor (_28243_, _28242_, _03020_);
  nor (_28244_, _28165_, _04838_);
  not (_28245_, _28244_);
  nor (_28246_, _28229_, _05274_);
  and (_28247_, _28246_, _28245_);
  nor (_28248_, _28247_, _28243_);
  nor (_28249_, _28248_, _10251_);
  nor (_28251_, _28178_, _03140_);
  and (_28252_, _28251_, _28245_);
  and (_28253_, _28182_, _02533_);
  nor (_28254_, _28253_, _28252_);
  and (_28255_, _28254_, _05781_);
  not (_28256_, _28255_);
  nor (_28257_, _28256_, _28249_);
  nor (_28258_, _11644_, _10307_);
  nor (_28259_, _28258_, _28165_);
  and (_28260_, _28259_, _03036_);
  nor (_28262_, _28260_, _28257_);
  and (_28263_, _28262_, _05786_);
  nor (_28264_, _11768_, _10307_);
  nor (_28265_, _28264_, _28165_);
  nor (_28266_, _28265_, _05786_);
  or (_28267_, _28266_, _28263_);
  and (_28268_, _28267_, _10250_);
  nor (_28269_, _10280_, _10276_);
  nor (_28270_, _28269_, _10281_);
  not (_28271_, _28270_);
  and (_28273_, _28271_, _03148_);
  or (_28274_, _28273_, _02531_);
  nor (_28275_, _28274_, _28268_);
  and (_28276_, _28183_, _02531_);
  or (_28277_, _28276_, _02897_);
  nor (_28278_, _28277_, _28275_);
  and (_28279_, _28271_, _02897_);
  or (_28280_, _28279_, _03166_);
  nor (_28281_, _28280_, _28278_);
  and (_28282_, _28175_, _03166_);
  nor (_28284_, _28282_, _04159_);
  not (_28285_, _28284_);
  nor (_28286_, _28285_, _28281_);
  nor (_28287_, _28183_, _03916_);
  nor (_28288_, _28287_, _03174_);
  not (_28289_, _28288_);
  nor (_28290_, _28289_, _28286_);
  and (_28291_, _11821_, _04650_);
  or (_28292_, _28165_, _03178_);
  nor (_28293_, _28292_, _28291_);
  nor (_28295_, _28293_, _28290_);
  or (_28296_, _28295_, _34702_);
  or (_28297_, _34698_, \oc8051_golden_model_1.SP [6]);
  and (_28298_, _28297_, _36029_);
  and (_35294_, _28298_, _28296_);
  and (_35295_, \oc8051_golden_model_1.TCON [0], _36029_);
  and (_35296_, \oc8051_golden_model_1.TCON [1], _36029_);
  and (_35297_, \oc8051_golden_model_1.TCON [2], _36029_);
  and (_35298_, \oc8051_golden_model_1.TCON [3], _36029_);
  and (_35299_, \oc8051_golden_model_1.TCON [4], _36029_);
  and (_35301_, \oc8051_golden_model_1.TCON [5], _36029_);
  and (_35302_, \oc8051_golden_model_1.TCON [6], _36029_);
  and (_35303_, \oc8051_golden_model_1.TH0 [0], _36029_);
  and (_35304_, \oc8051_golden_model_1.TH0 [1], _36029_);
  and (_35305_, \oc8051_golden_model_1.TH0 [2], _36029_);
  and (_35306_, \oc8051_golden_model_1.TH0 [3], _36029_);
  and (_35307_, \oc8051_golden_model_1.TH0 [4], _36029_);
  and (_35308_, \oc8051_golden_model_1.TH0 [5], _36029_);
  and (_35309_, \oc8051_golden_model_1.TH0 [6], _36029_);
  and (_35310_, \oc8051_golden_model_1.TH1 [0], _36029_);
  and (_35312_, \oc8051_golden_model_1.TH1 [1], _36029_);
  and (_35313_, \oc8051_golden_model_1.TH1 [2], _36029_);
  and (_35314_, \oc8051_golden_model_1.TH1 [3], _36029_);
  and (_35315_, \oc8051_golden_model_1.TH1 [4], _36029_);
  and (_35316_, \oc8051_golden_model_1.TH1 [5], _36029_);
  and (_35317_, \oc8051_golden_model_1.TH1 [6], _36029_);
  and (_35318_, \oc8051_golden_model_1.TL0 [0], _36029_);
  and (_35319_, \oc8051_golden_model_1.TL0 [1], _36029_);
  and (_35320_, \oc8051_golden_model_1.TL0 [2], _36029_);
  and (_35321_, \oc8051_golden_model_1.TL0 [3], _36029_);
  and (_35323_, \oc8051_golden_model_1.TL0 [4], _36029_);
  and (_35324_, \oc8051_golden_model_1.TL0 [5], _36029_);
  and (_35325_, \oc8051_golden_model_1.TL0 [6], _36029_);
  and (_35326_, \oc8051_golden_model_1.TL1 [0], _36029_);
  and (_35327_, \oc8051_golden_model_1.TL1 [1], _36029_);
  and (_35328_, \oc8051_golden_model_1.TL1 [2], _36029_);
  and (_35329_, \oc8051_golden_model_1.TL1 [3], _36029_);
  and (_35330_, \oc8051_golden_model_1.TL1 [4], _36029_);
  and (_35331_, \oc8051_golden_model_1.TL1 [5], _36029_);
  and (_35332_, \oc8051_golden_model_1.TL1 [6], _36029_);
  and (_35334_, \oc8051_golden_model_1.TMOD [0], _36029_);
  and (_35335_, \oc8051_golden_model_1.TMOD [1], _36029_);
  and (_35336_, \oc8051_golden_model_1.TMOD [2], _36029_);
  and (_35337_, \oc8051_golden_model_1.TMOD [3], _36029_);
  and (_35338_, \oc8051_golden_model_1.TMOD [4], _36029_);
  and (_35339_, \oc8051_golden_model_1.TMOD [5], _36029_);
  and (_35340_, \oc8051_golden_model_1.TMOD [6], _36029_);
  and (_28303_, _34702_, \oc8051_golden_model_1.P0INREG [0]);
  or (_28304_, _28303_, _00760_);
  and (_35342_, _28304_, _36029_);
  and (_28306_, _34702_, \oc8051_golden_model_1.P0INREG [1]);
  or (_28307_, _28306_, _00753_);
  and (_35343_, _28307_, _36029_);
  and (_28308_, _34702_, \oc8051_golden_model_1.P0INREG [2]);
  or (_28309_, _28308_, _00738_);
  and (_35344_, _28309_, _36029_);
  and (_28310_, _34702_, \oc8051_golden_model_1.P0INREG [3]);
  or (_28311_, _28310_, _00746_);
  and (_35345_, _28311_, _36029_);
  and (_28312_, _34702_, \oc8051_golden_model_1.P0INREG [4]);
  or (_28314_, _28312_, _00725_);
  and (_35346_, _28314_, _36029_);
  and (_28315_, _34702_, \oc8051_golden_model_1.P0INREG [5]);
  or (_28316_, _28315_, _00718_);
  and (_35347_, _28316_, _36029_);
  and (_28317_, _34702_, \oc8051_golden_model_1.P0INREG [6]);
  or (_28318_, _28317_, _00703_);
  and (_35349_, _28318_, _36029_);
  and (_28319_, _34702_, \oc8051_golden_model_1.P1INREG [0]);
  or (_28320_, _28319_, _00513_);
  and (_35350_, _28320_, _36029_);
  and (_28321_, _34702_, \oc8051_golden_model_1.P1INREG [1]);
  or (_28322_, _28321_, _00486_);
  and (_35351_, _28322_, _36029_);
  and (_28323_, _34702_, \oc8051_golden_model_1.P1INREG [2]);
  or (_28324_, _28323_, _00504_);
  and (_35353_, _28324_, _36029_);
  and (_28325_, _34702_, \oc8051_golden_model_1.P1INREG [3]);
  or (_28326_, _28325_, _00494_);
  and (_35354_, _28326_, _36029_);
  and (_28329_, _34702_, \oc8051_golden_model_1.P1INREG [4]);
  or (_28330_, _28329_, _00474_);
  and (_35355_, _28330_, _36029_);
  and (_28331_, _34702_, \oc8051_golden_model_1.P1INREG [5]);
  or (_28332_, _28331_, _00443_);
  and (_35356_, _28332_, _36029_);
  and (_28333_, _34702_, \oc8051_golden_model_1.P1INREG [6]);
  or (_28334_, _28333_, _00464_);
  and (_35357_, _28334_, _36029_);
  and (_28335_, _34702_, \oc8051_golden_model_1.P2INREG [0]);
  or (_28337_, _28335_, _00536_);
  and (_35359_, _28337_, _36029_);
  and (_28338_, _34702_, \oc8051_golden_model_1.P2INREG [1]);
  or (_28339_, _28338_, _00544_);
  and (_35360_, _28339_, _36029_);
  and (_28340_, _34702_, \oc8051_golden_model_1.P2INREG [2]);
  or (_28341_, _28340_, _00529_);
  and (_35361_, _28341_, _36029_);
  and (_28342_, _34702_, \oc8051_golden_model_1.P2INREG [3]);
  or (_28343_, _28342_, _00553_);
  and (_35362_, _28343_, _36029_);
  and (_28345_, _34702_, \oc8051_golden_model_1.P2INREG [4]);
  or (_28346_, _28345_, _00576_);
  and (_35363_, _28346_, _36029_);
  and (_28347_, _34702_, \oc8051_golden_model_1.P2INREG [5]);
  or (_28348_, _28347_, _00585_);
  and (_35364_, _28348_, _36029_);
  and (_28349_, _34702_, \oc8051_golden_model_1.P2INREG [6]);
  or (_28350_, _28349_, _00566_);
  and (_35365_, _28350_, _36029_);
  and (_28352_, _34702_, \oc8051_golden_model_1.P3INREG [0]);
  or (_28353_, _28352_, _00611_);
  and (_35367_, _28353_, _36029_);
  and (_28354_, _34702_, \oc8051_golden_model_1.P3INREG [1]);
  or (_28355_, _28354_, _00631_);
  and (_35368_, _28355_, _36029_);
  and (_28356_, _34702_, \oc8051_golden_model_1.P3INREG [2]);
  or (_28357_, _28356_, _00621_);
  and (_35369_, _28357_, _36029_);
  and (_28358_, _34702_, \oc8051_golden_model_1.P3INREG [3]);
  or (_28360_, _28358_, _00639_);
  and (_35370_, _28360_, _36029_);
  and (_28361_, _34702_, \oc8051_golden_model_1.P3INREG [4]);
  or (_28362_, _28361_, _00649_);
  and (_35372_, _28362_, _36029_);
  and (_28363_, _34702_, \oc8051_golden_model_1.P3INREG [5]);
  or (_28364_, _28363_, _00664_);
  and (_35373_, _28364_, _36029_);
  and (_28365_, _34702_, \oc8051_golden_model_1.P3INREG [6]);
  or (_28366_, _28365_, _00656_);
  and (_35374_, _28366_, _36029_);
  and (_00005_[6], _00657_, _36029_);
  and (_00005_[5], _00665_, _36029_);
  and (_00005_[4], _00650_, _36029_);
  and (_00005_[3], _00640_, _36029_);
  and (_00005_[2], _00622_, _36029_);
  and (_00005_[1], _00633_, _36029_);
  and (_00005_[0], _00613_, _36029_);
  and (_00004_[6], _00568_, _36029_);
  and (_00004_[5], _00586_, _36029_);
  and (_00004_[4], _00577_, _36029_);
  and (_00004_[3], _00554_, _36029_);
  and (_00004_[2], _00530_, _36029_);
  and (_00004_[1], _00545_, _36029_);
  and (_00004_[0], _00537_, _36029_);
  and (_00003_[6], _00466_, _36029_);
  and (_00003_[5], _00444_, _36029_);
  and (_00003_[4], _00475_, _36029_);
  and (_00003_[3], _00496_, _36029_);
  and (_00003_[2], _00505_, _36029_);
  and (_00003_[1], _00487_, _36029_);
  and (_00003_[0], _00515_, _36029_);
  and (_00002_[6], _00704_, _36029_);
  and (_00002_[5], _00719_, _36029_);
  and (_00002_[4], _00726_, _36029_);
  and (_00002_[3], _00747_, _36029_);
  and (_00002_[2], _00739_, _36029_);
  and (_00002_[1], _00754_, _36029_);
  and (_00002_[0], _00761_, _36029_);
  or (_28370_, _09384_, _02304_);
  and (_28372_, _28370_, op0_cnst);
  and (_28373_, _28372_, _34698_);
  and (_28374_, _28373_, _36029_);
  or (_28375_, _27524_, _32054_);
  nand (_28376_, _27524_, _32054_);
  and (_28377_, _28376_, _28375_);
  and (_28378_, _27645_, _32183_);
  nor (_28379_, _27645_, _32183_);
  or (_28380_, _28379_, _28378_);
  or (_28381_, _28380_, _28377_);
  and (_28383_, _27893_, _30514_);
  nor (_28384_, _27893_, _30514_);
  or (_28385_, _28384_, _28383_);
  and (_28386_, _27769_, _30508_);
  nor (_28387_, _27769_, _30508_);
  or (_28388_, _28387_, _28386_);
  or (_28389_, _28388_, _28385_);
  or (_28390_, _28389_, _28381_);
  nor (_28391_, _28160_, _30526_);
  and (_28392_, _28160_, _30526_);
  or (_28393_, _28392_, _28391_);
  and (_28394_, _28026_, _30520_);
  nor (_28395_, _28026_, _30520_);
  or (_28396_, _28395_, _28394_);
  or (_28397_, _28396_, _28393_);
  nor (_28398_, _10389_, _30488_);
  and (_28399_, _10389_, _30488_);
  or (_28400_, _28399_, _28398_);
  nor (_28401_, _28295_, _30532_);
  and (_28402_, _28295_, _30532_);
  or (_28404_, _28402_, _28401_);
  or (_28405_, _28404_, _28400_);
  or (_28406_, _28405_, _28397_);
  or (_28407_, _28406_, _28390_);
  and (_00007_, _28407_, _28374_);
  or (_28408_, _10239_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_28409_, _10239_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_28410_, _28409_, _28408_);
  nor (_28411_, _26906_, _31004_);
  and (_28412_, _26906_, _31004_);
  or (_28414_, _28412_, _28411_);
  and (_28415_, _27437_, _29741_);
  nor (_28416_, _27437_, _29741_);
  nor (_28417_, _27022_, _31040_);
  and (_28418_, _27022_, _31040_);
  or (_28419_, _28418_, _28417_);
  not (_28420_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_28421_, _27251_, _28420_);
  and (_28422_, _27251_, _28420_);
  or (_28423_, _28422_, _28421_);
  or (_28425_, _28423_, _28419_);
  and (_28426_, _27136_, _31054_);
  nor (_28427_, _26658_, _30996_);
  and (_28428_, _26658_, _30996_);
  or (_28429_, _28428_, _28427_);
  nor (_28430_, _27136_, _31054_);
  or (_28431_, _28430_, _28429_);
  or (_28432_, _28431_, _28426_);
  or (_28433_, _28432_, _28425_);
  or (_28434_, _28433_, _28416_);
  or (_28436_, _28434_, _28415_);
  or (_28437_, _28436_, _28414_);
  or (_28438_, _28437_, _28410_);
  and (_00006_, _28438_, _28374_);
  or (_00001_, _28372_, rst);
  and (_00005_[7], _00672_, _36029_);
  and (_00004_[7], _00593_, _36029_);
  and (_00003_[7], _00456_, _36029_);
  and (_00002_[7], _00712_, _36029_);
  not (_28439_, _34658_);
  nor (_28441_, _05630_, _28439_);
  and (_28442_, _05630_, _28439_);
  or (_28443_, _28442_, _28441_);
  not (_28444_, _34675_);
  nor (_28445_, _05661_, _28444_);
  and (_28446_, _05661_, _28444_);
  or (_28447_, _28446_, _28445_);
  or (_28448_, _28447_, _28443_);
  nand (_28449_, _05598_, _34692_);
  or (_28450_, _05598_, _34692_);
  and (_28451_, _28450_, _28449_);
  nor (_28452_, _05563_, _34573_);
  and (_28453_, _05563_, _34573_);
  or (_28454_, _28453_, _28452_);
  or (_28455_, _28454_, _28451_);
  or (_28456_, _28455_, _28448_);
  or (_28457_, _03120_, _34641_);
  nand (_28458_, _03120_, _34641_);
  and (_28459_, _28458_, _28457_);
  nand (_28460_, _03302_, _34624_);
  or (_28463_, _03302_, _34624_);
  and (_28464_, _28463_, _28460_);
  or (_28465_, _28464_, _28459_);
  nand (_28466_, _03492_, _34590_);
  or (_28467_, _03492_, _34590_);
  and (_28468_, _28467_, _28466_);
  or (_28469_, _03705_, _34607_);
  nand (_28470_, _03705_, _34607_);
  and (_28471_, _28470_, _28469_);
  or (_28472_, _28471_, _28468_);
  or (_28474_, _28472_, _28465_);
  or (_28475_, _28474_, _28456_);
  and (_28476_, _34939_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28477_, _28476_, _35492_);
  nor (_28478_, _28476_, _35492_);
  or (_28479_, _28478_, _28477_);
  or (_28480_, _28479_, _02711_);
  nand (_28481_, _03047_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_28482_, _02496_, _30104_);
  and (_28483_, _02496_, _30104_);
  or (_28485_, _28483_, _28482_);
  or (_28486_, _02465_, _30202_);
  nand (_28487_, _02465_, _30202_);
  and (_28488_, _28487_, _28486_);
  or (_28489_, _28488_, _28485_);
  or (_28490_, _02506_, _30032_);
  nand (_28491_, _02506_, _30032_);
  and (_28492_, _28491_, _28490_);
  or (_28493_, _02336_, _30170_);
  or (_28494_, _02505_, _35421_);
  and (_28496_, _28494_, _28493_);
  or (_28497_, _28496_, _28492_);
  or (_28498_, _28497_, _28489_);
  and (_28499_, _02432_, _30149_);
  nor (_28500_, _02432_, _30149_);
  or (_28501_, _28500_, _28499_);
  nor (_28502_, _02401_, _30126_);
  and (_28503_, _02401_, _30126_);
  or (_28504_, _28503_, _28502_);
  or (_28505_, _28504_, _28501_);
  and (_28507_, _02509_, _30056_);
  nor (_28508_, _02509_, _30056_);
  or (_28509_, _28508_, _28507_);
  not (_28510_, _02304_);
  nor (_28511_, _28510_, _30078_);
  and (_28512_, _28510_, _30078_);
  or (_28513_, _28512_, _28511_);
  or (_28514_, _28513_, _28509_);
  or (_28515_, _28514_, _28505_);
  or (_28516_, _28515_, _28498_);
  nor (_28518_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28519_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_28520_, _28519_, _28518_);
  nor (_28521_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_28522_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_28523_, _28522_, _28521_);
  and (_28524_, _28523_, _28520_);
  or (_28525_, \oc8051_golden_model_1.PC [12], _30567_);
  or (_28526_, _24108_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28527_, _28526_, _28525_);
  or (_28529_, \oc8051_golden_model_1.PC [13], _30542_);
  or (_28530_, _08887_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_28531_, _28530_, _28529_);
  and (_28532_, _28531_, _28527_);
  and (_28533_, _28532_, _28524_);
  and (_28534_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28535_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_28536_, _28535_, _28534_);
  nor (_28537_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_28538_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_28540_, _28538_, _28537_);
  and (_28541_, _28540_, _28536_);
  and (_28542_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28543_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_28544_, _28543_, _28542_);
  nor (_28545_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_28546_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_28547_, _28546_, _28545_);
  and (_28548_, _28547_, _28544_);
  and (_28549_, _28548_, _28541_);
  and (_28551_, _28549_, _28533_);
  or (_28552_, \oc8051_golden_model_1.PC [0], _35481_);
  or (_28553_, _02247_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28554_, _28553_, _28552_);
  or (_28555_, _02218_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_28556_, \oc8051_golden_model_1.PC [1], _35485_);
  and (_28557_, _28556_, _28555_);
  and (_28558_, _28557_, _28554_);
  and (_28559_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_28560_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_28562_, _28560_, _28559_);
  or (_28563_, \oc8051_golden_model_1.PC [3], _35492_);
  or (_28564_, _02214_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28565_, _28564_, _28563_);
  and (_28566_, _28565_, _28562_);
  and (_28567_, _28566_, _28558_);
  or (_28568_, \oc8051_golden_model_1.PC [4], _35496_);
  nand (_28569_, \oc8051_golden_model_1.PC [4], _35496_);
  and (_28570_, _28569_, _28568_);
  or (_28571_, _21725_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_28573_, \oc8051_golden_model_1.PC [5], _35500_);
  and (_28574_, _28573_, _28571_);
  and (_28575_, _28574_, _28570_);
  or (_28576_, \oc8051_golden_model_1.PC [6], _35504_);
  nand (_28577_, \oc8051_golden_model_1.PC [6], _35504_);
  and (_28578_, _28577_, _28576_);
  and (_28579_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_28580_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_28581_, _28580_, _28579_);
  and (_28582_, _28581_, _28578_);
  and (_28584_, _28582_, _28575_);
  and (_28585_, _28584_, _28567_);
  and (_28586_, _28585_, _28551_);
  and (_28587_, _28586_, _34698_);
  and (_28588_, _28587_, _28516_);
  and (_28589_, _28588_, _28481_);
  and (_28590_, _28589_, _28480_);
  nor (_28591_, _34945_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_28592_, _28591_, _34946_);
  nor (_28593_, _23124_, _03044_);
  and (_28595_, _23109_, _03044_);
  nor (_28596_, _28595_, _28593_);
  or (_28597_, _28596_, _28592_);
  nand (_28598_, _28596_, _28592_);
  and (_28599_, _28598_, _28597_);
  and (_28600_, _28599_, _28590_);
  nor (_28601_, _23823_, _03044_);
  and (_28602_, _23755_, _03044_);
  nor (_28603_, _28602_, _28601_);
  nand (_28604_, _28603_, _35902_);
  or (_28606_, _28603_, _35902_);
  and (_28607_, _28606_, _28604_);
  nand (_28608_, _03051_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_28609_, _03047_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_28610_, _03051_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_28611_, _28610_, _28609_);
  and (_28612_, _28611_, _28608_);
  and (_28613_, _28612_, _28607_);
  and (_28614_, _28613_, _28600_);
  and (_28615_, _28614_, _28475_);
  or (_28617_, _02832_, _32048_);
  nand (_28618_, _02832_, _32048_);
  and (_28619_, _28618_, _28617_);
  nor (_28620_, _03672_, _32164_);
  and (_28621_, _03672_, _32164_);
  or (_28622_, _28621_, _28620_);
  or (_28623_, _28622_, _28619_);
  or (_28624_, _03215_, _31930_);
  nand (_28625_, _03215_, _31930_);
  and (_28626_, _28625_, _28624_);
  nor (_28628_, _04662_, _32203_);
  and (_28629_, _04662_, _32203_);
  or (_28630_, _28629_, _28628_);
  or (_28631_, _28630_, _28626_);
  or (_28632_, _28631_, _28623_);
  or (_28633_, _03260_, _31870_);
  nand (_28634_, _03260_, _31870_);
  and (_28635_, _28634_, _28633_);
  or (_28636_, _02799_, _32073_);
  nand (_28637_, _02799_, _32073_);
  and (_28639_, _28637_, _28636_);
  or (_28640_, _28639_, _28635_);
  or (_28641_, _02932_, _32135_);
  nand (_28642_, _02932_, _32135_);
  and (_28643_, _28642_, _28641_);
  and (_28644_, _02768_, _31991_);
  nor (_28645_, _02768_, _31991_);
  or (_28646_, _28645_, _28644_);
  or (_28647_, _28646_, _28643_);
  or (_28648_, _28647_, _28640_);
  or (_28650_, _28648_, _28632_);
  and (_28651_, _22409_, \oc8051_golden_model_1.ACC [7]);
  nor (_28652_, _22409_, \oc8051_golden_model_1.ACC [7]);
  nor (_28653_, _28652_, _28651_);
  and (_28654_, _22055_, \oc8051_golden_model_1.ACC [6]);
  nor (_28655_, _22055_, \oc8051_golden_model_1.ACC [6]);
  nor (_28656_, _28655_, _28654_);
  and (_28657_, _21685_, \oc8051_golden_model_1.ACC [5]);
  nor (_28658_, _21685_, \oc8051_golden_model_1.ACC [5]);
  nor (_28659_, _28658_, _28657_);
  and (_28661_, _21325_, \oc8051_golden_model_1.ACC [4]);
  and (_28662_, _28661_, _28659_);
  nor (_28663_, _28662_, _28657_);
  nor (_28664_, _02703_, _02700_);
  nor (_28665_, _28664_, _02702_);
  not (_28666_, _28665_);
  nor (_28667_, _21325_, \oc8051_golden_model_1.ACC [4]);
  nor (_28668_, _28667_, _28661_);
  and (_28669_, _28668_, _28659_);
  nand (_28670_, _28669_, _28666_);
  nand (_28672_, _28670_, _28663_);
  and (_28673_, _28672_, _28656_);
  or (_28674_, _28673_, _28654_);
  and (_28675_, _28674_, _28653_);
  nor (_28676_, _28675_, _28651_);
  and (_28677_, _23109_, _22771_);
  and (_28678_, _23755_, _23446_);
  and (_28679_, _28678_, _28677_);
  not (_28680_, _28679_);
  nor (_28681_, _28680_, _28676_);
  and (_28684_, _24420_, _24089_);
  and (_28686_, _28684_, _28681_);
  and (_28688_, _28686_, _24747_);
  and (_28690_, _28688_, _09008_);
  nor (_28692_, _28688_, _09008_);
  nor (_28694_, _28692_, _28690_);
  nor (_28696_, _28694_, _02584_);
  and (_28698_, _09436_, _02585_);
  and (_28700_, _09008_, _02600_);
  and (_28702_, _09351_, _02571_);
  nor (_28705_, _28702_, _28700_);
  and (_28706_, _28705_, _02586_);
  or (_28707_, _28706_, _02580_);
  nor (_28708_, _28707_, _28698_);
  nor (_28709_, _06227_, _02579_);
  nor (_28710_, _28709_, _02548_);
  not (_28711_, _28710_);
  nor (_28712_, _28711_, _28708_);
  nor (_28713_, _28712_, _28696_);
  nor (_28714_, _28713_, _02583_);
  nor (_28716_, _09351_, _02543_);
  or (_28717_, _28716_, _28714_);
  and (_28718_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28719_, _28476_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28720_, _28719_, _34943_);
  and (_28721_, _28720_, _35924_);
  and (_28722_, _28721_, _28718_);
  and (_28723_, _28722_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28724_, _28723_, _30578_);
  and (_28725_, _28723_, _30578_);
  or (_28727_, _28725_, _28724_);
  and (_28728_, _28727_, _28717_);
  nor (_28729_, _28727_, _28717_);
  or (_28730_, _28729_, _28728_);
  and (_28731_, _28730_, _28650_);
  and (property_invalid_rom_pc, _28731_, _28615_);
  nor (_28732_, _30488_, \oc8051_golden_model_1.SP [7]);
  and (_28733_, _30488_, \oc8051_golden_model_1.SP [7]);
  or (_28734_, _28733_, _28732_);
  nor (_28735_, _30532_, \oc8051_golden_model_1.SP [6]);
  and (_28737_, _30532_, \oc8051_golden_model_1.SP [6]);
  or (_28738_, _28737_, _28735_);
  and (_28739_, _30526_, \oc8051_golden_model_1.SP [5]);
  nor (_28740_, _30526_, \oc8051_golden_model_1.SP [5]);
  or (_28741_, _28740_, _28739_);
  and (_28742_, _30514_, \oc8051_golden_model_1.SP [3]);
  nor (_28743_, _30514_, \oc8051_golden_model_1.SP [3]);
  or (_28744_, _28743_, _28742_);
  and (_28745_, _30502_, \oc8051_golden_model_1.SP [1]);
  or (_28746_, _30496_, _02877_);
  nand (_28748_, _30496_, _02877_);
  and (_28749_, _28748_, _28746_);
  nor (_28750_, _30502_, \oc8051_golden_model_1.SP [1]);
  or (_28751_, _28750_, _28749_);
  or (_28752_, _28751_, _28745_);
  nor (_28753_, _30508_, \oc8051_golden_model_1.SP [2]);
  and (_28754_, _30508_, \oc8051_golden_model_1.SP [2]);
  or (_28755_, _28754_, _28753_);
  or (_28756_, _28755_, _28752_);
  or (_28757_, _28756_, _28744_);
  and (_28759_, _30520_, \oc8051_golden_model_1.SP [4]);
  nor (_28760_, _30520_, \oc8051_golden_model_1.SP [4]);
  or (_28761_, _28760_, _28759_);
  or (_28762_, _28761_, _28757_);
  or (_28763_, _28762_, _28741_);
  or (_28764_, _28763_, _28738_);
  or (_28765_, _28764_, _28734_);
  and (_28766_, _28372_, inst_finished_r);
  and (_28767_, _28766_, property_invalid_sp_1_r);
  and (property_invalid_sp, _28767_, _28765_);
  nand (_28769_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_28770_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_28771_, _28770_, _28769_);
  and (_28772_, _26563_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_28773_, \oc8051_golden_model_1.PSW [1], _30996_);
  or (_28774_, _28773_, _28772_);
  or (_28775_, _28774_, _28771_);
  and (_28776_, _27026_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_28777_, \oc8051_golden_model_1.PSW [4], _31054_);
  or (_28778_, _28777_, _28776_);
  and (_28780_, _26911_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_28781_, \oc8051_golden_model_1.PSW [3], _31040_);
  or (_28782_, _28781_, _28780_);
  or (_28783_, _28782_, _28778_);
  or (_28784_, _28783_, _28775_);
  and (_28785_, _07319_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_28786_, \oc8051_golden_model_1.PSW [7], _30969_);
  or (_28787_, _28786_, _28785_);
  and (_28788_, _27141_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_28789_, \oc8051_golden_model_1.PSW [5], _28420_);
  or (_28791_, _28789_, _28788_);
  nand (_28792_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_28793_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_28794_, _28793_, _28792_);
  or (_28795_, _28794_, _28791_);
  or (_28796_, _28795_, _28787_);
  or (_28797_, _28796_, _28784_);
  and (_28798_, _28797_, property_invalid_psw_1_r);
  and (property_invalid_psw, _28798_, _28766_);
  nand (_28799_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_28801_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_28802_, _28801_, _28799_);
  and (_28803_, _19392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_28804_, \oc8051_golden_model_1.P3 [2], _31782_);
  or (_28805_, _28804_, _28803_);
  or (_28806_, _28805_, _28802_);
  and (_28807_, \oc8051_golden_model_1.P3 [0], _31756_);
  and (_28808_, _19173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_28809_, _28808_, _28807_);
  and (_28810_, _19278_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_28812_, \oc8051_golden_model_1.P3 [1], _31769_);
  or (_28813_, _28812_, _28810_);
  or (_28814_, _28813_, _28809_);
  or (_28815_, _28814_, _28806_);
  or (_28816_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_28817_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_28818_, _28817_, _28816_);
  or (_28819_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_28820_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_28821_, _28820_, _28819_);
  or (_28823_, _28821_, _28818_);
  and (_28824_, _08738_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_28825_, \oc8051_golden_model_1.P3 [7], _31451_);
  or (_28826_, _28825_, _28824_);
  nand (_28827_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_28828_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_28829_, _28828_, _28827_);
  or (_28830_, _28829_, _28826_);
  or (_28831_, _28830_, _28823_);
  or (_28832_, _28831_, _28815_);
  and (property_invalid_p3, _28832_, _28766_);
  nand (_28834_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_28835_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_28836_, _28835_, _28834_);
  and (_28837_, _18613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_28838_, \oc8051_golden_model_1.P2 [2], _31681_);
  or (_28839_, _28838_, _28837_);
  or (_28840_, _28839_, _28836_);
  and (_28841_, \oc8051_golden_model_1.P2 [0], _31648_);
  and (_28842_, _18394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_28844_, _28842_, _28841_);
  and (_28845_, _18500_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_28846_, \oc8051_golden_model_1.P2 [1], _31661_);
  or (_28847_, _28846_, _28845_);
  or (_28848_, _28847_, _28844_);
  or (_28849_, _28848_, _28840_);
  or (_28850_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_28851_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_28852_, _28851_, _28850_);
  or (_28853_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_28855_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_28856_, _28855_, _28853_);
  or (_28857_, _28856_, _28852_);
  and (_28858_, _08635_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_28859_, \oc8051_golden_model_1.P2 [7], _31435_);
  or (_28860_, _28859_, _28858_);
  nand (_28861_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_28862_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_28863_, _28862_, _28861_);
  or (_28864_, _28863_, _28860_);
  or (_28866_, _28864_, _28857_);
  or (_28867_, _28866_, _28849_);
  and (property_invalid_p2, _28867_, _28766_);
  nand (_28868_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_28869_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_28870_, _28869_, _28868_);
  and (_28871_, _17835_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_28872_, \oc8051_golden_model_1.P1 [2], _31582_);
  or (_28873_, _28872_, _28871_);
  or (_28874_, _28873_, _28870_);
  and (_28876_, \oc8051_golden_model_1.P1 [0], _31555_);
  and (_28877_, _17616_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_28878_, _28877_, _28876_);
  and (_28879_, _17721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_28880_, \oc8051_golden_model_1.P1 [1], _31568_);
  or (_28881_, _28880_, _28879_);
  or (_28882_, _28881_, _28878_);
  or (_28883_, _28882_, _28874_);
  or (_28884_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_28885_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_28887_, _28885_, _28884_);
  or (_28888_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_28889_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_28890_, _28889_, _28888_);
  or (_28891_, _28890_, _28887_);
  and (_28892_, _08532_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_28893_, \oc8051_golden_model_1.P1 [7], _31417_);
  or (_28894_, _28893_, _28892_);
  nand (_28895_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_28896_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_28898_, _28896_, _28895_);
  or (_28899_, _28898_, _28894_);
  or (_28900_, _28899_, _28891_);
  or (_28901_, _28900_, _28883_);
  and (property_invalid_p1, _28901_, _28766_);
  nand (_28902_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_28903_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_28904_, _28903_, _28902_);
  and (_28905_, _16987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_28906_, \oc8051_golden_model_1.P0 [2], _31481_);
  or (_28908_, _28906_, _28905_);
  or (_28909_, _28908_, _28904_);
  and (_28910_, \oc8051_golden_model_1.P0 [0], _31458_);
  and (_28911_, _16742_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_28912_, _28911_, _28910_);
  and (_28913_, _16861_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_28914_, \oc8051_golden_model_1.P0 [1], _31477_);
  or (_28915_, _28914_, _28913_);
  or (_28916_, _28915_, _28912_);
  or (_28917_, _28916_, _28909_);
  or (_28919_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_28920_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_28921_, _28920_, _28919_);
  or (_28922_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_28923_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_28924_, _28923_, _28922_);
  or (_28925_, _28924_, _28921_);
  and (_28926_, _08417_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_28927_, \oc8051_golden_model_1.P0 [7], _31403_);
  or (_28928_, _28927_, _28926_);
  nand (_28930_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_28931_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_28932_, _28931_, _28930_);
  or (_28933_, _28932_, _28928_);
  or (_28934_, _28933_, _28925_);
  or (_28935_, _28934_, _28917_);
  and (property_invalid_p0, _28935_, _28766_);
  or (_28936_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_28937_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_28938_, _28937_, _28936_);
  or (_28940_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nand (_28941_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_28942_, _28941_, _28940_);
  or (_28943_, _28942_, _28938_);
  and (_28944_, _03375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_28945_, \oc8051_golden_model_1.IRAM[0] [0], _32339_);
  or (_28946_, _28945_, _28944_);
  and (_28947_, \oc8051_golden_model_1.IRAM[0] [1], _32352_);
  and (_28948_, _03949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_28949_, _28948_, _28947_);
  or (_28951_, _28949_, _28946_);
  or (_28952_, _28951_, _28943_);
  or (_28953_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_28954_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_28955_, _28954_, _28953_);
  or (_28956_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_28957_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_28958_, _28957_, _28956_);
  or (_28959_, _28958_, _28955_);
  or (_28960_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_28962_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_28963_, _28962_, _28960_);
  or (_28964_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_28965_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_28966_, _28965_, _28964_);
  or (_28967_, _28966_, _28963_);
  or (_28968_, _28967_, _28959_);
  or (_28969_, _28968_, _28952_);
  or (_28970_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_28971_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_28973_, _28971_, _28970_);
  or (_28974_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_28975_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_28976_, _28975_, _28974_);
  or (_28977_, _28976_, _28973_);
  or (_28978_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_28979_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_28980_, _28979_, _28978_);
  or (_28981_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand (_28982_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_28984_, _28982_, _28981_);
  or (_28985_, _28984_, _28980_);
  or (_28986_, _28985_, _28977_);
  and (_28987_, _05148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_28988_, \oc8051_golden_model_1.IRAM[1] [4], _32423_);
  or (_28989_, _28988_, _28987_);
  and (_28990_, \oc8051_golden_model_1.IRAM[1] [5], _32427_);
  and (_28991_, _04841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_28992_, _28991_, _28990_);
  or (_28993_, _28992_, _28989_);
  or (_28994_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_28995_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_28996_, _28995_, _28994_);
  or (_28997_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand (_28998_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_28999_, _28998_, _28997_);
  or (_29000_, _28999_, _28996_);
  or (_29001_, _29000_, _28993_);
  or (_29002_, _29001_, _28986_);
  or (_29003_, _29002_, _28969_);
  or (_29006_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_29007_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_29008_, _29007_, _29006_);
  or (_29009_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_29010_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_29011_, _29010_, _29009_);
  or (_29012_, _29011_, _29008_);
  and (_29013_, \oc8051_golden_model_1.IRAM[2] [2], _32442_);
  and (_29014_, _04384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_29015_, _29014_, _29013_);
  nand (_29017_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_29018_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_29019_, _29018_, _29017_);
  or (_29020_, _29019_, _29015_);
  or (_29021_, _29020_, _29012_);
  and (_29022_, _05154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_29023_, \oc8051_golden_model_1.IRAM[2] [4], _32447_);
  or (_29024_, _29023_, _29022_);
  and (_29025_, \oc8051_golden_model_1.IRAM[2] [5], _32450_);
  and (_29026_, _04847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_29028_, _29026_, _29025_);
  or (_29029_, _29028_, _29024_);
  or (_29030_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand (_29031_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_29032_, _29031_, _29030_);
  and (_29033_, _04573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_29034_, \oc8051_golden_model_1.IRAM[2] [7], _32455_);
  or (_29035_, _29034_, _29033_);
  or (_29036_, _29035_, _29032_);
  or (_29037_, _29036_, _29029_);
  or (_29039_, _29037_, _29021_);
  and (_29040_, \oc8051_golden_model_1.IRAM[3] [1], _32462_);
  and (_29041_, _03955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_29042_, _29041_, _29040_);
  and (_29043_, _03764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_29044_, \oc8051_golden_model_1.IRAM[3] [0], _32459_);
  or (_29045_, _29044_, _29043_);
  or (_29046_, _29045_, _29042_);
  and (_29047_, \oc8051_golden_model_1.IRAM[3] [2], _32465_);
  and (_29048_, _04381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_29050_, _29048_, _29047_);
  nand (_29051_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_29052_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_29053_, _29052_, _29051_);
  or (_29054_, _29053_, _29050_);
  or (_29055_, _29054_, _29046_);
  or (_29056_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand (_29057_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_29058_, _29057_, _29056_);
  and (_29059_, _04571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_29061_, \oc8051_golden_model_1.IRAM[3] [7], _32254_);
  or (_29062_, _29061_, _29059_);
  or (_29063_, _29062_, _29058_);
  or (_29064_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_29065_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_29066_, _29065_, _29064_);
  or (_29067_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_29068_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_29069_, _29068_, _29067_);
  or (_29070_, _29069_, _29066_);
  or (_29072_, _29070_, _29063_);
  or (_29073_, _29072_, _29055_);
  or (_29074_, _29073_, _29039_);
  or (_29075_, _29074_, _29003_);
  and (_29076_, _03780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_29077_, \oc8051_golden_model_1.IRAM[4] [0], _32482_);
  or (_29078_, _29077_, _29076_);
  and (_29079_, _03969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_29080_, \oc8051_golden_model_1.IRAM[4] [1], _32502_);
  or (_29081_, _29080_, _29079_);
  or (_29083_, _29081_, _29078_);
  or (_29084_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_29085_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_29086_, _29085_, _29084_);
  nand (_29087_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_29088_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_29089_, _29088_, _29087_);
  or (_29090_, _29089_, _29086_);
  or (_29091_, _29090_, _29083_);
  or (_29092_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_29094_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_29095_, _29094_, _29092_);
  or (_29096_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_29097_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_29098_, _29097_, _29096_);
  or (_29099_, _29098_, _29095_);
  or (_29100_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_29101_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_29102_, _29101_, _29100_);
  nand (_29103_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_29105_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_29106_, _29105_, _29103_);
  or (_29107_, _29106_, _29102_);
  or (_29108_, _29107_, _29099_);
  or (_29109_, _29108_, _29091_);
  or (_29110_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_29111_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_29112_, _29111_, _29110_);
  nand (_29113_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_29114_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_29115_, _29114_, _29113_);
  or (_29116_, _29115_, _29112_);
  or (_29117_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_29118_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_29119_, _29118_, _29117_);
  or (_29120_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_29121_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_29122_, _29121_, _29120_);
  or (_29123_, _29122_, _29119_);
  or (_29124_, _29123_, _29116_);
  or (_29126_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_29127_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_29128_, _29127_, _29126_);
  nand (_29129_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_29130_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_29131_, _29130_, _29129_);
  or (_29132_, _29131_, _29128_);
  and (_29133_, _05168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_29134_, \oc8051_golden_model_1.IRAM[5] [4], _32539_);
  or (_29135_, _29134_, _29133_);
  and (_29137_, \oc8051_golden_model_1.IRAM[5] [5], _32550_);
  and (_29138_, _04862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_29139_, _29138_, _29137_);
  or (_29140_, _29139_, _29135_);
  or (_29141_, _29140_, _29132_);
  or (_29142_, _29141_, _29124_);
  or (_29143_, _29142_, _29109_);
  nand (_29144_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_29145_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_29146_, _29145_, _29144_);
  and (_29148_, \oc8051_golden_model_1.IRAM[6] [2], _32596_);
  and (_29149_, _04396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_29150_, _29149_, _29148_);
  or (_29151_, _29150_, _29146_);
  or (_29152_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_29153_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_29154_, _29153_, _29152_);
  or (_29155_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_29156_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_29157_, _29156_, _29155_);
  or (_29159_, _29157_, _29154_);
  or (_29160_, _29159_, _29151_);
  and (_29161_, _04581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_29162_, \oc8051_golden_model_1.IRAM[6] [7], _32641_);
  or (_29163_, _29162_, _29161_);
  nand (_29164_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_29165_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_29166_, _29165_, _29164_);
  or (_29167_, _29166_, _29163_);
  and (_29168_, _05162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_29170_, \oc8051_golden_model_1.IRAM[6] [4], _32617_);
  or (_29171_, _29170_, _29168_);
  and (_29172_, \oc8051_golden_model_1.IRAM[6] [5], _32628_);
  and (_29173_, _04856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_29174_, _29173_, _29172_);
  or (_29175_, _29174_, _29171_);
  or (_29176_, _29175_, _29167_);
  or (_29177_, _29176_, _29160_);
  and (_29178_, _03963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_29179_, \oc8051_golden_model_1.IRAM[7] [1], _32667_);
  or (_29181_, _29179_, _29178_);
  and (_29182_, _03774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_29183_, \oc8051_golden_model_1.IRAM[7] [0], _32657_);
  or (_29184_, _29183_, _29182_);
  or (_29185_, _29184_, _29181_);
  nand (_29186_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_29187_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_29188_, _29187_, _29186_);
  and (_29189_, _04393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_29190_, \oc8051_golden_model_1.IRAM[7] [2], _32677_);
  or (_29192_, _29190_, _29189_);
  or (_29193_, _29192_, _29188_);
  or (_29194_, _29193_, _29185_);
  or (_29195_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_29196_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_29197_, _29196_, _29195_);
  or (_29198_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_29199_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_29200_, _29199_, _29198_);
  or (_29201_, _29200_, _29197_);
  and (_29203_, \oc8051_golden_model_1.IRAM[7] [7], _32266_);
  and (_29204_, _04579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_29205_, _29204_, _29203_);
  nand (_29206_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_29207_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_29208_, _29207_, _29206_);
  or (_29209_, _29208_, _29205_);
  or (_29210_, _29209_, _29201_);
  or (_29211_, _29210_, _29194_);
  or (_29212_, _29211_, _29177_);
  or (_29214_, _29212_, _29143_);
  or (_29215_, _29214_, _29075_);
  and (_29216_, _03796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_29217_, \oc8051_golden_model_1.IRAM[8] [0], _32723_);
  or (_29218_, _29217_, _29216_);
  and (_29219_, _03984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_29220_, \oc8051_golden_model_1.IRAM[8] [1], _32726_);
  or (_29221_, _29220_, _29219_);
  or (_29222_, _29221_, _29218_);
  or (_29223_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_29225_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_29226_, _29225_, _29223_);
  nand (_29227_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_29228_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_29229_, _29228_, _29227_);
  or (_29230_, _29229_, _29226_);
  or (_29231_, _29230_, _29222_);
  or (_29232_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_29233_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_29234_, _29233_, _29232_);
  or (_29236_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand (_29237_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_29238_, _29237_, _29236_);
  or (_29239_, _29238_, _29234_);
  or (_29240_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_29241_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_29242_, _29241_, _29240_);
  nand (_29243_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_29244_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_29245_, _29244_, _29243_);
  or (_29247_, _29245_, _29242_);
  or (_29248_, _29247_, _29239_);
  or (_29249_, _29248_, _29231_);
  or (_29250_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_29251_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_29252_, _29251_, _29250_);
  nand (_29253_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_29254_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_29255_, _29254_, _29253_);
  or (_29256_, _29255_, _29252_);
  or (_29258_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_29259_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_29260_, _29259_, _29258_);
  or (_29261_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_29262_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_29263_, _29262_, _29261_);
  or (_29264_, _29263_, _29260_);
  or (_29265_, _29264_, _29256_);
  or (_29266_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_29267_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_29269_, _29267_, _29266_);
  nand (_29270_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_29271_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_29272_, _29271_, _29270_);
  or (_29273_, _29272_, _29269_);
  and (_29274_, _05182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_29275_, \oc8051_golden_model_1.IRAM[9] [4], _32753_);
  or (_29276_, _29275_, _29274_);
  and (_29277_, _04876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_29278_, \oc8051_golden_model_1.IRAM[9] [5], _32756_);
  or (_29280_, _29278_, _29277_);
  or (_29281_, _29280_, _29276_);
  or (_29282_, _29281_, _29273_);
  or (_29283_, _29282_, _29265_);
  or (_29284_, _29283_, _29249_);
  or (_29285_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nand (_29286_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_29287_, _29286_, _29285_);
  and (_29288_, \oc8051_golden_model_1.IRAM[10] [2], _32770_);
  and (_29289_, _04415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_29291_, _29289_, _29288_);
  or (_29292_, _29291_, _29287_);
  or (_29293_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand (_29294_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_29295_, _29294_, _29293_);
  or (_29296_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand (_29297_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_29298_, _29297_, _29296_);
  or (_29299_, _29298_, _29295_);
  or (_29300_, _29299_, _29292_);
  and (_29302_, _04595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_29303_, \oc8051_golden_model_1.IRAM[10] [7], _32280_);
  or (_29304_, _29303_, _29302_);
  nand (_29305_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_29306_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_29307_, _29306_, _29305_);
  or (_29308_, _29307_, _29304_);
  and (_29309_, _05177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_29310_, \oc8051_golden_model_1.IRAM[10] [4], _32775_);
  or (_29311_, _29310_, _29309_);
  and (_29313_, _04871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_29314_, \oc8051_golden_model_1.IRAM[10] [5], _32778_);
  or (_29315_, _29314_, _29313_);
  or (_29316_, _29315_, _29311_);
  or (_29317_, _29316_, _29308_);
  or (_29318_, _29317_, _29300_);
  and (_29319_, _03791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_29320_, \oc8051_golden_model_1.IRAM[11] [0], _32787_);
  or (_29321_, _29320_, _29319_);
  and (_29322_, \oc8051_golden_model_1.IRAM[11] [1], _32790_);
  and (_29324_, _03979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_29325_, _29324_, _29322_);
  or (_29326_, _29325_, _29321_);
  nand (_29327_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_29328_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_29329_, _29328_, _29327_);
  and (_29330_, _04413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_29331_, \oc8051_golden_model_1.IRAM[11] [2], _32793_);
  or (_29332_, _29331_, _29330_);
  or (_29333_, _29332_, _29329_);
  or (_29335_, _29333_, _29326_);
  or (_29336_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_29337_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_29338_, _29337_, _29336_);
  or (_29339_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_29340_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_29341_, _29340_, _29339_);
  or (_29342_, _29341_, _29338_);
  and (_29343_, _04593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_29344_, \oc8051_golden_model_1.IRAM[11] [7], _32805_);
  or (_29346_, _29344_, _29343_);
  nand (_29347_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_29348_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_29349_, _29348_, _29347_);
  or (_29350_, _29349_, _29346_);
  or (_29351_, _29350_, _29342_);
  or (_29352_, _29351_, _29335_);
  or (_29353_, _29352_, _29318_);
  or (_29354_, _29353_, _29284_);
  or (_29355_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_29357_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_29358_, _29357_, _29355_);
  nand (_29359_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_29360_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_29361_, _29360_, _29359_);
  or (_29362_, _29361_, _29358_);
  and (_29363_, _03808_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_29364_, \oc8051_golden_model_1.IRAM[12] [0], _32809_);
  or (_29365_, _29364_, _29363_);
  and (_29366_, \oc8051_golden_model_1.IRAM[12] [1], _32812_);
  and (_29368_, _03996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_29369_, _29368_, _29366_);
  or (_29370_, _29369_, _29365_);
  or (_29371_, _29370_, _29362_);
  or (_29372_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_29373_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_29374_, _29373_, _29372_);
  nand (_29375_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_29376_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_29377_, _29376_, _29375_);
  or (_29379_, _29377_, _29374_);
  or (_29380_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_29381_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_29382_, _29381_, _29380_);
  or (_29383_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand (_29384_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_29385_, _29384_, _29383_);
  or (_29386_, _29385_, _29382_);
  or (_29387_, _29386_, _29379_);
  or (_29388_, _29387_, _29371_);
  or (_29390_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_29391_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_29392_, _29391_, _29390_);
  or (_29393_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_29394_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_29395_, _29394_, _29393_);
  or (_29396_, _29395_, _29392_);
  or (_29397_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_29398_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_29399_, _29398_, _29397_);
  nand (_29401_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_29402_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_29403_, _29402_, _29401_);
  or (_29404_, _29403_, _29399_);
  or (_29405_, _29404_, _29396_);
  and (_29406_, _05194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_29407_, \oc8051_golden_model_1.IRAM[13] [4], _32838_);
  or (_29408_, _29407_, _29406_);
  and (_29409_, _04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_29410_, \oc8051_golden_model_1.IRAM[13] [5], _32841_);
  or (_29412_, _29410_, _29409_);
  or (_29413_, _29412_, _29408_);
  or (_29414_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_29415_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_29416_, _29415_, _29414_);
  nand (_29417_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_29418_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_29419_, _29418_, _29417_);
  or (_29420_, _29419_, _29416_);
  or (_29421_, _29420_, _29413_);
  or (_29423_, _29421_, _29405_);
  or (_29424_, _29423_, _29388_);
  or (_29425_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand (_29426_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_29427_, _29426_, _29425_);
  or (_29428_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand (_29429_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_29430_, _29429_, _29428_);
  or (_29431_, _29430_, _29427_);
  and (_29432_, \oc8051_golden_model_1.IRAM[14] [2], _32855_);
  and (_29434_, _04427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_29435_, _29434_, _29432_);
  nand (_29436_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_29437_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_29438_, _29437_, _29436_);
  or (_29439_, _29438_, _29435_);
  or (_29440_, _29439_, _29431_);
  and (_29441_, \oc8051_golden_model_1.IRAM[14] [5], _32864_);
  and (_29442_, _04883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_29443_, _29442_, _29441_);
  and (_29445_, _05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_29446_, \oc8051_golden_model_1.IRAM[14] [4], _32861_);
  or (_29447_, _29446_, _29445_);
  or (_29448_, _29447_, _29443_);
  and (_29449_, \oc8051_golden_model_1.IRAM[14] [7], _32291_);
  and (_29450_, _04609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_29451_, _29450_, _29449_);
  nand (_29452_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_29453_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_29454_, _29453_, _29452_);
  or (_29456_, _29454_, _29451_);
  or (_29457_, _29456_, _29448_);
  or (_29458_, _29457_, _29440_);
  and (_29459_, _03991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_29460_, \oc8051_golden_model_1.IRAM[15] [1], _32875_);
  or (_29461_, _29460_, _29459_);
  and (_29462_, _03803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_29463_, \oc8051_golden_model_1.IRAM[15] [0], _32872_);
  or (_29464_, _29463_, _29462_);
  or (_29465_, _29464_, _29461_);
  or (_29467_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_29468_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_29469_, _29468_, _29467_);
  and (_29470_, _04425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_29471_, \oc8051_golden_model_1.IRAM[15] [2], _32878_);
  or (_29472_, _29471_, _29470_);
  or (_29473_, _29472_, _29469_);
  or (_29474_, _29473_, _29465_);
  nand (_29475_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_29476_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_29478_, _29476_, _29475_);
  and (_29479_, _04607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_29480_, \oc8051_golden_model_1.IRAM[15] [7], _32322_);
  or (_29481_, _29480_, _29479_);
  or (_29482_, _29481_, _29478_);
  or (_29483_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_29484_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_29485_, _29484_, _29483_);
  or (_29486_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_29487_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_29489_, _29487_, _29486_);
  or (_29490_, _29489_, _29485_);
  or (_29491_, _29490_, _29482_);
  or (_29492_, _29491_, _29474_);
  or (_29493_, _29492_, _29458_);
  or (_29494_, _29493_, _29424_);
  or (_29495_, _29494_, _29354_);
  or (_29496_, _29495_, _29215_);
  and (property_invalid_iram, _29496_, _28766_);
  nand (_29497_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_29499_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_29500_, _29499_, _29497_);
  and (_29501_, _16266_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_29502_, _16266_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_29503_, _29502_, _29501_);
  or (_29504_, _29503_, _29500_);
  nor (_29505_, _09403_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_29506_, _09403_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_29507_, _29506_, _29505_);
  and (_29508_, _16171_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_29510_, _16171_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_29511_, _29510_, _29508_);
  or (_29512_, _29511_, _29507_);
  or (_29513_, _29512_, _29504_);
  or (_29514_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_29515_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_29516_, _29515_, _29514_);
  or (_29517_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_29518_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_29519_, _29518_, _29517_);
  or (_29521_, _29519_, _29516_);
  and (_29522_, _08323_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_29523_, _08323_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_29524_, _29523_, _29522_);
  nand (_29525_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_29526_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_29527_, _29526_, _29525_);
  or (_29528_, _29527_, _29524_);
  or (_29529_, _29528_, _29521_);
  or (_29530_, _29529_, _29513_);
  and (property_invalid_dph, _29530_, _28766_);
  nand (_29532_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_29533_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_29534_, _29533_, _29532_);
  and (_29535_, _15613_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_29536_, \oc8051_golden_model_1.DPL [2], _30926_);
  or (_29537_, _29536_, _29535_);
  or (_29538_, _29537_, _29534_);
  and (_29539_, \oc8051_golden_model_1.DPL [0], _30918_);
  and (_29540_, _15429_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_29541_, _29540_, _29539_);
  and (_29542_, _15517_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_29543_, \oc8051_golden_model_1.DPL [1], _30922_);
  or (_29544_, _29543_, _29542_);
  or (_29545_, _29544_, _29541_);
  or (_29546_, _29545_, _29538_);
  or (_29547_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_29548_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_29549_, _29548_, _29547_);
  or (_29550_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_29553_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_29554_, _29553_, _29550_);
  or (_29555_, _29554_, _29549_);
  and (_29556_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_29557_, \oc8051_golden_model_1.DPL [7], _30637_);
  or (_29558_, _29557_, _29556_);
  nand (_29559_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_29560_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_29561_, _29560_, _29559_);
  or (_29562_, _29561_, _29558_);
  or (_29564_, _29562_, _29555_);
  or (_29565_, _29564_, _29546_);
  and (property_invalid_dpl, _29565_, _28766_);
  nand (_29566_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_29567_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_29568_, _29567_, _29566_);
  and (_29569_, _06826_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_29570_, \oc8051_golden_model_1.B [2], _29616_);
  or (_29571_, _29570_, _29569_);
  or (_29572_, _29571_, _29568_);
  and (_29574_, \oc8051_golden_model_1.B [0], _28327_);
  and (_29575_, _06820_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_29576_, _29575_, _29574_);
  and (_29577_, _06814_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29578_, \oc8051_golden_model_1.B [1], _28972_);
  or (_29579_, _29578_, _29577_);
  or (_29580_, _29579_, _29576_);
  or (_29581_, _29580_, _29572_);
  or (_29582_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_29583_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_29585_, _29583_, _29582_);
  or (_29586_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_29587_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_29588_, _29587_, _29586_);
  or (_29589_, _29588_, _29585_);
  and (_29590_, _06232_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_29591_, \oc8051_golden_model_1.B [7], _27213_);
  or (_29592_, _29591_, _29590_);
  nand (_29593_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_29594_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_29596_, _29594_, _29593_);
  or (_29597_, _29596_, _29592_);
  or (_29598_, _29597_, _29589_);
  or (_29599_, _29598_, _29581_);
  and (property_invalid_b_reg, _29599_, _28766_);
  nand (_29600_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_29601_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_29602_, _29601_, _29600_);
  and (_29603_, _06984_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_29604_, \oc8051_golden_model_1.ACC [2], _31140_);
  or (_29606_, _29604_, _29603_);
  or (_29607_, _29606_, _29602_);
  nor (_29608_, _02618_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_29609_, _02618_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_29610_, _29609_, _29608_);
  and (_29611_, _02549_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_29612_, _02549_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_29613_, _29612_, _29611_);
  or (_29614_, _29613_, _29610_);
  or (_29615_, _29614_, _29607_);
  or (_29617_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_29618_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_29619_, _29618_, _29617_);
  or (_29620_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_29621_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_29622_, _29621_, _29620_);
  or (_29623_, _29622_, _29619_);
  and (_29624_, _06833_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_29625_, _06833_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_29626_, _29625_, _29624_);
  nand (_29628_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_29629_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_29630_, _29629_, _29628_);
  or (_29631_, _29630_, _29626_);
  or (_29632_, _29631_, _29623_);
  or (_29633_, _29632_, _29615_);
  and (property_invalid_acc, _29633_, _28766_);
  nor (_29634_, _20594_, _35485_);
  and (_29635_, _20594_, _35485_);
  nand (_29636_, _20956_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_29638_, _20956_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_29639_, _29638_, _29636_);
  nand (_29640_, _22763_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_29641_, _22763_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_29642_, _29641_, _29640_);
  and (_29643_, _23440_, _30556_);
  nor (_29644_, _23440_, _30556_);
  and (_29645_, _23101_, _30550_);
  nor (_29646_, _23101_, _30550_);
  and (_29647_, _24741_, _30542_);
  and (_29649_, _25049_, _30573_);
  nor (_29650_, _25049_, _30573_);
  nand (_29651_, _09783_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_29652_, _09783_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_29653_, _29652_, _29651_);
  nand (_29654_, _24411_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_29655_, _24411_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_29656_, _29655_, _29654_);
  or (_29657_, _20195_, _35481_);
  nand (_29658_, _20195_, _35481_);
  and (_29660_, _29658_, _29657_);
  or (_29661_, _29660_, _29656_);
  or (_29662_, _29661_, _29653_);
  or (_29663_, _29662_, _29650_);
  or (_29664_, _29663_, _29649_);
  and (_29665_, _23748_, _30561_);
  nor (_29666_, _23748_, _30561_);
  or (_29667_, _29666_, _29665_);
  or (_29668_, _29667_, _29664_);
  or (_29669_, _29668_, _29647_);
  nor (_29671_, _24083_, _30546_);
  nor (_29672_, _24741_, _30542_);
  and (_29673_, _24083_, _30546_);
  or (_29674_, _29673_, _29672_);
  or (_29675_, _29674_, _29671_);
  or (_29676_, _29675_, _29669_);
  or (_29677_, _29676_, _29646_);
  or (_29678_, _29677_, _29645_);
  or (_29679_, _29678_, _29644_);
  or (_29680_, _29679_, _29643_);
  or (_29682_, _29680_, _29642_);
  nand (_29683_, _22048_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_29684_, _22048_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_29685_, _29684_, _29683_);
  nand (_29686_, _21318_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_29687_, _21318_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_29688_, _29687_, _29686_);
  or (_29689_, _29688_, _29685_);
  or (_29690_, _29689_, _29682_);
  and (_29691_, _21679_, _35496_);
  nor (_29693_, _21679_, _35496_);
  or (_29694_, _29693_, _29691_);
  or (_29695_, _29694_, _29690_);
  or (_29696_, _29695_, _29639_);
  nor (_29697_, _22404_, _35504_);
  and (_29698_, _22404_, _35504_);
  or (_29699_, _29698_, _29697_);
  or (_29700_, _29699_, _29696_);
  or (_29701_, _29700_, _29635_);
  or (_29702_, _29701_, _29634_);
  and (property_invalid_pc, _29702_, _28373_);
  buf (_36077_, _36029_);
  buf (_36118_, _36029_);
  buf (_00036_, _36029_);
  buf (_00078_, _36029_);
  buf (_00120_, _36029_);
  buf (_00162_, _36029_);
  buf (_00207_, _36029_);
  buf (_00253_, _36029_);
  buf (_00295_, _36029_);
  buf (_00339_, _36029_);
  buf (_00392_, _36029_);
  buf (_00445_, _36029_);
  buf (_00498_, _36029_);
  buf (_00551_, _36029_);
  buf (_00604_, _36029_);
  buf (_30875_, _30770_);
  buf (_30877_, _30771_);
  buf (_30890_, _30770_);
  buf (_30891_, _30771_);
  buf (_31200_, _30791_);
  buf (_31201_, _30792_);
  buf (_31202_, _30793_);
  buf (_31203_, _30794_);
  buf (_31204_, _30795_);
  buf (_31205_, _30797_);
  buf (_31206_, _30798_);
  buf (_31207_, _30799_);
  buf (_31209_, _30800_);
  buf (_31210_, _30801_);
  buf (_31211_, _30803_);
  buf (_31212_, _30804_);
  buf (_31213_, _30805_);
  buf (_31214_, _30806_);
  buf (_31266_, _30791_);
  buf (_31267_, _30792_);
  buf (_31268_, _30793_);
  buf (_31269_, _30794_);
  buf (_31270_, _30795_);
  buf (_31271_, _30797_);
  buf (_31272_, _30798_);
  buf (_31273_, _30799_);
  buf (_31275_, _30800_);
  buf (_31276_, _30801_);
  buf (_31277_, _30803_);
  buf (_31278_, _30804_);
  buf (_31279_, _30805_);
  buf (_31280_, _30806_);
  buf (_31605_, _31573_);
  buf (_31717_, _31573_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _36033_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _36036_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _36040_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _36043_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _36047_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _36051_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _36054_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _36026_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _36029_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _36080_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _36084_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _36087_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _36091_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _36095_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _36098_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _36102_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _36074_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _36077_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00343_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00347_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00351_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00355_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00359_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00363_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00367_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00336_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00339_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00396_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00400_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00404_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00408_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00412_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00416_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00420_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00389_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00392_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00449_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00453_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00457_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00461_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00465_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00469_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00473_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00442_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00445_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00502_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00506_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00510_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00514_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00518_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00522_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00526_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00495_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00498_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00555_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00559_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00563_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00567_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00571_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00575_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00579_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00548_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00551_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00608_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00612_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00616_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00620_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00624_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00628_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00632_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00601_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00604_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _36121_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _36125_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _36128_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00009_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00012_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00016_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00019_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _36115_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _36118_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00039_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00042_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00045_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00049_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00052_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00055_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00058_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00033_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00036_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00081_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00084_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00087_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00091_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00094_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00097_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00100_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00075_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00078_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00123_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00126_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00129_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00133_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00136_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00139_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00142_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00117_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00120_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00165_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00168_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00171_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00175_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00178_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00182_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00185_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00159_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00162_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00211_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00214_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00218_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00221_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00225_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00228_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00232_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00204_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00207_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00256_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00259_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00263_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00266_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00270_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00273_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00276_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00250_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00253_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00299_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00302_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00305_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00308_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00312_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00315_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00318_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00293_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00295_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _32708_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _32709_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _32710_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _32711_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _32712_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _32713_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _32715_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _32484_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _32697_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _32699_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _32700_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _32701_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _32702_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _32703_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _32704_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _32705_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _32686_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _32688_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _32689_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _32690_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _32691_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _32692_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _32694_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _32695_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _32675_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _32676_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _32678_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _32679_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _32680_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _32681_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _32682_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _32684_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _32664_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _32665_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _32666_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _32668_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _32669_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _32670_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _32671_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _32672_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _32653_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _32654_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _32655_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _32656_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _32658_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _32659_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _32660_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _32661_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _32642_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _32643_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _32644_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _32645_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _32647_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _32648_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _32649_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _32650_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _32631_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _32632_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _32633_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _32634_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _32635_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _32637_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _32638_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _32639_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _32619_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _32620_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _32621_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _32623_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _32624_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _32625_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _32626_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _32627_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _32608_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _32609_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _32610_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _32611_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _32613_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _32614_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _32615_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _32616_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _32598_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _32599_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _32600_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _32601_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _32602_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _32603_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _32604_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _32605_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _32587_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _32588_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _32589_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _32590_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _32591_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _32592_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _32593_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _32594_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _32575_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _32576_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _32577_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _32579_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _32580_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _32581_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _32582_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _32583_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _32564_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _32565_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _32566_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _32567_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _32568_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _32570_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _32571_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _32572_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _32552_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _32553_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _32554_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _32556_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _32557_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _32558_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _32559_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _32560_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _32540_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _32541_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _32543_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _32544_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _32545_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _32546_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _32547_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _32549_);
  dff (\oc8051_golden_model_1.B [0], _35155_);
  dff (\oc8051_golden_model_1.B [1], _35156_);
  dff (\oc8051_golden_model_1.B [2], _35157_);
  dff (\oc8051_golden_model_1.B [3], _35159_);
  dff (\oc8051_golden_model_1.B [4], _35160_);
  dff (\oc8051_golden_model_1.B [5], _35161_);
  dff (\oc8051_golden_model_1.B [6], _35162_);
  dff (\oc8051_golden_model_1.B [7], _32485_);
  dff (\oc8051_golden_model_1.ACC [0], _35164_);
  dff (\oc8051_golden_model_1.ACC [1], _35165_);
  dff (\oc8051_golden_model_1.ACC [2], _35166_);
  dff (\oc8051_golden_model_1.ACC [3], _35167_);
  dff (\oc8051_golden_model_1.ACC [4], _35168_);
  dff (\oc8051_golden_model_1.ACC [5], _35169_);
  dff (\oc8051_golden_model_1.ACC [6], _35170_);
  dff (\oc8051_golden_model_1.ACC [7], _32486_);
  dff (\oc8051_golden_model_1.DPL [0], _35172_);
  dff (\oc8051_golden_model_1.DPL [1], _35173_);
  dff (\oc8051_golden_model_1.DPL [2], _35174_);
  dff (\oc8051_golden_model_1.DPL [3], _35175_);
  dff (\oc8051_golden_model_1.DPL [4], _35176_);
  dff (\oc8051_golden_model_1.DPL [5], _35178_);
  dff (\oc8051_golden_model_1.DPL [6], _35179_);
  dff (\oc8051_golden_model_1.DPL [7], _32487_);
  dff (\oc8051_golden_model_1.DPH [0], _35180_);
  dff (\oc8051_golden_model_1.DPH [1], _35182_);
  dff (\oc8051_golden_model_1.DPH [2], _35183_);
  dff (\oc8051_golden_model_1.DPH [3], _35184_);
  dff (\oc8051_golden_model_1.DPH [4], _35185_);
  dff (\oc8051_golden_model_1.DPH [5], _35186_);
  dff (\oc8051_golden_model_1.DPH [6], _35187_);
  dff (\oc8051_golden_model_1.DPH [7], _32488_);
  dff (\oc8051_golden_model_1.IE [0], _35188_);
  dff (\oc8051_golden_model_1.IE [1], _35189_);
  dff (\oc8051_golden_model_1.IE [2], _35190_);
  dff (\oc8051_golden_model_1.IE [3], _35191_);
  dff (\oc8051_golden_model_1.IE [4], _35193_);
  dff (\oc8051_golden_model_1.IE [5], _35194_);
  dff (\oc8051_golden_model_1.IE [6], _35195_);
  dff (\oc8051_golden_model_1.IE [7], _32489_);
  dff (\oc8051_golden_model_1.IP [0], _35196_);
  dff (\oc8051_golden_model_1.IP [1], _35197_);
  dff (\oc8051_golden_model_1.IP [2], _35198_);
  dff (\oc8051_golden_model_1.IP [3], _35199_);
  dff (\oc8051_golden_model_1.IP [4], _35200_);
  dff (\oc8051_golden_model_1.IP [5], _35201_);
  dff (\oc8051_golden_model_1.IP [6], _35202_);
  dff (\oc8051_golden_model_1.IP [7], _32490_);
  dff (\oc8051_golden_model_1.P0 [0], _35204_);
  dff (\oc8051_golden_model_1.P0 [1], _35205_);
  dff (\oc8051_golden_model_1.P0 [2], _35206_);
  dff (\oc8051_golden_model_1.P0 [3], _35208_);
  dff (\oc8051_golden_model_1.P0 [4], _35209_);
  dff (\oc8051_golden_model_1.P0 [5], _35210_);
  dff (\oc8051_golden_model_1.P0 [6], _35211_);
  dff (\oc8051_golden_model_1.P0 [7], _32491_);
  dff (\oc8051_golden_model_1.P1 [0], _35213_);
  dff (\oc8051_golden_model_1.P1 [1], _35214_);
  dff (\oc8051_golden_model_1.P1 [2], _35215_);
  dff (\oc8051_golden_model_1.P1 [3], _35216_);
  dff (\oc8051_golden_model_1.P1 [4], _35217_);
  dff (\oc8051_golden_model_1.P1 [5], _35218_);
  dff (\oc8051_golden_model_1.P1 [6], _35219_);
  dff (\oc8051_golden_model_1.P1 [7], _32492_);
  dff (\oc8051_golden_model_1.P2 [0], _35221_);
  dff (\oc8051_golden_model_1.P2 [1], _35222_);
  dff (\oc8051_golden_model_1.P2 [2], _35223_);
  dff (\oc8051_golden_model_1.P2 [3], _35224_);
  dff (\oc8051_golden_model_1.P2 [4], _35225_);
  dff (\oc8051_golden_model_1.P2 [5], _35227_);
  dff (\oc8051_golden_model_1.P2 [6], _35228_);
  dff (\oc8051_golden_model_1.P2 [7], _32493_);
  dff (\oc8051_golden_model_1.P3 [0], _35229_);
  dff (\oc8051_golden_model_1.P3 [1], _35231_);
  dff (\oc8051_golden_model_1.P3 [2], _35232_);
  dff (\oc8051_golden_model_1.P3 [3], _35233_);
  dff (\oc8051_golden_model_1.P3 [4], _35234_);
  dff (\oc8051_golden_model_1.P3 [5], _35235_);
  dff (\oc8051_golden_model_1.P3 [6], _35236_);
  dff (\oc8051_golden_model_1.P3 [7], _32495_);
  dff (\oc8051_golden_model_1.PC [0], _35239_);
  dff (\oc8051_golden_model_1.PC [1], _35240_);
  dff (\oc8051_golden_model_1.PC [2], _35241_);
  dff (\oc8051_golden_model_1.PC [3], _35242_);
  dff (\oc8051_golden_model_1.PC [4], _35243_);
  dff (\oc8051_golden_model_1.PC [5], _35244_);
  dff (\oc8051_golden_model_1.PC [6], _35245_);
  dff (\oc8051_golden_model_1.PC [7], _35246_);
  dff (\oc8051_golden_model_1.PC [8], _35247_);
  dff (\oc8051_golden_model_1.PC [9], _35249_);
  dff (\oc8051_golden_model_1.PC [10], _35250_);
  dff (\oc8051_golden_model_1.PC [11], _35251_);
  dff (\oc8051_golden_model_1.PC [12], _35252_);
  dff (\oc8051_golden_model_1.PC [13], _35253_);
  dff (\oc8051_golden_model_1.PC [14], _35254_);
  dff (\oc8051_golden_model_1.PC [15], _32496_);
  dff (\oc8051_golden_model_1.PSW [0], _35256_);
  dff (\oc8051_golden_model_1.PSW [1], _35257_);
  dff (\oc8051_golden_model_1.PSW [2], _35258_);
  dff (\oc8051_golden_model_1.PSW [3], _35259_);
  dff (\oc8051_golden_model_1.PSW [4], _35260_);
  dff (\oc8051_golden_model_1.PSW [5], _35261_);
  dff (\oc8051_golden_model_1.PSW [6], _35262_);
  dff (\oc8051_golden_model_1.PSW [7], _32497_);
  dff (\oc8051_golden_model_1.PCON [0], _35264_);
  dff (\oc8051_golden_model_1.PCON [1], _35265_);
  dff (\oc8051_golden_model_1.PCON [2], _35266_);
  dff (\oc8051_golden_model_1.PCON [3], _35267_);
  dff (\oc8051_golden_model_1.PCON [4], _35268_);
  dff (\oc8051_golden_model_1.PCON [5], _35269_);
  dff (\oc8051_golden_model_1.PCON [6], _35270_);
  dff (\oc8051_golden_model_1.PCON [7], _32498_);
  dff (\oc8051_golden_model_1.SBUF [0], _35271_);
  dff (\oc8051_golden_model_1.SBUF [1], _35272_);
  dff (\oc8051_golden_model_1.SBUF [2], _35273_);
  dff (\oc8051_golden_model_1.SBUF [3], _35275_);
  dff (\oc8051_golden_model_1.SBUF [4], _35276_);
  dff (\oc8051_golden_model_1.SBUF [5], _35277_);
  dff (\oc8051_golden_model_1.SBUF [6], _35278_);
  dff (\oc8051_golden_model_1.SBUF [7], _32499_);
  dff (\oc8051_golden_model_1.SCON [0], _35279_);
  dff (\oc8051_golden_model_1.SCON [1], _35280_);
  dff (\oc8051_golden_model_1.SCON [2], _35281_);
  dff (\oc8051_golden_model_1.SCON [3], _35282_);
  dff (\oc8051_golden_model_1.SCON [4], _35283_);
  dff (\oc8051_golden_model_1.SCON [5], _35284_);
  dff (\oc8051_golden_model_1.SCON [6], _35286_);
  dff (\oc8051_golden_model_1.SCON [7], _32500_);
  dff (\oc8051_golden_model_1.SP [0], _35287_);
  dff (\oc8051_golden_model_1.SP [1], _35288_);
  dff (\oc8051_golden_model_1.SP [2], _35290_);
  dff (\oc8051_golden_model_1.SP [3], _35291_);
  dff (\oc8051_golden_model_1.SP [4], _35292_);
  dff (\oc8051_golden_model_1.SP [5], _35293_);
  dff (\oc8051_golden_model_1.SP [6], _35294_);
  dff (\oc8051_golden_model_1.SP [7], _32501_);
  dff (\oc8051_golden_model_1.TCON [0], _35295_);
  dff (\oc8051_golden_model_1.TCON [1], _35296_);
  dff (\oc8051_golden_model_1.TCON [2], _35297_);
  dff (\oc8051_golden_model_1.TCON [3], _35298_);
  dff (\oc8051_golden_model_1.TCON [4], _35299_);
  dff (\oc8051_golden_model_1.TCON [5], _35301_);
  dff (\oc8051_golden_model_1.TCON [6], _35302_);
  dff (\oc8051_golden_model_1.TCON [7], _32503_);
  dff (\oc8051_golden_model_1.TH0 [0], _35303_);
  dff (\oc8051_golden_model_1.TH0 [1], _35304_);
  dff (\oc8051_golden_model_1.TH0 [2], _35305_);
  dff (\oc8051_golden_model_1.TH0 [3], _35306_);
  dff (\oc8051_golden_model_1.TH0 [4], _35307_);
  dff (\oc8051_golden_model_1.TH0 [5], _35308_);
  dff (\oc8051_golden_model_1.TH0 [6], _35309_);
  dff (\oc8051_golden_model_1.TH0 [7], _32504_);
  dff (\oc8051_golden_model_1.TH1 [0], _35310_);
  dff (\oc8051_golden_model_1.TH1 [1], _35312_);
  dff (\oc8051_golden_model_1.TH1 [2], _35313_);
  dff (\oc8051_golden_model_1.TH1 [3], _35314_);
  dff (\oc8051_golden_model_1.TH1 [4], _35315_);
  dff (\oc8051_golden_model_1.TH1 [5], _35316_);
  dff (\oc8051_golden_model_1.TH1 [6], _35317_);
  dff (\oc8051_golden_model_1.TH1 [7], _32505_);
  dff (\oc8051_golden_model_1.TL0 [0], _35318_);
  dff (\oc8051_golden_model_1.TL0 [1], _35319_);
  dff (\oc8051_golden_model_1.TL0 [2], _35320_);
  dff (\oc8051_golden_model_1.TL0 [3], _35321_);
  dff (\oc8051_golden_model_1.TL0 [4], _35323_);
  dff (\oc8051_golden_model_1.TL0 [5], _35324_);
  dff (\oc8051_golden_model_1.TL0 [6], _35325_);
  dff (\oc8051_golden_model_1.TL0 [7], _32506_);
  dff (\oc8051_golden_model_1.TL1 [0], _35326_);
  dff (\oc8051_golden_model_1.TL1 [1], _35327_);
  dff (\oc8051_golden_model_1.TL1 [2], _35328_);
  dff (\oc8051_golden_model_1.TL1 [3], _35329_);
  dff (\oc8051_golden_model_1.TL1 [4], _35330_);
  dff (\oc8051_golden_model_1.TL1 [5], _35331_);
  dff (\oc8051_golden_model_1.TL1 [6], _35332_);
  dff (\oc8051_golden_model_1.TL1 [7], _32507_);
  dff (\oc8051_golden_model_1.TMOD [0], _35334_);
  dff (\oc8051_golden_model_1.TMOD [1], _35335_);
  dff (\oc8051_golden_model_1.TMOD [2], _35336_);
  dff (\oc8051_golden_model_1.TMOD [3], _35337_);
  dff (\oc8051_golden_model_1.TMOD [4], _35338_);
  dff (\oc8051_golden_model_1.TMOD [5], _35339_);
  dff (\oc8051_golden_model_1.TMOD [6], _35340_);
  dff (\oc8051_golden_model_1.TMOD [7], _32508_);
  dff (\oc8051_golden_model_1.P0INREG [0], _35342_);
  dff (\oc8051_golden_model_1.P0INREG [1], _35343_);
  dff (\oc8051_golden_model_1.P0INREG [2], _35344_);
  dff (\oc8051_golden_model_1.P0INREG [3], _35345_);
  dff (\oc8051_golden_model_1.P0INREG [4], _35346_);
  dff (\oc8051_golden_model_1.P0INREG [5], _35347_);
  dff (\oc8051_golden_model_1.P0INREG [6], _35349_);
  dff (\oc8051_golden_model_1.P0INREG [7], _32509_);
  dff (\oc8051_golden_model_1.P1INREG [0], _35350_);
  dff (\oc8051_golden_model_1.P1INREG [1], _35351_);
  dff (\oc8051_golden_model_1.P1INREG [2], _35353_);
  dff (\oc8051_golden_model_1.P1INREG [3], _35354_);
  dff (\oc8051_golden_model_1.P1INREG [4], _35355_);
  dff (\oc8051_golden_model_1.P1INREG [5], _35356_);
  dff (\oc8051_golden_model_1.P1INREG [6], _35357_);
  dff (\oc8051_golden_model_1.P1INREG [7], _32510_);
  dff (\oc8051_golden_model_1.P2INREG [0], _35359_);
  dff (\oc8051_golden_model_1.P2INREG [1], _35360_);
  dff (\oc8051_golden_model_1.P2INREG [2], _35361_);
  dff (\oc8051_golden_model_1.P2INREG [3], _35362_);
  dff (\oc8051_golden_model_1.P2INREG [4], _35363_);
  dff (\oc8051_golden_model_1.P2INREG [5], _35364_);
  dff (\oc8051_golden_model_1.P2INREG [6], _35365_);
  dff (\oc8051_golden_model_1.P2INREG [7], _32512_);
  dff (\oc8051_golden_model_1.P3INREG [0], _35367_);
  dff (\oc8051_golden_model_1.P3INREG [1], _35368_);
  dff (\oc8051_golden_model_1.P3INREG [2], _35369_);
  dff (\oc8051_golden_model_1.P3INREG [3], _35370_);
  dff (\oc8051_golden_model_1.P3INREG [4], _35372_);
  dff (\oc8051_golden_model_1.P3INREG [5], _35373_);
  dff (\oc8051_golden_model_1.P3INREG [6], _35374_);
  dff (\oc8051_golden_model_1.P3INREG [7], _32513_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03061_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03072_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03093_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03115_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03136_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _01083_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03147_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _01053_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03158_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03169_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03180_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03191_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03202_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03213_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03224_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01090_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02699_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _24753_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02900_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03104_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03315_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03516_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03717_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03918_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _04119_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04320_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04434_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04547_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04648_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04749_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04850_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04951_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _05052_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _26950_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _30783_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _30784_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _30785_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _30786_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _30787_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _30788_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _30789_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _30768_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _30791_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _30792_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _30793_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _30794_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _30795_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _30797_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _30798_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _30770_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _30799_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _30800_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _30801_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _30803_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _30804_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _30805_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _30806_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _30771_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04380_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _28683_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04383_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _28685_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04386_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _28687_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _28689_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04389_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _28691_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _28693_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04392_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _28695_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04395_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _28697_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _28699_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _28701_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04398_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _28704_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04401_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _04404_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _04464_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _04466_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04368_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _04469_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _04472_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04371_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _04475_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _04374_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _04478_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _04481_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _04484_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _04487_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _04490_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _04493_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _04496_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _04377_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _31573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _30941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _30942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _30943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _30944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _30945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _30946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _30947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _30948_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _30949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _30950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _30951_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _30952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _30953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _30954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _30956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _30832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _30960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _30961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _30962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _30963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _30964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _30965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _30966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _30967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _30968_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _30970_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _30971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _30972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _30973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _30974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _30975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _30833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _31153_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _31154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _31155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _31156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _31157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _31158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _31159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _31161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _31162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _31163_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _31164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _31165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _31166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _31167_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _31168_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _31169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _31170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _31172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _31173_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _31174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _31175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _31176_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _31177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _31178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _31179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _31180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _31181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _31183_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _31184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _31185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _31186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _30898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _30871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _31187_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _31188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _31189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _31190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _30873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _31191_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _31193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _31194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _31195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _31196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _31197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _31199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _30874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _31200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _31201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _31202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _31203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _31204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _31205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _31206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _30875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _31207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _31209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _31210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _31211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _31212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _31213_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _31214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _30877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _30878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _30879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _31215_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _31216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _31217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _31218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _31220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _31221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _31222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _30880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _31223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _31224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _31225_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _31226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _31227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _31228_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _31229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _31231_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _31232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _31233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _31234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _31235_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _31236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _31237_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _31238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _30881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _31239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _31240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _31242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _31243_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _31244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _31245_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _31246_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _31247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _31248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _31249_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _31250_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _31251_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _31253_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _31254_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _31255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _30883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _30884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _30886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _30885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _31256_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _31257_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _31258_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _31259_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _31260_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _31261_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _31262_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _30888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _31264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _31265_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _30889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _31266_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _31267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _31268_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _31269_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _31270_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _31271_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _31272_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _30890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _31273_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _31275_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _31276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _31277_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _31278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _31279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _31280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _30891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _30892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _31281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _31282_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _31283_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _31284_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _31286_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _31287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _31288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _30893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _30895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _30896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _31289_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _31290_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _31291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _30897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _31292_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _31293_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _31294_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _31295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _31296_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _31297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _31298_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _31299_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _31300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _31301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _31302_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _31303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _31304_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _31305_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _31307_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _31308_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _31309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _31310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _31311_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _31312_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _31313_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _31314_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _31315_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _31316_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _31318_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _31319_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _31320_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _31321_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _31322_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _31323_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _31324_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _30899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _31325_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _31326_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _31327_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _31329_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _31330_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _31331_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _31332_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _30900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _30901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _30903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _31333_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _31334_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _31335_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _31336_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _31337_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _31338_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _31340_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _31341_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _31342_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _31343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _31344_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _31345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _31346_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _31347_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _31348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _30904_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _30905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _30906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _30907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _31349_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _31351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _31352_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _31353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _31354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _31355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _31356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _31357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _31358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _31359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _31360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _31362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _31363_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _31364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _31365_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _30908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _30909_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _31715_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _31733_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _31734_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _31736_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _31737_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _31738_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _31739_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _31740_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _31716_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _31717_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _31741_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _31742_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _31718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _33693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _33698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _33703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _33709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _33714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _33719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _33724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _33727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _33764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _33768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _33771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _33775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _33778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _33782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _33785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _33788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _33939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _33942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _33946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _33949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _33953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _33956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _33960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _33962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _33908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _33912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _33915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _33919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _33922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _33926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _33929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _33932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _33880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _33884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _33887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _33891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _33894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _33898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _33901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _33904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _33852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _33855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _33859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _33862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _33866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _33869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _33873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _33876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _33824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _33827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _33831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _33834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _33838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _33841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _33845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _33848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _33793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _33797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _33800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _33804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _33807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _33811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _33814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _33817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _33734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _33737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _33741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _33744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _33748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _33751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _33755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _33757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _33967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _33970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _33974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _33977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _33981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _33984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _33988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _33990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _34120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _34124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _34128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _34132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _34136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _34139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _34143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _34146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _34090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _34094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _34098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _34102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _34106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _34109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _34113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _34115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _34058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _34062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _34066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _34070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _34074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _34078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _34082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _34085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _34025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _34029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _34033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _34037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _34041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _34045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _34049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _34052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _33994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _33997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _34001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _34005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _34009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _34013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _34017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _34020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _34151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _34155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _34159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _34162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _34166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _34170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _34174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _33450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _36008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _36010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _36012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _36013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _36015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _36017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _36019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _33440_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _31601_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _31603_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _31664_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _31666_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _31667_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _31668_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _31669_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _31670_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _31671_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _31604_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _31605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24356_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24368_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24380_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _09006_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _09017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _09028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _09039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13659_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _33315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _33317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _33319_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _33321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _33322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _33324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _33326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _30230_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _33328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _33330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _33332_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _33333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _33335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _33337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _33339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _30233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _33341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _33343_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _33344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _33346_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _33348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _33350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _33352_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _30236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _33354_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _33355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _33357_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _33359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _33361_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _33363_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _33365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _30239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21654_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09611_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.SBUF_next [0], \oc8051_golden_model_1.SBUF [0]);
  buf(\oc8051_golden_model_1.SBUF_next [1], \oc8051_golden_model_1.SBUF [1]);
  buf(\oc8051_golden_model_1.SBUF_next [2], \oc8051_golden_model_1.SBUF [2]);
  buf(\oc8051_golden_model_1.SBUF_next [3], \oc8051_golden_model_1.SBUF [3]);
  buf(\oc8051_golden_model_1.SBUF_next [4], \oc8051_golden_model_1.SBUF [4]);
  buf(\oc8051_golden_model_1.SBUF_next [5], \oc8051_golden_model_1.SBUF [5]);
  buf(\oc8051_golden_model_1.SBUF_next [6], \oc8051_golden_model_1.SBUF [6]);
  buf(\oc8051_golden_model_1.SBUF_next [7], \oc8051_golden_model_1.SBUF [7]);
  buf(\oc8051_golden_model_1.SCON_next [0], \oc8051_golden_model_1.SCON [0]);
  buf(\oc8051_golden_model_1.SCON_next [1], \oc8051_golden_model_1.SCON [1]);
  buf(\oc8051_golden_model_1.SCON_next [2], \oc8051_golden_model_1.SCON [2]);
  buf(\oc8051_golden_model_1.SCON_next [3], \oc8051_golden_model_1.SCON [3]);
  buf(\oc8051_golden_model_1.SCON_next [4], \oc8051_golden_model_1.SCON [4]);
  buf(\oc8051_golden_model_1.SCON_next [5], \oc8051_golden_model_1.SCON [5]);
  buf(\oc8051_golden_model_1.SCON_next [6], \oc8051_golden_model_1.SCON [6]);
  buf(\oc8051_golden_model_1.SCON_next [7], \oc8051_golden_model_1.SCON [7]);
  buf(\oc8051_golden_model_1.PCON_next [0], \oc8051_golden_model_1.PCON [0]);
  buf(\oc8051_golden_model_1.PCON_next [1], \oc8051_golden_model_1.PCON [1]);
  buf(\oc8051_golden_model_1.PCON_next [2], \oc8051_golden_model_1.PCON [2]);
  buf(\oc8051_golden_model_1.PCON_next [3], \oc8051_golden_model_1.PCON [3]);
  buf(\oc8051_golden_model_1.PCON_next [4], \oc8051_golden_model_1.PCON [4]);
  buf(\oc8051_golden_model_1.PCON_next [5], \oc8051_golden_model_1.PCON [5]);
  buf(\oc8051_golden_model_1.PCON_next [6], \oc8051_golden_model_1.PCON [6]);
  buf(\oc8051_golden_model_1.PCON_next [7], \oc8051_golden_model_1.PCON [7]);
  buf(\oc8051_golden_model_1.TCON_next [0], \oc8051_golden_model_1.TCON [0]);
  buf(\oc8051_golden_model_1.TCON_next [1], \oc8051_golden_model_1.TCON [1]);
  buf(\oc8051_golden_model_1.TCON_next [2], \oc8051_golden_model_1.TCON [2]);
  buf(\oc8051_golden_model_1.TCON_next [3], \oc8051_golden_model_1.TCON [3]);
  buf(\oc8051_golden_model_1.TCON_next [4], \oc8051_golden_model_1.TCON [4]);
  buf(\oc8051_golden_model_1.TCON_next [5], \oc8051_golden_model_1.TCON [5]);
  buf(\oc8051_golden_model_1.TCON_next [6], \oc8051_golden_model_1.TCON [6]);
  buf(\oc8051_golden_model_1.TCON_next [7], \oc8051_golden_model_1.TCON [7]);
  buf(\oc8051_golden_model_1.TL0_next [0], \oc8051_golden_model_1.TL0 [0]);
  buf(\oc8051_golden_model_1.TL0_next [1], \oc8051_golden_model_1.TL0 [1]);
  buf(\oc8051_golden_model_1.TL0_next [2], \oc8051_golden_model_1.TL0 [2]);
  buf(\oc8051_golden_model_1.TL0_next [3], \oc8051_golden_model_1.TL0 [3]);
  buf(\oc8051_golden_model_1.TL0_next [4], \oc8051_golden_model_1.TL0 [4]);
  buf(\oc8051_golden_model_1.TL0_next [5], \oc8051_golden_model_1.TL0 [5]);
  buf(\oc8051_golden_model_1.TL0_next [6], \oc8051_golden_model_1.TL0 [6]);
  buf(\oc8051_golden_model_1.TL0_next [7], \oc8051_golden_model_1.TL0 [7]);
  buf(\oc8051_golden_model_1.TL1_next [0], \oc8051_golden_model_1.TL1 [0]);
  buf(\oc8051_golden_model_1.TL1_next [1], \oc8051_golden_model_1.TL1 [1]);
  buf(\oc8051_golden_model_1.TL1_next [2], \oc8051_golden_model_1.TL1 [2]);
  buf(\oc8051_golden_model_1.TL1_next [3], \oc8051_golden_model_1.TL1 [3]);
  buf(\oc8051_golden_model_1.TL1_next [4], \oc8051_golden_model_1.TL1 [4]);
  buf(\oc8051_golden_model_1.TL1_next [5], \oc8051_golden_model_1.TL1 [5]);
  buf(\oc8051_golden_model_1.TL1_next [6], \oc8051_golden_model_1.TL1 [6]);
  buf(\oc8051_golden_model_1.TL1_next [7], \oc8051_golden_model_1.TL1 [7]);
  buf(\oc8051_golden_model_1.TH0_next [0], \oc8051_golden_model_1.TH0 [0]);
  buf(\oc8051_golden_model_1.TH0_next [1], \oc8051_golden_model_1.TH0 [1]);
  buf(\oc8051_golden_model_1.TH0_next [2], \oc8051_golden_model_1.TH0 [2]);
  buf(\oc8051_golden_model_1.TH0_next [3], \oc8051_golden_model_1.TH0 [3]);
  buf(\oc8051_golden_model_1.TH0_next [4], \oc8051_golden_model_1.TH0 [4]);
  buf(\oc8051_golden_model_1.TH0_next [5], \oc8051_golden_model_1.TH0 [5]);
  buf(\oc8051_golden_model_1.TH0_next [6], \oc8051_golden_model_1.TH0 [6]);
  buf(\oc8051_golden_model_1.TH0_next [7], \oc8051_golden_model_1.TH0 [7]);
  buf(\oc8051_golden_model_1.TH1_next [0], \oc8051_golden_model_1.TH1 [0]);
  buf(\oc8051_golden_model_1.TH1_next [1], \oc8051_golden_model_1.TH1 [1]);
  buf(\oc8051_golden_model_1.TH1_next [2], \oc8051_golden_model_1.TH1 [2]);
  buf(\oc8051_golden_model_1.TH1_next [3], \oc8051_golden_model_1.TH1 [3]);
  buf(\oc8051_golden_model_1.TH1_next [4], \oc8051_golden_model_1.TH1 [4]);
  buf(\oc8051_golden_model_1.TH1_next [5], \oc8051_golden_model_1.TH1 [5]);
  buf(\oc8051_golden_model_1.TH1_next [6], \oc8051_golden_model_1.TH1 [6]);
  buf(\oc8051_golden_model_1.TH1_next [7], \oc8051_golden_model_1.TH1 [7]);
  buf(\oc8051_golden_model_1.TMOD_next [0], \oc8051_golden_model_1.TMOD [0]);
  buf(\oc8051_golden_model_1.TMOD_next [1], \oc8051_golden_model_1.TMOD [1]);
  buf(\oc8051_golden_model_1.TMOD_next [2], \oc8051_golden_model_1.TMOD [2]);
  buf(\oc8051_golden_model_1.TMOD_next [3], \oc8051_golden_model_1.TMOD [3]);
  buf(\oc8051_golden_model_1.TMOD_next [4], \oc8051_golden_model_1.TMOD [4]);
  buf(\oc8051_golden_model_1.TMOD_next [5], \oc8051_golden_model_1.TMOD [5]);
  buf(\oc8051_golden_model_1.TMOD_next [6], \oc8051_golden_model_1.TMOD [6]);
  buf(\oc8051_golden_model_1.TMOD_next [7], \oc8051_golden_model_1.TMOD [7]);
  buf(\oc8051_golden_model_1.IE_next [0], \oc8051_golden_model_1.IE [0]);
  buf(\oc8051_golden_model_1.IE_next [1], \oc8051_golden_model_1.IE [1]);
  buf(\oc8051_golden_model_1.IE_next [2], \oc8051_golden_model_1.IE [2]);
  buf(\oc8051_golden_model_1.IE_next [3], \oc8051_golden_model_1.IE [3]);
  buf(\oc8051_golden_model_1.IE_next [4], \oc8051_golden_model_1.IE [4]);
  buf(\oc8051_golden_model_1.IE_next [5], \oc8051_golden_model_1.IE [5]);
  buf(\oc8051_golden_model_1.IE_next [6], \oc8051_golden_model_1.IE [6]);
  buf(\oc8051_golden_model_1.IE_next [7], \oc8051_golden_model_1.IE [7]);
  buf(\oc8051_golden_model_1.IP_next [0], \oc8051_golden_model_1.IP [0]);
  buf(\oc8051_golden_model_1.IP_next [1], \oc8051_golden_model_1.IP [1]);
  buf(\oc8051_golden_model_1.IP_next [2], \oc8051_golden_model_1.IP [2]);
  buf(\oc8051_golden_model_1.IP_next [3], \oc8051_golden_model_1.IP [3]);
  buf(\oc8051_golden_model_1.IP_next [4], \oc8051_golden_model_1.IP [4]);
  buf(\oc8051_golden_model_1.IP_next [5], \oc8051_golden_model_1.IP [5]);
  buf(\oc8051_golden_model_1.IP_next [6], \oc8051_golden_model_1.IP [6]);
  buf(\oc8051_golden_model_1.IP_next [7], \oc8051_golden_model_1.IP [7]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1269 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1286 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1335 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1376 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1376 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1376 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1376 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1431 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1431 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1431 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1431 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1481 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1467 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1467 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1481 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1481 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1481 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1561 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1597 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1597 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1597 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1597 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1630 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1630 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1630 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1630 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1663 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1663 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1663 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1663 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1712 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1712 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1712 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1712 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1712 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1712 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1712 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1757 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1774 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1791 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1791 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1822 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1822 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1822 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1822 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1822 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1822 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1822 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1867 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1884 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1901 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1901 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n1994 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2011 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2028 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2028 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2053 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2069 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2100 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2069 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2126 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2126 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2069 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2330 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2330 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2330 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2330 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2360 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2360 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2360 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2360 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2390 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2390 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2390 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2390 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2390 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2390 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2390 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2390 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2425 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2428 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2456 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2456 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2462 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2493 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2501 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2509 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2566 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2608 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2608 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2691 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2691 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2713 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2713 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2732 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2733 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2608 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2608 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2750 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2751 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2751 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2751 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2751 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2751 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2751 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2751 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1046 , \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1063 , \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1146 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1146 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1146 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1148 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1148 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1148 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1150 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1150 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1150 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1150 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1151 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1151 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1151 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1151 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1152 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1152 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1152 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1153 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1153 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1153 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1153 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1154 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1154 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1154 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1154 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1155 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1155 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1156 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1156 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1156 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1156 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1202 , \oc8051_golden_model_1.n2428 [7]);
  buf(\oc8051_golden_model_1.n1244 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1245 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1245 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1245 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1245 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1245 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1245 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1245 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1245 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1245 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1246 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1246 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1246 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1247 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1247 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1247 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1247 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1247 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1247 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1247 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1249 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1249 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1249 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1251 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1251 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1252 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1252 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1252 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1252 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1252 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1252 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1252 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1252 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1253 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1253 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1253 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1253 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1253 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1253 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1253 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1255 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1258 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1268 , \oc8051_golden_model_1.n1269 [0]);
  buf(\oc8051_golden_model_1.n1269 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1269 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1269 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1269 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1269 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1269 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1269 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1285 , \oc8051_golden_model_1.n1286 [0]);
  buf(\oc8051_golden_model_1.n1286 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1286 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1286 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1286 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1286 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1286 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1286 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1317 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n1317 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n1317 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n1317 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n1317 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n1317 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n1317 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n1317 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n1317 [8], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1317 [9], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1317 [10], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1317 [11], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1317 [12], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.n1317 [13], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.n1317 [14], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.n1317 [15], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n1319 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1319 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1319 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1319 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1319 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1319 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1319 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1319 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1321 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1322 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1324 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1334 , \oc8051_golden_model_1.n1335 [0]);
  buf(\oc8051_golden_model_1.n1335 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1335 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1335 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1335 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1335 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1335 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1335 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1337 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1337 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1337 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1337 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1337 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1337 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1337 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1337 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1341 [8], \oc8051_golden_model_1.n1376 [7]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1376 [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1344 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1344 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1344 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1344 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1344 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1348 [4], \oc8051_golden_model_1.n1376 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1376 [6]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1350 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1350 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1350 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1350 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1376 [2]);
  buf(\oc8051_golden_model_1.n1359 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1359 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1359 [2], \oc8051_golden_model_1.n1376 [2]);
  buf(\oc8051_golden_model_1.n1359 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1359 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1359 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1359 [6], \oc8051_golden_model_1.n1376 [6]);
  buf(\oc8051_golden_model_1.n1359 [7], \oc8051_golden_model_1.n1376 [7]);
  buf(\oc8051_golden_model_1.n1360 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1360 [1], \oc8051_golden_model_1.n1376 [2]);
  buf(\oc8051_golden_model_1.n1360 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1360 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1360 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1360 [5], \oc8051_golden_model_1.n1376 [6]);
  buf(\oc8051_golden_model_1.n1360 [6], \oc8051_golden_model_1.n1376 [7]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1376 [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1398 [8], \oc8051_golden_model_1.n1431 [7]);
  buf(\oc8051_golden_model_1.n1399 , \oc8051_golden_model_1.n1431 [7]);
  buf(\oc8051_golden_model_1.n1404 [4], \oc8051_golden_model_1.n1431 [6]);
  buf(\oc8051_golden_model_1.n1405 , \oc8051_golden_model_1.n1431 [6]);
  buf(\oc8051_golden_model_1.n1413 , \oc8051_golden_model_1.n1431 [2]);
  buf(\oc8051_golden_model_1.n1414 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1414 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1414 [2], \oc8051_golden_model_1.n1431 [2]);
  buf(\oc8051_golden_model_1.n1414 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1414 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1414 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1414 [6], \oc8051_golden_model_1.n1431 [6]);
  buf(\oc8051_golden_model_1.n1414 [7], \oc8051_golden_model_1.n1431 [7]);
  buf(\oc8051_golden_model_1.n1415 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1415 [1], \oc8051_golden_model_1.n1431 [2]);
  buf(\oc8051_golden_model_1.n1415 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1415 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1415 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1415 [5], \oc8051_golden_model_1.n1431 [6]);
  buf(\oc8051_golden_model_1.n1415 [6], \oc8051_golden_model_1.n1431 [7]);
  buf(\oc8051_golden_model_1.n1430 , \oc8051_golden_model_1.n1431 [0]);
  buf(\oc8051_golden_model_1.n1431 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1431 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1431 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1431 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1433 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n1433 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n1433 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n1433 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n1433 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n1433 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n1433 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n1433 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n1433 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1435 [8], \oc8051_golden_model_1.n1467 [7]);
  buf(\oc8051_golden_model_1.n1436 , \oc8051_golden_model_1.n1467 [7]);
  buf(\oc8051_golden_model_1.n1437 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n1437 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n1437 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n1437 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n1438 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n1438 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n1438 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n1438 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n1438 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1441 , \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1442 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n1442 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n1442 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n1442 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n1442 [4], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n1442 [5], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n1442 [6], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n1442 [7], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n1442 [8], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n1449 , \oc8051_golden_model_1.n1467 [2]);
  buf(\oc8051_golden_model_1.n1450 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1450 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1450 [2], \oc8051_golden_model_1.n1467 [2]);
  buf(\oc8051_golden_model_1.n1450 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1450 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1450 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1450 [6], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1450 [7], \oc8051_golden_model_1.n1467 [7]);
  buf(\oc8051_golden_model_1.n1451 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1451 [1], \oc8051_golden_model_1.n1467 [2]);
  buf(\oc8051_golden_model_1.n1451 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1451 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1451 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1451 [5], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1451 [6], \oc8051_golden_model_1.n1467 [7]);
  buf(\oc8051_golden_model_1.n1466 , \oc8051_golden_model_1.n1481 [0]);
  buf(\oc8051_golden_model_1.n1467 [0], \oc8051_golden_model_1.n1481 [0]);
  buf(\oc8051_golden_model_1.n1467 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1467 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1467 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1467 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1467 [6], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1470 [8], \oc8051_golden_model_1.n1481 [7]);
  buf(\oc8051_golden_model_1.n1471 , \oc8051_golden_model_1.n1481 [7]);
  buf(\oc8051_golden_model_1.n1478 , \oc8051_golden_model_1.n1481 [2]);
  buf(\oc8051_golden_model_1.n1479 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1479 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1479 [2], \oc8051_golden_model_1.n1481 [2]);
  buf(\oc8051_golden_model_1.n1479 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1479 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1479 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1479 [6], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1479 [7], \oc8051_golden_model_1.n1481 [7]);
  buf(\oc8051_golden_model_1.n1480 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1480 [1], \oc8051_golden_model_1.n1481 [2]);
  buf(\oc8051_golden_model_1.n1480 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1480 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1480 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1480 [5], \oc8051_golden_model_1.n1481 [6]);
  buf(\oc8051_golden_model_1.n1480 [6], \oc8051_golden_model_1.n1481 [7]);
  buf(\oc8051_golden_model_1.n1481 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1481 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1481 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1481 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1483 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1483 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1483 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1483 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1483 [4], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.n1483 [5], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.n1483 [6], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.n1483 [7], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n1483 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1485 [8], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1486 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1487 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1487 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1487 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1490 , \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1491 [0], \oc8051_golden_model_1.n2616 );
  buf(\oc8051_golden_model_1.n1491 [1], \oc8051_golden_model_1.n2615 );
  buf(\oc8051_golden_model_1.n1491 [2], \oc8051_golden_model_1.n2614 );
  buf(\oc8051_golden_model_1.n1491 [3], \oc8051_golden_model_1.n2613 );
  buf(\oc8051_golden_model_1.n1491 [4], \oc8051_golden_model_1.n2612 );
  buf(\oc8051_golden_model_1.n1491 [5], \oc8051_golden_model_1.n2611 );
  buf(\oc8051_golden_model_1.n1491 [6], \oc8051_golden_model_1.n2610 );
  buf(\oc8051_golden_model_1.n1491 [7], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n1491 [8], \oc8051_golden_model_1.n2609 );
  buf(\oc8051_golden_model_1.n1498 , \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1499 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1499 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1499 [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1499 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1499 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1499 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1499 [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1499 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1500 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1500 [1], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1500 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1500 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1500 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1500 [5], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1500 [6], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1515 , \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.n1516 [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.n1516 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1516 [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1516 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1516 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1516 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1516 [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1516 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1518 [4], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1519 , \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1520 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1520 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1520 [2], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1520 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1520 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1520 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1520 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.n1522 [2]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1524 [8], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1532 , \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1533 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1533 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1533 [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1533 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1533 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1533 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1533 [6], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1533 [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1534 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1534 [1], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1534 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1534 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1534 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1534 [5], \oc8051_golden_model_1.n1535 [6]);
  buf(\oc8051_golden_model_1.n1534 [6], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1535 [0], \oc8051_golden_model_1.n1538 [0]);
  buf(\oc8051_golden_model_1.n1535 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1535 [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1535 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1535 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1535 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1535 [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1536 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1536 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1536 [2], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1536 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1536 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1536 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1536 [6], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1536 [7], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1537 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1537 [1], \oc8051_golden_model_1.n1538 [2]);
  buf(\oc8051_golden_model_1.n1537 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1537 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1537 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1537 [5], \oc8051_golden_model_1.n1538 [6]);
  buf(\oc8051_golden_model_1.n1537 [6], \oc8051_golden_model_1.n1538 [7]);
  buf(\oc8051_golden_model_1.n1538 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1538 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1538 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1538 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1541 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1541 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1542 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1543 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1543 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1544 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1544 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1544 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1545 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1545 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1545 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1545 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1545 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1545 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1546 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1547 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1548 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1550 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1552 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1553 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1560 , \oc8051_golden_model_1.n1561 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1562 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1562 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1565 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1565 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.n1597 [7]);
  buf(\oc8051_golden_model_1.n1568 , \oc8051_golden_model_1.n1597 [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1569 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1569 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1569 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.n1597 [6]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.n1597 [6]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.n1597 [2]);
  buf(\oc8051_golden_model_1.n1580 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1580 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1580 [2], \oc8051_golden_model_1.n1597 [2]);
  buf(\oc8051_golden_model_1.n1580 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1580 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1580 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1580 [6], \oc8051_golden_model_1.n1597 [6]);
  buf(\oc8051_golden_model_1.n1580 [7], \oc8051_golden_model_1.n1597 [7]);
  buf(\oc8051_golden_model_1.n1581 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1581 [1], \oc8051_golden_model_1.n1597 [2]);
  buf(\oc8051_golden_model_1.n1581 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1581 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1581 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1581 [5], \oc8051_golden_model_1.n1597 [6]);
  buf(\oc8051_golden_model_1.n1581 [6], \oc8051_golden_model_1.n1597 [7]);
  buf(\oc8051_golden_model_1.n1596 , \oc8051_golden_model_1.n1597 [0]);
  buf(\oc8051_golden_model_1.n1597 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1597 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1597 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1597 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1601 [8], \oc8051_golden_model_1.n1630 [7]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1630 [7]);
  buf(\oc8051_golden_model_1.n1604 [4], \oc8051_golden_model_1.n1630 [6]);
  buf(\oc8051_golden_model_1.n1605 , \oc8051_golden_model_1.n1630 [6]);
  buf(\oc8051_golden_model_1.n1612 , \oc8051_golden_model_1.n1630 [2]);
  buf(\oc8051_golden_model_1.n1613 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1613 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1613 [2], \oc8051_golden_model_1.n1630 [2]);
  buf(\oc8051_golden_model_1.n1613 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1613 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1613 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1613 [6], \oc8051_golden_model_1.n1630 [6]);
  buf(\oc8051_golden_model_1.n1613 [7], \oc8051_golden_model_1.n1630 [7]);
  buf(\oc8051_golden_model_1.n1614 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1614 [1], \oc8051_golden_model_1.n1630 [2]);
  buf(\oc8051_golden_model_1.n1614 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1614 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1614 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1614 [5], \oc8051_golden_model_1.n1630 [6]);
  buf(\oc8051_golden_model_1.n1614 [6], \oc8051_golden_model_1.n1630 [7]);
  buf(\oc8051_golden_model_1.n1629 , \oc8051_golden_model_1.n1630 [0]);
  buf(\oc8051_golden_model_1.n1630 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1630 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1630 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1630 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1634 [8], \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.n1637 [4], \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.n1638 , \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.n1645 , \oc8051_golden_model_1.n1663 [2]);
  buf(\oc8051_golden_model_1.n1646 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1646 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1646 [2], \oc8051_golden_model_1.n1663 [2]);
  buf(\oc8051_golden_model_1.n1646 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1646 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1646 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1646 [6], \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.n1646 [7], \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.n1647 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1647 [1], \oc8051_golden_model_1.n1663 [2]);
  buf(\oc8051_golden_model_1.n1647 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1647 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1647 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1647 [5], \oc8051_golden_model_1.n1663 [6]);
  buf(\oc8051_golden_model_1.n1647 [6], \oc8051_golden_model_1.n1663 [7]);
  buf(\oc8051_golden_model_1.n1662 , \oc8051_golden_model_1.n1663 [0]);
  buf(\oc8051_golden_model_1.n1663 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1663 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1663 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1667 [8], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.n1670 [4], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.n1678 , \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.n1679 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1679 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1679 [2], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.n1679 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1679 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1679 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1679 [6], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.n1679 [7], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.n1696 [2]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.n1696 [6]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.n1696 [7]);
  buf(\oc8051_golden_model_1.n1695 , \oc8051_golden_model_1.n1696 [0]);
  buf(\oc8051_golden_model_1.n1696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1710 [1], \oc8051_golden_model_1.n1712 [1]);
  buf(\oc8051_golden_model_1.n1710 [2], \oc8051_golden_model_1.n1712 [2]);
  buf(\oc8051_golden_model_1.n1710 [3], \oc8051_golden_model_1.n1712 [3]);
  buf(\oc8051_golden_model_1.n1710 [4], \oc8051_golden_model_1.n1712 [4]);
  buf(\oc8051_golden_model_1.n1710 [5], \oc8051_golden_model_1.n1712 [5]);
  buf(\oc8051_golden_model_1.n1710 [6], \oc8051_golden_model_1.n1712 [6]);
  buf(\oc8051_golden_model_1.n1710 [7], \oc8051_golden_model_1.n1712 [7]);
  buf(\oc8051_golden_model_1.n1711 [0], \oc8051_golden_model_1.n1712 [1]);
  buf(\oc8051_golden_model_1.n1711 [1], \oc8051_golden_model_1.n1712 [2]);
  buf(\oc8051_golden_model_1.n1711 [2], \oc8051_golden_model_1.n1712 [3]);
  buf(\oc8051_golden_model_1.n1711 [3], \oc8051_golden_model_1.n1712 [4]);
  buf(\oc8051_golden_model_1.n1711 [4], \oc8051_golden_model_1.n1712 [5]);
  buf(\oc8051_golden_model_1.n1711 [5], \oc8051_golden_model_1.n1712 [6]);
  buf(\oc8051_golden_model_1.n1711 [6], \oc8051_golden_model_1.n1712 [7]);
  buf(\oc8051_golden_model_1.n1712 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n1756 , \oc8051_golden_model_1.n1757 [0]);
  buf(\oc8051_golden_model_1.n1757 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1757 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1757 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1757 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1757 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1757 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1757 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1773 , \oc8051_golden_model_1.n1774 [0]);
  buf(\oc8051_golden_model_1.n1774 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1774 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1774 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1774 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1774 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1774 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1774 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1790 , \oc8051_golden_model_1.n1791 [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1807 , \oc8051_golden_model_1.n1808 [0]);
  buf(\oc8051_golden_model_1.n1808 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1808 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1808 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1808 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1808 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1808 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1808 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1820 [1], \oc8051_golden_model_1.n1822 [1]);
  buf(\oc8051_golden_model_1.n1820 [2], \oc8051_golden_model_1.n1822 [2]);
  buf(\oc8051_golden_model_1.n1820 [3], \oc8051_golden_model_1.n1822 [3]);
  buf(\oc8051_golden_model_1.n1820 [4], \oc8051_golden_model_1.n1822 [4]);
  buf(\oc8051_golden_model_1.n1820 [5], \oc8051_golden_model_1.n1822 [5]);
  buf(\oc8051_golden_model_1.n1820 [6], \oc8051_golden_model_1.n1822 [6]);
  buf(\oc8051_golden_model_1.n1820 [7], \oc8051_golden_model_1.n1822 [7]);
  buf(\oc8051_golden_model_1.n1821 [0], \oc8051_golden_model_1.n1822 [1]);
  buf(\oc8051_golden_model_1.n1821 [1], \oc8051_golden_model_1.n1822 [2]);
  buf(\oc8051_golden_model_1.n1821 [2], \oc8051_golden_model_1.n1822 [3]);
  buf(\oc8051_golden_model_1.n1821 [3], \oc8051_golden_model_1.n1822 [4]);
  buf(\oc8051_golden_model_1.n1821 [4], \oc8051_golden_model_1.n1822 [5]);
  buf(\oc8051_golden_model_1.n1821 [5], \oc8051_golden_model_1.n1822 [6]);
  buf(\oc8051_golden_model_1.n1821 [6], \oc8051_golden_model_1.n1822 [7]);
  buf(\oc8051_golden_model_1.n1822 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n1866 , \oc8051_golden_model_1.n1867 [0]);
  buf(\oc8051_golden_model_1.n1867 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1867 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1867 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1867 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1867 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1867 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1867 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1883 , \oc8051_golden_model_1.n1884 [0]);
  buf(\oc8051_golden_model_1.n1884 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1884 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1884 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1884 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1884 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1884 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1884 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1900 , \oc8051_golden_model_1.n1901 [0]);
  buf(\oc8051_golden_model_1.n1901 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1901 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1901 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1901 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1901 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1901 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1901 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1917 , \oc8051_golden_model_1.n1918 [0]);
  buf(\oc8051_golden_model_1.n1918 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1918 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1918 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1918 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1918 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1918 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1918 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1993 , \oc8051_golden_model_1.n1994 [0]);
  buf(\oc8051_golden_model_1.n1994 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1994 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1994 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1994 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1994 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1994 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1994 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2010 , \oc8051_golden_model_1.n2011 [0]);
  buf(\oc8051_golden_model_1.n2011 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2011 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2011 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2011 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2011 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2027 , \oc8051_golden_model_1.n2028 [0]);
  buf(\oc8051_golden_model_1.n2028 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2028 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2028 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2028 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2028 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2028 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2028 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2044 , \oc8051_golden_model_1.n2045 [0]);
  buf(\oc8051_golden_model_1.n2045 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2045 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2045 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2045 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2045 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2045 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2045 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2049 , \oc8051_golden_model_1.n2053 [7]);
  buf(\oc8051_golden_model_1.n2050 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2050 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2050 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2050 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2050 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2050 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2050 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2051 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2051 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2051 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2051 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2051 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2051 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2051 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2051 [7], \oc8051_golden_model_1.n2053 [7]);
  buf(\oc8051_golden_model_1.n2052 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2052 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2052 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2052 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2052 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2052 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2052 [6], \oc8051_golden_model_1.n2053 [7]);
  buf(\oc8051_golden_model_1.n2053 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2053 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2053 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2053 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2053 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2053 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2053 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2068 , \oc8051_golden_model_1.n2069 [0]);
  buf(\oc8051_golden_model_1.n2069 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2069 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2069 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2069 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2069 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2069 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2069 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2097 , \oc8051_golden_model_1.n2100 [7]);
  buf(\oc8051_golden_model_1.n2098 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2098 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2098 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2098 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2098 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2098 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2098 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2098 [7], \oc8051_golden_model_1.n2100 [7]);
  buf(\oc8051_golden_model_1.n2099 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2099 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2099 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2099 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2099 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2099 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2099 [6], \oc8051_golden_model_1.n2100 [7]);
  buf(\oc8051_golden_model_1.n2100 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2107 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2107 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2107 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2107 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2108 , \oc8051_golden_model_1.n2126 [2]);
  buf(\oc8051_golden_model_1.n2109 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2109 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2109 [2], \oc8051_golden_model_1.n2126 [2]);
  buf(\oc8051_golden_model_1.n2109 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2109 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2109 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2109 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2109 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2110 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2110 [1], \oc8051_golden_model_1.n2126 [2]);
  buf(\oc8051_golden_model_1.n2110 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2110 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2110 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2110 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2110 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2125 , \oc8051_golden_model_1.n2126 [0]);
  buf(\oc8051_golden_model_1.n2126 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2126 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2126 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2126 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2126 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2126 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2301 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2304 , \oc8051_golden_model_1.n2330 [7]);
  buf(\oc8051_golden_model_1.n2306 , \oc8051_golden_model_1.n2330 [6]);
  buf(\oc8051_golden_model_1.n2312 , \oc8051_golden_model_1.n2330 [2]);
  buf(\oc8051_golden_model_1.n2313 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2313 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2313 [2], \oc8051_golden_model_1.n2330 [2]);
  buf(\oc8051_golden_model_1.n2313 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2313 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2313 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2313 [6], \oc8051_golden_model_1.n2330 [6]);
  buf(\oc8051_golden_model_1.n2313 [7], \oc8051_golden_model_1.n2330 [7]);
  buf(\oc8051_golden_model_1.n2314 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2314 [1], \oc8051_golden_model_1.n2330 [2]);
  buf(\oc8051_golden_model_1.n2314 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2314 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2314 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2314 [5], \oc8051_golden_model_1.n2330 [6]);
  buf(\oc8051_golden_model_1.n2314 [6], \oc8051_golden_model_1.n2330 [7]);
  buf(\oc8051_golden_model_1.n2329 , \oc8051_golden_model_1.n2330 [0]);
  buf(\oc8051_golden_model_1.n2330 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2330 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2330 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2330 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2334 , \oc8051_golden_model_1.n2360 [7]);
  buf(\oc8051_golden_model_1.n2336 , \oc8051_golden_model_1.n2360 [6]);
  buf(\oc8051_golden_model_1.n2342 , \oc8051_golden_model_1.n2360 [2]);
  buf(\oc8051_golden_model_1.n2343 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2343 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2343 [2], \oc8051_golden_model_1.n2360 [2]);
  buf(\oc8051_golden_model_1.n2343 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2343 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2343 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2343 [6], \oc8051_golden_model_1.n2360 [6]);
  buf(\oc8051_golden_model_1.n2343 [7], \oc8051_golden_model_1.n2360 [7]);
  buf(\oc8051_golden_model_1.n2344 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2344 [1], \oc8051_golden_model_1.n2360 [2]);
  buf(\oc8051_golden_model_1.n2344 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2344 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2344 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2344 [5], \oc8051_golden_model_1.n2360 [6]);
  buf(\oc8051_golden_model_1.n2344 [6], \oc8051_golden_model_1.n2360 [7]);
  buf(\oc8051_golden_model_1.n2359 , \oc8051_golden_model_1.n2360 [0]);
  buf(\oc8051_golden_model_1.n2360 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2360 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2360 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2360 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2364 , \oc8051_golden_model_1.n2390 [7]);
  buf(\oc8051_golden_model_1.n2366 , \oc8051_golden_model_1.n2390 [6]);
  buf(\oc8051_golden_model_1.n2372 , \oc8051_golden_model_1.n2390 [2]);
  buf(\oc8051_golden_model_1.n2373 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2373 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2373 [2], \oc8051_golden_model_1.n2390 [2]);
  buf(\oc8051_golden_model_1.n2373 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2373 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2373 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2373 [6], \oc8051_golden_model_1.n2390 [6]);
  buf(\oc8051_golden_model_1.n2373 [7], \oc8051_golden_model_1.n2390 [7]);
  buf(\oc8051_golden_model_1.n2374 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2374 [1], \oc8051_golden_model_1.n2390 [2]);
  buf(\oc8051_golden_model_1.n2374 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2374 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2374 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2374 [5], \oc8051_golden_model_1.n2390 [6]);
  buf(\oc8051_golden_model_1.n2374 [6], \oc8051_golden_model_1.n2390 [7]);
  buf(\oc8051_golden_model_1.n2389 , \oc8051_golden_model_1.n2390 [0]);
  buf(\oc8051_golden_model_1.n2390 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2390 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2390 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2390 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2394 , \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.n2396 , \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.n2402 , \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.n2403 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2403 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2403 [2], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.n2403 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2403 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2403 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2403 [6], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.n2403 [7], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.n2404 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2404 [1], \oc8051_golden_model_1.n2420 [2]);
  buf(\oc8051_golden_model_1.n2404 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2404 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2404 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2404 [5], \oc8051_golden_model_1.n2420 [6]);
  buf(\oc8051_golden_model_1.n2404 [6], \oc8051_golden_model_1.n2420 [7]);
  buf(\oc8051_golden_model_1.n2419 , \oc8051_golden_model_1.n2420 [0]);
  buf(\oc8051_golden_model_1.n2420 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2420 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2420 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2420 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2422 , \oc8051_golden_model_1.n2425 [7]);
  buf(\oc8051_golden_model_1.n2423 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2423 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2423 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2423 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2423 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2423 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2423 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2423 [7], \oc8051_golden_model_1.n2425 [7]);
  buf(\oc8051_golden_model_1.n2424 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2424 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2424 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2424 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2424 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2424 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2424 [6], \oc8051_golden_model_1.n2425 [7]);
  buf(\oc8051_golden_model_1.n2425 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2425 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2425 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2425 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2425 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2425 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2425 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2426 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2426 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2426 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2426 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2426 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2426 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2426 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2426 [7], \oc8051_golden_model_1.n2428 [7]);
  buf(\oc8051_golden_model_1.n2427 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2427 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2427 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2427 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2427 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2427 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2427 [6], \oc8051_golden_model_1.n2428 [7]);
  buf(\oc8051_golden_model_1.n2428 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2428 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2428 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2428 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2428 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2428 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2428 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2432 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2432 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2432 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2432 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2432 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2432 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2432 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2432 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2432 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2432 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2438 , \oc8051_golden_model_1.n2456 [2]);
  buf(\oc8051_golden_model_1.n2439 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2439 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2439 [2], \oc8051_golden_model_1.n2456 [2]);
  buf(\oc8051_golden_model_1.n2439 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2439 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2439 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2439 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2439 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2440 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2440 [1], \oc8051_golden_model_1.n2456 [2]);
  buf(\oc8051_golden_model_1.n2440 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2440 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2440 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2440 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2440 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2455 , \oc8051_golden_model_1.n2456 [0]);
  buf(\oc8051_golden_model_1.n2456 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2456 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2456 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2456 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2456 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2456 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2459 , \oc8051_golden_model_1.n2462 [7]);
  buf(\oc8051_golden_model_1.n2460 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2460 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2460 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2460 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2460 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2460 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2460 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2460 [7], \oc8051_golden_model_1.n2462 [7]);
  buf(\oc8051_golden_model_1.n2461 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2461 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2461 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2461 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2461 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2461 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2461 [6], \oc8051_golden_model_1.n2462 [7]);
  buf(\oc8051_golden_model_1.n2462 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2462 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2462 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2462 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2462 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2462 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2462 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2490 , \oc8051_golden_model_1.n2493 [7]);
  buf(\oc8051_golden_model_1.n2491 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2491 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2491 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2491 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2491 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2491 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2491 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2491 [7], \oc8051_golden_model_1.n2493 [7]);
  buf(\oc8051_golden_model_1.n2492 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2492 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2492 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2492 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2492 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2492 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2492 [6], \oc8051_golden_model_1.n2493 [7]);
  buf(\oc8051_golden_model_1.n2493 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2493 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2493 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2498 , \oc8051_golden_model_1.n2501 [7]);
  buf(\oc8051_golden_model_1.n2499 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2499 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2499 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2499 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2499 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2499 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2499 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2499 [7], \oc8051_golden_model_1.n2501 [7]);
  buf(\oc8051_golden_model_1.n2500 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2500 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2500 [6], \oc8051_golden_model_1.n2501 [7]);
  buf(\oc8051_golden_model_1.n2501 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2501 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2501 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2501 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2501 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2501 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2501 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2509 [7]);
  buf(\oc8051_golden_model_1.n2507 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2507 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2507 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2507 [7], \oc8051_golden_model_1.n2509 [7]);
  buf(\oc8051_golden_model_1.n2508 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2508 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2508 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2508 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2508 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2508 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2508 [6], \oc8051_golden_model_1.n2509 [7]);
  buf(\oc8051_golden_model_1.n2509 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2509 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2509 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2509 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2509 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2509 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2509 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2514 , \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2515 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2515 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2515 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2515 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2515 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2515 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2515 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2515 [7], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2516 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2516 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2516 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2516 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2516 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2516 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2516 [6], \oc8051_golden_model_1.n2517 [7]);
  buf(\oc8051_golden_model_1.n2517 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2517 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2517 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2517 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2517 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2517 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2517 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.n2523 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2523 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2523 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2523 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2523 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2523 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2523 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2523 [7], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.n2524 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2524 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2524 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2524 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2524 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2524 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2524 [6], \oc8051_golden_model_1.n2525 [7]);
  buf(\oc8051_golden_model_1.n2525 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2525 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2525 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2547 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2548 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2548 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2548 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2548 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2549 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2549 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2549 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2549 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2550 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2550 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2550 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2550 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2550 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2550 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2550 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2550 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2551 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2552 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2553 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2554 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2555 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2556 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2557 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2558 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2565 , \oc8051_golden_model_1.n2566 [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2575 [1], \oc8051_golden_model_1.n2751 [1]);
  buf(\oc8051_golden_model_1.n2575 [2], \oc8051_golden_model_1.n2751 [2]);
  buf(\oc8051_golden_model_1.n2575 [3], \oc8051_golden_model_1.n2751 [3]);
  buf(\oc8051_golden_model_1.n2575 [4], \oc8051_golden_model_1.n2751 [4]);
  buf(\oc8051_golden_model_1.n2575 [5], \oc8051_golden_model_1.n2751 [5]);
  buf(\oc8051_golden_model_1.n2575 [6], \oc8051_golden_model_1.n2751 [6]);
  buf(\oc8051_golden_model_1.n2575 [7], \oc8051_golden_model_1.n2751 [7]);
  buf(\oc8051_golden_model_1.n2576 [0], \oc8051_golden_model_1.n2751 [1]);
  buf(\oc8051_golden_model_1.n2576 [1], \oc8051_golden_model_1.n2751 [2]);
  buf(\oc8051_golden_model_1.n2576 [2], \oc8051_golden_model_1.n2751 [3]);
  buf(\oc8051_golden_model_1.n2576 [3], \oc8051_golden_model_1.n2751 [4]);
  buf(\oc8051_golden_model_1.n2576 [4], \oc8051_golden_model_1.n2751 [5]);
  buf(\oc8051_golden_model_1.n2576 [5], \oc8051_golden_model_1.n2751 [6]);
  buf(\oc8051_golden_model_1.n2576 [6], \oc8051_golden_model_1.n2751 [7]);
  buf(\oc8051_golden_model_1.n2591 , \oc8051_golden_model_1.n2733 [0]);
  buf(\oc8051_golden_model_1.n2592 [0], \oc8051_golden_model_1.n2733 [0]);
  buf(\oc8051_golden_model_1.n2592 [1], \oc8051_golden_model_1.n2751 [1]);
  buf(\oc8051_golden_model_1.n2592 [2], \oc8051_golden_model_1.n2751 [2]);
  buf(\oc8051_golden_model_1.n2592 [3], \oc8051_golden_model_1.n2751 [3]);
  buf(\oc8051_golden_model_1.n2592 [4], \oc8051_golden_model_1.n2751 [4]);
  buf(\oc8051_golden_model_1.n2592 [5], \oc8051_golden_model_1.n2751 [5]);
  buf(\oc8051_golden_model_1.n2592 [6], \oc8051_golden_model_1.n2751 [6]);
  buf(\oc8051_golden_model_1.n2592 [7], \oc8051_golden_model_1.n2751 [7]);
  buf(\oc8051_golden_model_1.n2593 , \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n2594 , \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n2596 , \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n2597 , \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n2598 , \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n2600 , \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n2607 , \oc8051_golden_model_1.n2608 [0]);
  buf(\oc8051_golden_model_1.n2608 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2608 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2608 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2608 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2608 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2608 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2608 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2623 , \oc8051_golden_model_1.n2624 [0]);
  buf(\oc8051_golden_model_1.n2624 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2624 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2624 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2624 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2624 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2624 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2624 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2653 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2654 [0], \oc8051_golden_model_1.n2751 [0]);
  buf(\oc8051_golden_model_1.n2654 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2654 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2654 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2654 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2654 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2654 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2654 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2673 , \oc8051_golden_model_1.n2691 [7]);
  buf(\oc8051_golden_model_1.n2674 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2674 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2674 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2674 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2674 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2674 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2674 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [7], \oc8051_golden_model_1.n2691 [7]);
  buf(\oc8051_golden_model_1.n2675 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2675 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2675 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2675 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2675 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2675 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2675 [6], \oc8051_golden_model_1.n2691 [7]);
  buf(\oc8051_golden_model_1.n2690 , \oc8051_golden_model_1.n2691 [0]);
  buf(\oc8051_golden_model_1.n2691 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2691 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2691 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2691 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2691 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2691 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.n2705 );
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.n2704 );
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.n2703 );
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.n2702 );
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2695 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2695 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.n2697 [4]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.n2697 [5]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.n2697 [6]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.n2697 [7]);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2698 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2712 , \oc8051_golden_model_1.n2713 [0]);
  buf(\oc8051_golden_model_1.n2713 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2713 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2713 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2713 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2713 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2713 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2713 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2731 , \oc8051_golden_model_1.n2732 [0]);
  buf(\oc8051_golden_model_1.n2732 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2732 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2732 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2732 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2732 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2732 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2732 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2733 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2733 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2733 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2733 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2733 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2733 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2733 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2749 , \oc8051_golden_model_1.n2750 [0]);
  buf(\oc8051_golden_model_1.n2750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2750 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm_next[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm_next[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm_next[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm_next[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm_next[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm_next[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm_next[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm_next[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm_next[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm_next[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm_next[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm_next[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm_next[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm_next[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm_next[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm_next[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm_next[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm_next[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm_next[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm_next[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm_next[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm_next[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm_next[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm_next[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm_next[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm_next[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm_next[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm_next[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm_next[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm_next[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm_next[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm_next[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm_next[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm_next[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm_next[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm_next[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm_next[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm_next[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm_next[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm_next[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm_next[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm_next[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm_next[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm_next[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm_next[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm_next[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm_next[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm_next[7], \oc8051_golden_model_1.TCON [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm_next[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm_next[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm_next[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm_next[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm_next[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm_next[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm_next[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm_next[7], \oc8051_golden_model_1.SCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm_next[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm_next[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm_next[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm_next[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm_next[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm_next[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm_next[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm_next[7], \oc8051_golden_model_1.SBUF [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm_next[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm_next[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm_next[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm_next[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm_next[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm_next[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm_next[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm_next[7], \oc8051_golden_model_1.PCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm_next[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm_next[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm_next[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm_next[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm_next[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm_next[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm_next[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm_next[7], \oc8051_golden_model_1.IP [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm_next[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm_next[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm_next[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm_next[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm_next[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm_next[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm_next[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm_next[7], \oc8051_golden_model_1.IE [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(PC_gm[0], \oc8051_golden_model_1.PC [0]);
  buf(PC_gm[1], \oc8051_golden_model_1.PC [1]);
  buf(PC_gm[2], \oc8051_golden_model_1.PC [2]);
  buf(PC_gm[3], \oc8051_golden_model_1.PC [3]);
  buf(PC_gm[4], \oc8051_golden_model_1.PC [4]);
  buf(PC_gm[5], \oc8051_golden_model_1.PC [5]);
  buf(PC_gm[6], \oc8051_golden_model_1.PC [6]);
  buf(PC_gm[7], \oc8051_golden_model_1.PC [7]);
  buf(PC_gm[8], \oc8051_golden_model_1.PC [8]);
  buf(PC_gm[9], \oc8051_golden_model_1.PC [9]);
  buf(PC_gm[10], \oc8051_golden_model_1.PC [10]);
  buf(PC_gm[11], \oc8051_golden_model_1.PC [11]);
  buf(PC_gm[12], \oc8051_golden_model_1.PC [12]);
  buf(PC_gm[13], \oc8051_golden_model_1.PC [13]);
  buf(PC_gm[14], \oc8051_golden_model_1.PC [14]);
  buf(PC_gm[15], \oc8051_golden_model_1.PC [15]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc_impl[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc_impl[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc_impl[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc_impl[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc_impl[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc_impl[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc_impl[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc_impl[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc_impl[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc_impl[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc_impl[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc_impl[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc_impl[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc_impl[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc_impl[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc_impl[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(property_invalid_dec_rom_pc, 1'b0);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
