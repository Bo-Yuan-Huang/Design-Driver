
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire _44007_;
  wire _44008_;
  wire _44009_;
  wire _44010_;
  wire _44011_;
  wire _44012_;
  wire _44013_;
  wire _44014_;
  wire _44015_;
  wire _44016_;
  wire _44017_;
  wire _44018_;
  wire _44019_;
  wire _44020_;
  wire _44021_;
  wire _44022_;
  wire _44023_;
  wire _44024_;
  wire _44025_;
  wire _44026_;
  wire _44027_;
  wire _44028_;
  wire _44029_;
  wire _44030_;
  wire _44031_;
  wire _44032_;
  wire _44033_;
  wire _44034_;
  wire _44035_;
  wire _44036_;
  wire _44037_;
  wire _44038_;
  wire _44039_;
  wire _44040_;
  wire _44041_;
  wire _44042_;
  wire _44043_;
  wire _44044_;
  wire _44045_;
  wire _44046_;
  wire _44047_;
  wire _44048_;
  wire _44049_;
  wire _44050_;
  wire _44051_;
  wire _44052_;
  wire _44053_;
  wire _44054_;
  wire _44055_;
  wire _44056_;
  wire _44057_;
  wire _44058_;
  wire _44059_;
  wire _44060_;
  wire _44061_;
  wire _44062_;
  wire _44063_;
  wire _44064_;
  wire _44065_;
  wire _44066_;
  wire _44067_;
  wire _44068_;
  wire _44069_;
  wire _44070_;
  wire _44071_;
  wire _44072_;
  wire _44073_;
  wire _44074_;
  wire _44075_;
  wire _44076_;
  wire _44077_;
  wire _44078_;
  wire _44079_;
  wire _44080_;
  wire _44081_;
  wire _44082_;
  wire _44083_;
  wire _44084_;
  wire _44085_;
  wire _44086_;
  wire _44087_;
  wire _44088_;
  wire _44089_;
  wire _44090_;
  wire _44091_;
  wire _44092_;
  wire _44093_;
  wire _44094_;
  wire _44095_;
  wire _44096_;
  wire _44097_;
  wire _44098_;
  wire _44099_;
  wire _44100_;
  wire _44101_;
  wire _44102_;
  wire _44103_;
  wire _44104_;
  wire _44105_;
  wire _44106_;
  wire _44107_;
  wire _44108_;
  wire _44109_;
  wire _44110_;
  wire _44111_;
  wire _44112_;
  wire _44113_;
  wire _44114_;
  wire _44115_;
  wire _44116_;
  wire _44117_;
  wire _44118_;
  wire _44119_;
  wire _44120_;
  wire _44121_;
  wire _44122_;
  wire _44123_;
  wire _44124_;
  wire _44125_;
  wire _44126_;
  wire _44127_;
  wire _44128_;
  wire _44129_;
  wire _44130_;
  wire _44131_;
  wire _44132_;
  wire _44133_;
  wire _44134_;
  wire _44135_;
  wire _44136_;
  wire _44137_;
  wire _44138_;
  wire _44139_;
  wire _44140_;
  wire _44141_;
  wire _44142_;
  wire _44143_;
  wire _44144_;
  wire _44145_;
  wire _44146_;
  wire _44147_;
  wire _44148_;
  wire _44149_;
  wire _44150_;
  wire _44151_;
  wire _44152_;
  wire _44153_;
  wire _44154_;
  wire _44155_;
  wire _44156_;
  wire _44157_;
  wire _44158_;
  wire _44159_;
  wire _44160_;
  wire _44161_;
  wire _44162_;
  wire _44163_;
  wire _44164_;
  wire _44165_;
  wire _44166_;
  wire _44167_;
  wire _44168_;
  wire _44169_;
  wire _44170_;
  wire _44171_;
  wire _44172_;
  wire _44173_;
  wire _44174_;
  wire _44175_;
  wire _44176_;
  wire _44177_;
  wire _44178_;
  wire _44179_;
  wire _44180_;
  wire _44181_;
  wire _44182_;
  wire _44183_;
  wire _44184_;
  wire _44185_;
  wire _44186_;
  wire _44187_;
  wire _44188_;
  wire _44189_;
  wire _44190_;
  wire _44191_;
  wire _44192_;
  wire _44193_;
  wire _44194_;
  wire _44195_;
  wire _44196_;
  wire _44197_;
  wire _44198_;
  wire _44199_;
  wire _44200_;
  wire _44201_;
  wire _44202_;
  wire _44203_;
  wire _44204_;
  wire _44205_;
  wire _44206_;
  wire _44207_;
  wire _44208_;
  wire _44209_;
  wire _44210_;
  wire _44211_;
  wire _44212_;
  wire _44213_;
  wire _44214_;
  wire _44215_;
  wire _44216_;
  wire _44217_;
  wire _44218_;
  wire _44219_;
  wire _44220_;
  wire _44221_;
  wire _44222_;
  wire _44223_;
  wire _44224_;
  wire _44225_;
  wire _44226_;
  wire _44227_;
  wire _44228_;
  wire _44229_;
  wire _44230_;
  wire _44231_;
  wire _44232_;
  wire _44233_;
  wire _44234_;
  wire _44235_;
  wire _44236_;
  wire _44237_;
  wire _44238_;
  wire _44239_;
  wire _44240_;
  wire _44241_;
  wire _44242_;
  wire _44243_;
  wire _44244_;
  wire _44245_;
  wire _44246_;
  wire _44247_;
  wire _44248_;
  wire _44249_;
  wire _44250_;
  wire _44251_;
  wire _44252_;
  wire _44253_;
  wire _44254_;
  wire _44255_;
  wire _44256_;
  wire _44257_;
  wire _44258_;
  wire _44259_;
  wire _44260_;
  wire _44261_;
  wire _44262_;
  wire _44263_;
  wire _44264_;
  wire _44265_;
  wire _44266_;
  wire _44267_;
  wire _44268_;
  wire _44269_;
  wire _44270_;
  wire _44271_;
  wire _44272_;
  wire _44273_;
  wire _44274_;
  wire _44275_;
  wire _44276_;
  wire _44277_;
  wire _44278_;
  wire _44279_;
  wire _44280_;
  wire _44281_;
  wire _44282_;
  wire _44283_;
  wire _44284_;
  wire _44285_;
  wire _44286_;
  wire _44287_;
  wire _44288_;
  wire _44289_;
  wire _44290_;
  wire _44291_;
  wire _44292_;
  wire _44293_;
  wire _44294_;
  wire _44295_;
  wire _44296_;
  wire _44297_;
  wire _44298_;
  wire _44299_;
  wire _44300_;
  wire _44301_;
  wire _44302_;
  wire _44303_;
  wire _44304_;
  wire _44305_;
  wire _44306_;
  wire _44307_;
  wire _44308_;
  wire _44309_;
  wire _44310_;
  wire _44311_;
  wire _44312_;
  wire _44313_;
  wire _44314_;
  wire _44315_;
  wire _44316_;
  wire _44317_;
  wire _44318_;
  wire _44319_;
  wire _44320_;
  wire _44321_;
  wire _44322_;
  wire _44323_;
  wire _44324_;
  wire _44325_;
  wire _44326_;
  wire _44327_;
  wire _44328_;
  wire _44329_;
  wire _44330_;
  wire _44331_;
  wire _44332_;
  wire _44333_;
  wire _44334_;
  wire _44335_;
  wire _44336_;
  wire _44337_;
  wire _44338_;
  wire _44339_;
  wire _44340_;
  wire _44341_;
  wire _44342_;
  wire _44343_;
  wire _44344_;
  wire _44345_;
  wire _44346_;
  wire _44347_;
  wire _44348_;
  wire _44349_;
  wire _44350_;
  wire _44351_;
  wire _44352_;
  wire _44353_;
  wire _44354_;
  wire _44355_;
  wire _44356_;
  wire _44357_;
  wire _44358_;
  wire _44359_;
  wire _44360_;
  wire _44361_;
  wire _44362_;
  wire _44363_;
  wire _44364_;
  wire _44365_;
  wire _44366_;
  wire _44367_;
  wire _44368_;
  wire _44369_;
  wire _44370_;
  wire _44371_;
  wire _44372_;
  wire _44373_;
  wire _44374_;
  wire _44375_;
  wire _44376_;
  wire _44377_;
  wire _44378_;
  wire _44379_;
  wire _44380_;
  wire _44381_;
  wire _44382_;
  wire _44383_;
  wire _44384_;
  wire _44385_;
  wire _44386_;
  wire _44387_;
  wire _44388_;
  wire _44389_;
  wire _44390_;
  wire _44391_;
  wire _44392_;
  wire _44393_;
  wire _44394_;
  wire _44395_;
  wire _44396_;
  wire _44397_;
  wire _44398_;
  wire _44399_;
  wire _44400_;
  wire _44401_;
  wire _44402_;
  wire _44403_;
  wire _44404_;
  wire _44405_;
  wire _44406_;
  wire _44407_;
  wire _44408_;
  wire _44409_;
  wire _44410_;
  wire _44411_;
  wire _44412_;
  wire _44413_;
  wire _44414_;
  wire _44415_;
  wire _44416_;
  wire _44417_;
  wire _44418_;
  wire _44419_;
  wire _44420_;
  wire _44421_;
  wire _44422_;
  wire _44423_;
  wire _44424_;
  wire _44425_;
  wire _44426_;
  wire _44427_;
  wire _44428_;
  wire _44429_;
  wire _44430_;
  wire _44431_;
  wire _44432_;
  wire _44433_;
  wire _44434_;
  wire _44435_;
  wire _44436_;
  wire _44437_;
  wire _44438_;
  wire _44439_;
  wire _44440_;
  wire _44441_;
  wire _44442_;
  wire _44443_;
  wire _44444_;
  wire _44445_;
  wire _44446_;
  wire _44447_;
  wire _44448_;
  wire _44449_;
  wire _44450_;
  wire _44451_;
  wire _44452_;
  wire _44453_;
  wire _44454_;
  wire _44455_;
  wire _44456_;
  wire _44457_;
  wire _44458_;
  wire _44459_;
  wire _44460_;
  wire _44461_;
  wire _44462_;
  wire _44463_;
  wire _44464_;
  wire _44465_;
  wire _44466_;
  wire _44467_;
  wire _44468_;
  wire _44469_;
  wire _44470_;
  wire _44471_;
  wire _44472_;
  wire _44473_;
  wire _44474_;
  wire _44475_;
  wire _44476_;
  wire _44477_;
  wire _44478_;
  wire _44479_;
  wire _44480_;
  wire _44481_;
  wire _44482_;
  wire _44483_;
  wire _44484_;
  wire _44485_;
  wire _44486_;
  wire _44487_;
  wire _44488_;
  wire _44489_;
  wire _44490_;
  wire _44491_;
  wire _44492_;
  wire _44493_;
  wire _44494_;
  wire _44495_;
  wire _44496_;
  wire _44497_;
  wire _44498_;
  wire _44499_;
  wire _44500_;
  wire _44501_;
  wire _44502_;
  wire _44503_;
  wire _44504_;
  wire _44505_;
  wire _44506_;
  wire _44507_;
  wire _44508_;
  wire _44509_;
  wire _44510_;
  wire _44511_;
  wire _44512_;
  wire _44513_;
  wire _44514_;
  wire _44515_;
  wire _44516_;
  wire _44517_;
  wire _44518_;
  wire _44519_;
  wire _44520_;
  wire _44521_;
  wire _44522_;
  wire _44523_;
  wire _44524_;
  wire _44525_;
  wire _44526_;
  wire _44527_;
  wire _44528_;
  wire _44529_;
  wire _44530_;
  wire _44531_;
  wire _44532_;
  wire _44533_;
  wire _44534_;
  wire _44535_;
  wire _44536_;
  wire _44537_;
  wire _44538_;
  wire _44539_;
  wire _44540_;
  wire _44541_;
  wire _44542_;
  wire _44543_;
  wire _44544_;
  wire _44545_;
  wire _44546_;
  wire _44547_;
  wire _44548_;
  wire _44549_;
  wire _44550_;
  wire _44551_;
  wire _44552_;
  wire _44553_;
  wire _44554_;
  wire _44555_;
  wire _44556_;
  wire _44557_;
  wire _44558_;
  wire _44559_;
  wire _44560_;
  wire _44561_;
  wire _44562_;
  wire _44563_;
  wire _44564_;
  wire _44565_;
  wire _44566_;
  wire _44567_;
  wire _44568_;
  wire _44569_;
  wire _44570_;
  wire _44571_;
  wire _44572_;
  wire _44573_;
  wire _44574_;
  wire _44575_;
  wire _44576_;
  wire _44577_;
  wire _44578_;
  wire _44579_;
  wire _44580_;
  wire _44581_;
  wire _44582_;
  wire _44583_;
  wire _44584_;
  wire _44585_;
  wire _44586_;
  wire _44587_;
  wire _44588_;
  wire _44589_;
  wire _44590_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1090 ;
  wire [3:0] \oc8051_golden_model_1.n1092 ;
  wire [3:0] \oc8051_golden_model_1.n1094 ;
  wire [3:0] \oc8051_golden_model_1.n1095 ;
  wire [3:0] \oc8051_golden_model_1.n1096 ;
  wire [3:0] \oc8051_golden_model_1.n1097 ;
  wire [3:0] \oc8051_golden_model_1.n1098 ;
  wire [3:0] \oc8051_golden_model_1.n1099 ;
  wire [3:0] \oc8051_golden_model_1.n1100 ;
  wire \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1175 ;
  wire [8:0] \oc8051_golden_model_1.n1176 ;
  wire [8:0] \oc8051_golden_model_1.n1177 ;
  wire [7:0] \oc8051_golden_model_1.n1178 ;
  wire \oc8051_golden_model_1.n1179 ;
  wire \oc8051_golden_model_1.n1180 ;
  wire [2:0] \oc8051_golden_model_1.n1181 ;
  wire \oc8051_golden_model_1.n1182 ;
  wire [1:0] \oc8051_golden_model_1.n1183 ;
  wire [7:0] \oc8051_golden_model_1.n1184 ;
  wire [15:0] \oc8051_golden_model_1.n1211 ;
  wire [7:0] \oc8051_golden_model_1.n1213 ;
  wire [8:0] \oc8051_golden_model_1.n1215 ;
  wire [8:0] \oc8051_golden_model_1.n1219 ;
  wire \oc8051_golden_model_1.n1220 ;
  wire [3:0] \oc8051_golden_model_1.n1221 ;
  wire [4:0] \oc8051_golden_model_1.n1222 ;
  wire [4:0] \oc8051_golden_model_1.n1226 ;
  wire \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1228 ;
  wire \oc8051_golden_model_1.n1236 ;
  wire [7:0] \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire \oc8051_golden_model_1.n1242 ;
  wire [4:0] \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire [7:0] \oc8051_golden_model_1.n1257 ;
  wire [8:0] \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire \oc8051_golden_model_1.n1262 ;
  wire [3:0] \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [8:0] \oc8051_golden_model_1.n1279 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire \oc8051_golden_model_1.n1287 ;
  wire [7:0] \oc8051_golden_model_1.n1288 ;
  wire [8:0] \oc8051_golden_model_1.n1290 ;
  wire [8:0] \oc8051_golden_model_1.n1292 ;
  wire \oc8051_golden_model_1.n1293 ;
  wire [4:0] \oc8051_golden_model_1.n1294 ;
  wire [4:0] \oc8051_golden_model_1.n1296 ;
  wire \oc8051_golden_model_1.n1297 ;
  wire [8:0] \oc8051_golden_model_1.n1298 ;
  wire \oc8051_golden_model_1.n1305 ;
  wire [7:0] \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1308 ;
  wire \oc8051_golden_model_1.n1309 ;
  wire [7:0] \oc8051_golden_model_1.n1310 ;
  wire [8:0] \oc8051_golden_model_1.n1312 ;
  wire \oc8051_golden_model_1.n1313 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire [7:0] \oc8051_golden_model_1.n1321 ;
  wire [7:0] \oc8051_golden_model_1.n1322 ;
  wire [8:0] \oc8051_golden_model_1.n1325 ;
  wire [8:0] \oc8051_golden_model_1.n1326 ;
  wire [7:0] \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire [7:0] \oc8051_golden_model_1.n1329 ;
  wire [7:0] \oc8051_golden_model_1.n1330 ;
  wire [8:0] \oc8051_golden_model_1.n1333 ;
  wire [8:0] \oc8051_golden_model_1.n1335 ;
  wire \oc8051_golden_model_1.n1336 ;
  wire [4:0] \oc8051_golden_model_1.n1337 ;
  wire [4:0] \oc8051_golden_model_1.n1339 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire [7:0] \oc8051_golden_model_1.n1348 ;
  wire [8:0] \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire [4:0] \oc8051_golden_model_1.n1355 ;
  wire \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1363 ;
  wire [7:0] \oc8051_golden_model_1.n1364 ;
  wire [8:0] \oc8051_golden_model_1.n1368 ;
  wire \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1371 ;
  wire \oc8051_golden_model_1.n1372 ;
  wire \oc8051_golden_model_1.n1379 ;
  wire [7:0] \oc8051_golden_model_1.n1380 ;
  wire [8:0] \oc8051_golden_model_1.n1384 ;
  wire \oc8051_golden_model_1.n1385 ;
  wire [4:0] \oc8051_golden_model_1.n1387 ;
  wire \oc8051_golden_model_1.n1388 ;
  wire \oc8051_golden_model_1.n1395 ;
  wire [7:0] \oc8051_golden_model_1.n1396 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire [6:0] \oc8051_golden_model_1.n1557 ;
  wire [7:0] \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1581 ;
  wire [7:0] \oc8051_golden_model_1.n1582 ;
  wire [3:0] \oc8051_golden_model_1.n1589 ;
  wire \oc8051_golden_model_1.n1590 ;
  wire [7:0] \oc8051_golden_model_1.n1591 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire \oc8051_golden_model_1.n1738 ;
  wire \oc8051_golden_model_1.n1740 ;
  wire \oc8051_golden_model_1.n1746 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire \oc8051_golden_model_1.n1751 ;
  wire \oc8051_golden_model_1.n1753 ;
  wire \oc8051_golden_model_1.n1759 ;
  wire [7:0] \oc8051_golden_model_1.n1760 ;
  wire \oc8051_golden_model_1.n1764 ;
  wire \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1772 ;
  wire [7:0] \oc8051_golden_model_1.n1773 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire \oc8051_golden_model_1.n1779 ;
  wire \oc8051_golden_model_1.n1785 ;
  wire [7:0] \oc8051_golden_model_1.n1786 ;
  wire \oc8051_golden_model_1.n1788 ;
  wire [7:0] \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [15:0] \oc8051_golden_model_1.n1794 ;
  wire \oc8051_golden_model_1.n1800 ;
  wire [7:0] \oc8051_golden_model_1.n1801 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1825 ;
  wire [7:0] \oc8051_golden_model_1.n1826 ;
  wire \oc8051_golden_model_1.n1831 ;
  wire [7:0] \oc8051_golden_model_1.n1832 ;
  wire \oc8051_golden_model_1.n1837 ;
  wire [7:0] \oc8051_golden_model_1.n1838 ;
  wire \oc8051_golden_model_1.n1843 ;
  wire [7:0] \oc8051_golden_model_1.n1844 ;
  wire \oc8051_golden_model_1.n1849 ;
  wire [7:0] \oc8051_golden_model_1.n1850 ;
  wire [7:0] \oc8051_golden_model_1.n1851 ;
  wire [3:0] \oc8051_golden_model_1.n1852 ;
  wire [7:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1889 ;
  wire \oc8051_golden_model_1.n1908 ;
  wire [7:0] \oc8051_golden_model_1.n1909 ;
  wire [7:0] \oc8051_golden_model_1.n1913 ;
  wire [3:0] \oc8051_golden_model_1.n1914 ;
  wire [7:0] \oc8051_golden_model_1.n1915 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _44591_ (_43634_, rst);
  not _44592_ (_19448_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _44593_ (_19459_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44594_ (_19470_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _19459_);
  and _44595_ (_19481_, _19470_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44596_ (_19492_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _19459_);
  and _44597_ (_19503_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _19459_);
  nor _44598_ (_19514_, _19503_, _19492_);
  and _44599_ (_19525_, _19514_, _19481_);
  nor _44600_ (_19536_, _19525_, _19448_);
  and _44601_ (_19547_, _19448_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44602_ (_19558_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _44603_ (_19569_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _19558_);
  nor _44604_ (_19579_, _19569_, _19547_);
  not _44605_ (_19590_, _19579_);
  and _44606_ (_19601_, _19590_, _19525_);
  or _44607_ (_19612_, _19601_, _19536_);
  and _44608_ (_22076_, _19612_, _43634_);
  nor _44609_ (_19633_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44610_ (_19644_, _19633_);
  and _44611_ (_19654_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _44612_ (_19665_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _44613_ (_19676_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _44614_ (_19687_, _19676_);
  not _44615_ (_19698_, _19569_);
  nor _44616_ (_19720_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _44617_ (_19732_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _44618_ (_19743_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _19732_);
  nor _44619_ (_19755_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _44620_ (_19767_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _44621_ (_19779_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _19767_);
  nor _44622_ (_19791_, _19779_, _19755_);
  nor _44623_ (_19792_, _19791_, _19743_);
  not _44624_ (_19803_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _44625_ (_19814_, _19743_, _19803_);
  nor _44626_ (_19825_, _19814_, _19792_);
  and _44627_ (_19835_, _19825_, _19720_);
  not _44628_ (_19846_, _19835_);
  and _44629_ (_19857_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44630_ (_19868_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _44631_ (_19879_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44632_ (_19890_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _19879_);
  and _44633_ (_19901_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _44634_ (_19912_, _19901_, _19868_);
  and _44635_ (_19922_, _19912_, _19846_);
  nor _44636_ (_19933_, _19922_, _19698_);
  not _44637_ (_19944_, _19547_);
  nor _44638_ (_19955_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _44639_ (_19966_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _19767_);
  nor _44640_ (_19977_, _19966_, _19955_);
  nor _44641_ (_19988_, _19977_, _19743_);
  not _44642_ (_19999_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _44643_ (_20009_, _19743_, _19999_);
  nor _44644_ (_20020_, _20009_, _19988_);
  and _44645_ (_20031_, _20020_, _19720_);
  not _44646_ (_20042_, _20031_);
  and _44647_ (_20053_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _44648_ (_20064_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _44649_ (_20075_, _20064_, _20053_);
  and _44650_ (_20085_, _20075_, _20042_);
  nor _44651_ (_20096_, _20085_, _19944_);
  nor _44652_ (_20107_, _20096_, _19933_);
  nor _44653_ (_20118_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _44654_ (_20129_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _19767_);
  nor _44655_ (_20140_, _20129_, _20118_);
  nor _44656_ (_20151_, _20140_, _19743_);
  not _44657_ (_20162_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _44658_ (_20172_, _19743_, _20162_);
  nor _44659_ (_20183_, _20172_, _20151_);
  and _44660_ (_20194_, _20183_, _19720_);
  not _44661_ (_20205_, _20194_);
  and _44662_ (_20216_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _44663_ (_20227_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44664_ (_20238_, _20227_, _20216_);
  and _44665_ (_20248_, _20238_, _20205_);
  nor _44666_ (_20259_, _20248_, _19590_);
  nor _44667_ (_20270_, _20259_, _19633_);
  and _44668_ (_20281_, _20270_, _20107_);
  nor _44669_ (_20292_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _44670_ (_20303_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _19767_);
  nor _44671_ (_20314_, _20303_, _20292_);
  nor _44672_ (_20325_, _20314_, _19743_);
  not _44673_ (_20335_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _44674_ (_20346_, _19743_, _20335_);
  nor _44675_ (_20357_, _20346_, _20325_);
  and _44676_ (_20368_, _20357_, _19720_);
  not _44677_ (_20379_, _20368_);
  and _44678_ (_20390_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _44679_ (_20401_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _44680_ (_20412_, _20401_, _20390_);
  and _44681_ (_20422_, _20412_, _20379_);
  and _44682_ (_20433_, _20422_, _19633_);
  nor _44683_ (_20444_, _20433_, _20281_);
  not _44684_ (_20455_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44685_ (_20466_, _20455_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44686_ (_20477_, _20466_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44687_ (_20488_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _44688_ (_20499_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44689_ (_20509_, _20499_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44690_ (_20520_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _44691_ (_20531_, _20520_, _20488_);
  nor _44692_ (_20542_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44693_ (_20553_, _20542_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44694_ (_20564_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _44695_ (_20575_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44696_ (_20586_, _20466_, _20575_);
  and _44697_ (_20596_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _44698_ (_20607_, _20596_, _20564_);
  and _44699_ (_20618_, _20607_, _20531_);
  and _44700_ (_20639_, _20542_, _20455_);
  and _44701_ (_20640_, _20639_, _20357_);
  and _44702_ (_20651_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44703_ (_20662_, _20651_, _20575_);
  and _44704_ (_20682_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _44705_ (_20683_, _20651_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44706_ (_20694_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _44707_ (_20715_, _20694_, _20682_);
  not _44708_ (_20716_, _20715_);
  nor _44709_ (_20727_, _20716_, _20640_);
  and _44710_ (_20738_, _20727_, _20618_);
  not _44711_ (_20749_, _20738_);
  and _44712_ (_20769_, _20749_, _20444_);
  not _44713_ (_20770_, _20769_);
  nor _44714_ (_20781_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _44715_ (_20792_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _19767_);
  nor _44716_ (_20803_, _20792_, _20781_);
  nor _44717_ (_20814_, _20803_, _19743_);
  not _44718_ (_20825_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _44719_ (_20836_, _19743_, _20825_);
  nor _44720_ (_20846_, _20836_, _20814_);
  and _44721_ (_20857_, _20846_, _19720_);
  not _44722_ (_20868_, _20857_);
  and _44723_ (_20879_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _44724_ (_20900_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44725_ (_20901_, _20900_, _20879_);
  and _44726_ (_20912_, _20901_, _20868_);
  nor _44727_ (_20923_, _20912_, _19698_);
  nor _44728_ (_20934_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _44729_ (_20944_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _19767_);
  nor _44730_ (_20955_, _20944_, _20934_);
  nor _44731_ (_20966_, _20955_, _19743_);
  not _44732_ (_20977_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _44733_ (_20988_, _19743_, _20977_);
  nor _44734_ (_20999_, _20988_, _20966_);
  and _44735_ (_21010_, _20999_, _19720_);
  not _44736_ (_21021_, _21010_);
  and _44737_ (_21032_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _44738_ (_21042_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44739_ (_21053_, _21042_, _21032_);
  and _44740_ (_21074_, _21053_, _21021_);
  nor _44741_ (_21075_, _21074_, _19944_);
  nor _44742_ (_21086_, _21075_, _20923_);
  nor _44743_ (_21097_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _44744_ (_21108_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _19767_);
  nor _44745_ (_21119_, _21108_, _21097_);
  nor _44746_ (_21129_, _21119_, _19743_);
  not _44747_ (_21140_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _44748_ (_21151_, _19743_, _21140_);
  nor _44749_ (_21162_, _21151_, _21129_);
  and _44750_ (_21173_, _21162_, _19720_);
  not _44751_ (_21184_, _21173_);
  and _44752_ (_21195_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _44753_ (_21206_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44754_ (_21217_, _21206_, _21195_);
  and _44755_ (_21227_, _21217_, _21184_);
  nor _44756_ (_21238_, _21227_, _19590_);
  nor _44757_ (_21249_, _21238_, _19633_);
  and _44758_ (_21270_, _21249_, _21086_);
  nor _44759_ (_21271_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _44760_ (_21282_, _19767_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _44761_ (_21293_, _21282_, _21271_);
  nor _44762_ (_21304_, _21293_, _19743_);
  not _44763_ (_21314_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _44764_ (_21325_, _19743_, _21314_);
  nor _44765_ (_21336_, _21325_, _21304_);
  and _44766_ (_21347_, _21336_, _19720_);
  not _44767_ (_21358_, _21347_);
  and _44768_ (_21369_, _19857_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44769_ (_21380_, _19890_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _44770_ (_21391_, _21380_, _21369_);
  and _44771_ (_21402_, _21391_, _21358_);
  and _44772_ (_21412_, _21402_, _19633_);
  nor _44773_ (_21423_, _21412_, _21270_);
  and _44774_ (_21434_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _44775_ (_21445_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _44776_ (_21456_, _21445_, _21434_);
  and _44777_ (_21467_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _44778_ (_21478_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor _44779_ (_21489_, _21478_, _21467_);
  and _44780_ (_21499_, _21489_, _21456_);
  and _44781_ (_21510_, _21336_, _20639_);
  and _44782_ (_21521_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _44783_ (_21532_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _44784_ (_21543_, _21532_, _21521_);
  not _44785_ (_21554_, _21543_);
  nor _44786_ (_21565_, _21554_, _21510_);
  and _44787_ (_21576_, _21565_, _21499_);
  not _44788_ (_21587_, _21576_);
  and _44789_ (_21597_, _21587_, _21423_);
  and _44790_ (_21618_, _21597_, _20770_);
  and _44791_ (_21619_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _44792_ (_21630_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _44793_ (_21641_, _21630_, _21619_);
  and _44794_ (_21652_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _44795_ (_21663_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _44796_ (_21674_, _21663_, _21652_);
  and _44797_ (_21684_, _21674_, _21641_);
  and _44798_ (_21695_, _20999_, _20639_);
  and _44799_ (_21706_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _44800_ (_21727_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44801_ (_21728_, _21727_, _21706_);
  not _44802_ (_21739_, _21728_);
  nor _44803_ (_21750_, _21739_, _21695_);
  and _44804_ (_21761_, _21750_, _21684_);
  not _44805_ (_21772_, _21761_);
  and _44806_ (_21782_, _21772_, _21423_);
  not _44807_ (_21793_, _21782_);
  and _44808_ (_21804_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _44809_ (_21815_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _44810_ (_21826_, _21815_, _21804_);
  and _44811_ (_21837_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _44812_ (_21848_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _44813_ (_21859_, _21848_, _21837_);
  and _44814_ (_21870_, _21859_, _21826_);
  and _44815_ (_21880_, _20639_, _20020_);
  and _44816_ (_21891_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _44817_ (_21902_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _44818_ (_21913_, _21902_, _21891_);
  not _44819_ (_21924_, _21913_);
  nor _44820_ (_21935_, _21924_, _21880_);
  and _44821_ (_21946_, _21935_, _21870_);
  not _44822_ (_21957_, _21946_);
  and _44823_ (_21967_, _21957_, _20444_);
  and _44824_ (_21978_, _21782_, _21967_);
  nor _44825_ (_21989_, _20769_, _21978_);
  nor _44826_ (_22000_, _21989_, _21793_);
  and _44827_ (_22011_, _21597_, _20769_);
  and _44828_ (_22022_, _20749_, _21423_);
  and _44829_ (_22033_, _21587_, _20444_);
  nor _44830_ (_22044_, _22033_, _22022_);
  nor _44831_ (_22055_, _22044_, _22011_);
  and _44832_ (_22065_, _22055_, _22000_);
  and _44833_ (_22077_, _22065_, _21618_);
  and _44834_ (_22088_, _21423_, _21957_);
  and _44835_ (_22099_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _44836_ (_22110_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nor _44837_ (_22121_, _22110_, _22099_);
  and _44838_ (_22132_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _44839_ (_22142_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _44840_ (_22153_, _22142_, _22132_);
  and _44841_ (_22174_, _22153_, _22121_);
  and _44842_ (_22175_, _20846_, _20639_);
  and _44843_ (_22186_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _44844_ (_22197_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44845_ (_22208_, _22197_, _22186_);
  not _44846_ (_22219_, _22208_);
  nor _44847_ (_22229_, _22219_, _22175_);
  and _44848_ (_22240_, _22229_, _22174_);
  not _44849_ (_22251_, _22240_);
  and _44850_ (_22262_, _22251_, _20444_);
  and _44851_ (_22273_, _22262_, _22088_);
  and _44852_ (_22284_, _21772_, _20444_);
  nor _44853_ (_22295_, _22284_, _22088_);
  nor _44854_ (_22306_, _22295_, _21978_);
  and _44855_ (_22316_, _22306_, _22273_);
  and _44856_ (_22327_, _20749_, _21978_);
  not _44857_ (_22338_, _22327_);
  and _44858_ (_22349_, _22000_, _22338_);
  nor _44859_ (_22360_, _20769_, _21782_);
  nor _44860_ (_22371_, _22360_, _22349_);
  and _44861_ (_22382_, _22371_, _22316_);
  not _44862_ (_22393_, _22055_);
  nor _44863_ (_22403_, _22393_, _22000_);
  and _44864_ (_22414_, _22393_, _22000_);
  nor _44865_ (_22425_, _22414_, _22403_);
  not _44866_ (_22436_, _22425_);
  and _44867_ (_22447_, _22436_, _22382_);
  nor _44868_ (_22468_, _22436_, _22382_);
  nor _44869_ (_22469_, _22468_, _22447_);
  not _44870_ (_22480_, _22469_);
  and _44871_ (_22490_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _44872_ (_22501_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _44873_ (_22512_, _22501_, _22490_);
  and _44874_ (_22523_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _44875_ (_22534_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _44876_ (_22545_, _22534_, _22523_);
  and _44877_ (_22556_, _22545_, _22512_);
  and _44878_ (_22576_, _21162_, _20639_);
  and _44879_ (_22577_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _44880_ (_22588_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44881_ (_22599_, _22588_, _22577_);
  not _44882_ (_22610_, _22599_);
  nor _44883_ (_22621_, _22610_, _22576_);
  and _44884_ (_22632_, _22621_, _22556_);
  not _44885_ (_22643_, _22632_);
  and _44886_ (_22653_, _22643_, _21423_);
  and _44887_ (_22664_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _44888_ (_22675_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _44889_ (_22686_, _22675_, _22664_);
  and _44890_ (_22697_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _44891_ (_22708_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _44892_ (_22719_, _22708_, _22697_);
  and _44893_ (_22729_, _22719_, _22686_);
  and _44894_ (_22740_, _20639_, _19825_);
  and _44895_ (_22751_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and _44896_ (_22762_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _44897_ (_22773_, _22762_, _22751_);
  not _44898_ (_22794_, _22773_);
  nor _44899_ (_22795_, _22794_, _22740_);
  and _44900_ (_22806_, _22795_, _22729_);
  not _44901_ (_22816_, _22806_);
  and _44902_ (_22827_, _22816_, _20444_);
  and _44903_ (_22838_, _22827_, _22653_);
  and _44904_ (_22849_, _22643_, _20444_);
  not _44905_ (_22860_, _22849_);
  and _44906_ (_22871_, _22816_, _21423_);
  and _44907_ (_22882_, _22871_, _22860_);
  and _44908_ (_22893_, _22882_, _22262_);
  nor _44909_ (_22903_, _22893_, _22838_);
  and _44910_ (_22914_, _22251_, _21423_);
  nor _44911_ (_22925_, _22914_, _21967_);
  nor _44912_ (_22936_, _22925_, _22273_);
  not _44913_ (_22947_, _22936_);
  nor _44914_ (_22958_, _22947_, _22903_);
  nor _44915_ (_22969_, _22306_, _22273_);
  nor _44916_ (_22980_, _22969_, _22316_);
  and _44917_ (_22990_, _22980_, _22958_);
  nor _44918_ (_23001_, _22371_, _22316_);
  nor _44919_ (_23012_, _23001_, _22382_);
  and _44920_ (_23023_, _23012_, _22990_);
  and _44921_ (_23034_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _44922_ (_23055_, _20509_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _44923_ (_23056_, _23055_, _23034_);
  and _44924_ (_23066_, _20586_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _44925_ (_23077_, _20553_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _44926_ (_23088_, _23077_, _23066_);
  and _44927_ (_23099_, _23088_, _23056_);
  and _44928_ (_23110_, _20639_, _20183_);
  and _44929_ (_23121_, _20662_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _44930_ (_23132_, _20683_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _44931_ (_23143_, _23132_, _23121_);
  not _44932_ (_23153_, _23143_);
  nor _44933_ (_23164_, _23153_, _23110_);
  and _44934_ (_23175_, _23164_, _23099_);
  not _44935_ (_23186_, _23175_);
  and _44936_ (_23197_, _23186_, _21423_);
  and _44937_ (_23208_, _23197_, _22849_);
  nor _44938_ (_23219_, _22827_, _22653_);
  nor _44939_ (_23230_, _23219_, _22838_);
  and _44940_ (_23240_, _23230_, _23208_);
  nor _44941_ (_23251_, _22882_, _22262_);
  nor _44942_ (_23262_, _23251_, _22893_);
  and _44943_ (_23273_, _23262_, _23240_);
  and _44944_ (_23284_, _22947_, _22903_);
  nor _44945_ (_23295_, _23284_, _22958_);
  and _44946_ (_23306_, _23295_, _23273_);
  nor _44947_ (_23317_, _22980_, _22958_);
  nor _44948_ (_23338_, _23317_, _22990_);
  and _44949_ (_23339_, _23338_, _23306_);
  nor _44950_ (_23349_, _23012_, _22990_);
  nor _44951_ (_23360_, _23349_, _23023_);
  and _44952_ (_23371_, _23360_, _23339_);
  nor _44953_ (_23382_, _23371_, _23023_);
  nor _44954_ (_23393_, _23382_, _22480_);
  nor _44955_ (_23404_, _23393_, _22447_);
  nor _44956_ (_23415_, _22065_, _21618_);
  nor _44957_ (_23426_, _23415_, _22077_);
  not _44958_ (_23437_, _23426_);
  nor _44959_ (_23448_, _23437_, _23404_);
  or _44960_ (_23458_, _23448_, _22011_);
  nor _44961_ (_23469_, _23458_, _22077_);
  nor _44962_ (_23480_, _23469_, _19687_);
  and _44963_ (_23491_, _23469_, _19687_);
  nor _44964_ (_23502_, _23491_, _23480_);
  not _44965_ (_23513_, _23502_);
  and _44966_ (_23524_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _44967_ (_23535_, _23437_, _23404_);
  nor _44968_ (_23546_, _23535_, _23448_);
  and _44969_ (_23557_, _23546_, _23524_);
  and _44970_ (_23567_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _44971_ (_23578_, _23382_, _22480_);
  nor _44972_ (_23589_, _23578_, _23393_);
  and _44973_ (_23600_, _23589_, _23567_);
  nor _44974_ (_23611_, _23589_, _23567_);
  nor _44975_ (_23622_, _23611_, _23600_);
  not _44976_ (_23633_, _23622_);
  and _44977_ (_23644_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _44978_ (_23655_, _23360_, _23339_);
  nor _44979_ (_23666_, _23655_, _23371_);
  and _44980_ (_23676_, _23666_, _23644_);
  nor _44981_ (_23687_, _23666_, _23644_);
  nor _44982_ (_23698_, _23687_, _23676_);
  not _44983_ (_23709_, _23698_);
  and _44984_ (_23720_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _44985_ (_23731_, _23338_, _23306_);
  nor _44986_ (_23742_, _23731_, _23339_);
  and _44987_ (_23753_, _23742_, _23720_);
  nor _44988_ (_23774_, _23742_, _23720_);
  nor _44989_ (_23775_, _23774_, _23753_);
  not _44990_ (_23786_, _23775_);
  and _44991_ (_23796_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _44992_ (_23807_, _23295_, _23273_);
  nor _44993_ (_23818_, _23807_, _23306_);
  and _44994_ (_23829_, _23818_, _23796_);
  and _44995_ (_23840_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _44996_ (_23851_, _23262_, _23240_);
  nor _44997_ (_23862_, _23851_, _23273_);
  and _44998_ (_23873_, _23862_, _23840_);
  and _44999_ (_23884_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _45000_ (_23895_, _23230_, _23208_);
  nor _45001_ (_23905_, _23895_, _23240_);
  and _45002_ (_23916_, _23905_, _23884_);
  nor _45003_ (_23927_, _23862_, _23840_);
  nor _45004_ (_23938_, _23927_, _23873_);
  and _45005_ (_23959_, _23938_, _23916_);
  nor _45006_ (_23960_, _23959_, _23873_);
  not _45007_ (_23971_, _23960_);
  nor _45008_ (_23982_, _23818_, _23796_);
  nor _45009_ (_23993_, _23982_, _23829_);
  and _45010_ (_24004_, _23993_, _23971_);
  nor _45011_ (_24014_, _24004_, _23829_);
  nor _45012_ (_24025_, _24014_, _23786_);
  nor _45013_ (_24036_, _24025_, _23753_);
  nor _45014_ (_24047_, _24036_, _23709_);
  nor _45015_ (_24058_, _24047_, _23676_);
  nor _45016_ (_24069_, _24058_, _23633_);
  nor _45017_ (_24080_, _24069_, _23600_);
  nor _45018_ (_24090_, _23546_, _23524_);
  nor _45019_ (_24101_, _24090_, _23557_);
  not _45020_ (_24112_, _24101_);
  nor _45021_ (_24123_, _24112_, _24080_);
  nor _45022_ (_24134_, _24123_, _23557_);
  nor _45023_ (_24145_, _24134_, _23513_);
  nor _45024_ (_24156_, _24145_, _23480_);
  not _45025_ (_24167_, _24156_);
  and _45026_ (_24177_, _24167_, _19665_);
  and _45027_ (_24188_, _24177_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _45028_ (_24199_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _45029_ (_24210_, _24199_, _24188_);
  and _45030_ (_24221_, _24210_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _45031_ (_24232_, _24221_, _19654_);
  and _45032_ (_24243_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _45033_ (_24255_, _24243_, _24232_);
  and _45034_ (_24265_, _24232_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _45035_ (_24276_, _24265_, _24255_);
  and _45036_ (_24254_, _24276_, _43634_);
  nor _45037_ (_24297_, _19525_, _19558_);
  and _45038_ (_24308_, _19525_, _19558_);
  or _45039_ (_24319_, _24308_, _24297_);
  and _45040_ (_02349_, _24319_, _43634_);
  and _45041_ (_24340_, _23186_, _20444_);
  and _45042_ (_02541_, _24340_, _43634_);
  nor _45043_ (_24360_, _23197_, _22849_);
  nor _45044_ (_24371_, _24360_, _23208_);
  and _45045_ (_02720_, _24371_, _43634_);
  nor _45046_ (_24392_, _23905_, _23884_);
  nor _45047_ (_24403_, _24392_, _23916_);
  and _45048_ (_02893_, _24403_, _43634_);
  nor _45049_ (_24423_, _23938_, _23916_);
  nor _45050_ (_24434_, _24423_, _23959_);
  and _45051_ (_03129_, _24434_, _43634_);
  nor _45052_ (_24455_, _23993_, _23971_);
  nor _45053_ (_24466_, _24455_, _24004_);
  and _45054_ (_03347_, _24466_, _43634_);
  and _45055_ (_24487_, _24014_, _23786_);
  nor _45056_ (_24498_, _24487_, _24025_);
  and _45057_ (_03548_, _24498_, _43634_);
  and _45058_ (_24518_, _24036_, _23709_);
  nor _45059_ (_24529_, _24518_, _24047_);
  and _45060_ (_03749_, _24529_, _43634_);
  and _45061_ (_24550_, _24058_, _23633_);
  nor _45062_ (_24561_, _24550_, _24069_);
  and _45063_ (_03948_, _24561_, _43634_);
  and _45064_ (_24582_, _24112_, _24080_);
  nor _45065_ (_24592_, _24582_, _24123_);
  and _45066_ (_04045_, _24592_, _43634_);
  and _45067_ (_24613_, _24134_, _23513_);
  nor _45068_ (_24624_, _24613_, _24145_);
  and _45069_ (_04144_, _24624_, _43634_);
  nor _45070_ (_24645_, _24167_, _19665_);
  nor _45071_ (_24656_, _24645_, _24177_);
  and _45072_ (_04243_, _24656_, _43634_);
  and _45073_ (_24676_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _45074_ (_24687_, _24676_, _24177_);
  nor _45075_ (_24698_, _24687_, _24188_);
  and _45076_ (_04343_, _24698_, _43634_);
  nor _45077_ (_24719_, _24199_, _24188_);
  nor _45078_ (_24730_, _24719_, _24210_);
  and _45079_ (_04436_, _24730_, _43634_);
  and _45080_ (_24750_, _19644_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _45081_ (_24761_, _24750_, _24210_);
  nor _45082_ (_24772_, _24761_, _24221_);
  and _45083_ (_04536_, _24772_, _43634_);
  nor _45084_ (_24793_, _24221_, _19654_);
  nor _45085_ (_24804_, _24793_, _24232_);
  and _45086_ (_04634_, _24804_, _43634_);
  and _45087_ (_24825_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _19459_);
  nor _45088_ (_24835_, _24825_, _19470_);
  not _45089_ (_24846_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _45090_ (_24857_, _19492_, _24846_);
  and _45091_ (_24868_, _24857_, _24835_);
  and _45092_ (_24879_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _45093_ (_24890_, _24879_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _45094_ (_24901_, _24879_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45095_ (_24912_, _24901_, _24890_);
  and _45096_ (_00926_, _24912_, _43634_);
  and _45097_ (_00956_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _43634_);
  not _45098_ (_24942_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _45099_ (_24953_, _21227_, _24942_);
  and _45100_ (_24964_, _20912_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45101_ (_24975_, _24964_, _24953_);
  nor _45102_ (_24986_, _24975_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45103_ (_24996_, _21074_, _24942_);
  and _45104_ (_25017_, _21402_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _45105_ (_25018_, _25017_, _24996_);
  and _45106_ (_25029_, _25018_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _45107_ (_25040_, _25029_, _24986_);
  nor _45108_ (_25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _45109_ (_25062_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  and _45110_ (_25073_, _25051_, _21576_);
  nor _45111_ (_25083_, _25073_, _25062_);
  not _45112_ (_25094_, _25083_);
  and _45113_ (_25105_, _20248_, _24942_);
  and _45114_ (_25116_, _19922_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45115_ (_25127_, _25116_, _25105_);
  nor _45116_ (_25138_, _25127_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _45117_ (_25149_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45118_ (_25160_, _20085_, _24942_);
  and _45119_ (_25170_, _20422_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45120_ (_25181_, _25170_, _25160_);
  nor _45121_ (_25192_, _25181_, _25149_);
  nor _45122_ (_25203_, _25192_, _25138_);
  nor _45123_ (_25214_, _25203_, _25094_);
  and _45124_ (_25225_, _25203_, _25094_);
  nor _45125_ (_25236_, _25225_, _25214_);
  and _45126_ (_25247_, _25051_, _20738_);
  nor _45127_ (_25258_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor _45128_ (_25279_, _25258_, _25247_);
  not _45129_ (_25280_, _25279_);
  nor _45130_ (_25291_, _21227_, _24942_);
  nor _45131_ (_25302_, _25291_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45132_ (_25313_, _20912_, _24942_);
  and _45133_ (_25324_, _21074_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45134_ (_25335_, _25324_, _25313_);
  nor _45135_ (_25346_, _25335_, _25149_);
  nor _45136_ (_25357_, _25346_, _25302_);
  nor _45137_ (_25368_, _25357_, _25280_);
  and _45138_ (_25379_, _25357_, _25280_);
  nor _45139_ (_25390_, _25379_, _25368_);
  not _45140_ (_25401_, _25390_);
  nor _45141_ (_25412_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and _45142_ (_25423_, _25051_, _21761_);
  nor _45143_ (_25433_, _25423_, _25412_);
  not _45144_ (_25444_, _25433_);
  nor _45145_ (_25455_, _20248_, _24942_);
  nor _45146_ (_25466_, _25455_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45147_ (_25477_, _19922_, _24942_);
  and _45148_ (_25488_, _20085_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45149_ (_25499_, _25488_, _25477_);
  nor _45150_ (_25510_, _25499_, _25149_);
  nor _45151_ (_25521_, _25510_, _25466_);
  nor _45152_ (_25532_, _25521_, _25444_);
  and _45153_ (_25543_, _25521_, _25444_);
  and _45154_ (_25554_, _24975_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _45155_ (_25565_, _25554_);
  nor _45156_ (_25586_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _45157_ (_25587_, _25051_, _21946_);
  nor _45158_ (_25598_, _25587_, _25586_);
  and _45159_ (_25609_, _25598_, _25565_);
  and _45160_ (_25620_, _25127_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _45161_ (_25631_, _25620_);
  nor _45162_ (_25642_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  and _45163_ (_25653_, _25051_, _22240_);
  nor _45164_ (_25664_, _25653_, _25642_);
  and _45165_ (_25675_, _25664_, _25631_);
  nor _45166_ (_25686_, _25664_, _25631_);
  nor _45167_ (_25697_, _25686_, _25675_);
  not _45168_ (_25708_, _25697_);
  and _45169_ (_25719_, _25291_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _45170_ (_25730_, _25719_);
  and _45171_ (_25741_, _25051_, _22806_);
  nor _45172_ (_25752_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _45173_ (_25763_, _25752_, _25741_);
  and _45174_ (_25774_, _25763_, _25730_);
  and _45175_ (_25785_, _25455_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _45176_ (_25796_, _25785_);
  nor _45177_ (_25807_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and _45178_ (_25818_, _25051_, _22632_);
  nor _45179_ (_25828_, _25818_, _25807_);
  nor _45180_ (_25839_, _25828_, _25796_);
  not _45181_ (_25850_, _25839_);
  nor _45182_ (_25861_, _25763_, _25730_);
  nor _45183_ (_25872_, _25861_, _25774_);
  and _45184_ (_25883_, _25872_, _25850_);
  nor _45185_ (_25894_, _25883_, _25774_);
  nor _45186_ (_25915_, _25894_, _25708_);
  nor _45187_ (_25916_, _25915_, _25675_);
  nor _45188_ (_25927_, _25598_, _25565_);
  nor _45189_ (_25938_, _25927_, _25609_);
  not _45190_ (_25949_, _25938_);
  nor _45191_ (_25960_, _25949_, _25916_);
  nor _45192_ (_25971_, _25960_, _25609_);
  nor _45193_ (_25982_, _25971_, _25543_);
  nor _45194_ (_25993_, _25982_, _25532_);
  nor _45195_ (_26004_, _25993_, _25401_);
  nor _45196_ (_26015_, _26004_, _25368_);
  not _45197_ (_26026_, _26015_);
  and _45198_ (_26037_, _26026_, _25236_);
  or _45199_ (_26048_, _26037_, _25214_);
  and _45200_ (_26059_, _21402_, _20422_);
  or _45201_ (_26070_, _26059_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _45202_ (_26081_, _25181_);
  and _45203_ (_26092_, _25018_, _26081_);
  nor _45204_ (_26103_, _25499_, _25335_);
  and _45205_ (_26114_, _26103_, _26092_);
  or _45206_ (_26125_, _26114_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _45207_ (_26136_, _26125_, _26070_);
  and _45208_ (_26147_, _26136_, _26048_);
  and _45209_ (_26158_, _26147_, _25040_);
  nor _45210_ (_26169_, _26026_, _25236_);
  or _45211_ (_26179_, _26169_, _26037_);
  and _45212_ (_26190_, _26179_, _26158_);
  nor _45213_ (_26201_, _26158_, _25083_);
  nor _45214_ (_26212_, _26201_, _26190_);
  not _45215_ (_26223_, _26212_);
  and _45216_ (_26234_, _26212_, _25040_);
  not _45217_ (_26245_, _25203_);
  nor _45218_ (_26256_, _26158_, _25280_);
  and _45219_ (_26267_, _25993_, _25401_);
  nor _45220_ (_26278_, _26267_, _26004_);
  and _45221_ (_26289_, _26278_, _26158_);
  or _45222_ (_26300_, _26289_, _26256_);
  and _45223_ (_26311_, _26300_, _26245_);
  nor _45224_ (_26322_, _26300_, _26245_);
  nor _45225_ (_26333_, _26322_, _26311_);
  not _45226_ (_26344_, _26333_);
  not _45227_ (_26355_, _25357_);
  nor _45228_ (_26366_, _26158_, _25444_);
  nor _45229_ (_26377_, _25543_, _25532_);
  nor _45230_ (_26398_, _26377_, _25971_);
  and _45231_ (_26399_, _26377_, _25971_);
  or _45232_ (_26410_, _26399_, _26398_);
  and _45233_ (_26421_, _26410_, _26158_);
  or _45234_ (_26432_, _26421_, _26366_);
  and _45235_ (_26443_, _26432_, _26355_);
  nor _45236_ (_26454_, _26432_, _26355_);
  not _45237_ (_26465_, _25521_);
  and _45238_ (_26476_, _25949_, _25916_);
  or _45239_ (_26487_, _26476_, _25960_);
  and _45240_ (_26498_, _26487_, _26158_);
  nor _45241_ (_26509_, _26158_, _25598_);
  nor _45242_ (_26520_, _26509_, _26498_);
  and _45243_ (_26530_, _26520_, _26465_);
  and _45244_ (_26541_, _25894_, _25708_);
  nor _45245_ (_26552_, _26541_, _25915_);
  not _45246_ (_26563_, _26552_);
  and _45247_ (_26574_, _26563_, _26158_);
  nor _45248_ (_26585_, _26158_, _25664_);
  nor _45249_ (_26596_, _26585_, _26574_);
  and _45250_ (_26607_, _26596_, _25565_);
  nor _45251_ (_26628_, _26596_, _25565_);
  nor _45252_ (_26629_, _26628_, _26607_);
  not _45253_ (_26640_, _26629_);
  nor _45254_ (_26651_, _25872_, _25850_);
  nor _45255_ (_26662_, _26651_, _25883_);
  not _45256_ (_26673_, _26662_);
  and _45257_ (_26684_, _26673_, _26158_);
  nor _45258_ (_26695_, _26158_, _25763_);
  nor _45259_ (_26706_, _26695_, _26684_);
  and _45260_ (_26717_, _26706_, _25631_);
  not _45261_ (_26728_, _25828_);
  and _45262_ (_26739_, _26158_, _25785_);
  or _45263_ (_26750_, _26739_, _26728_);
  nand _45264_ (_26761_, _26158_, _25785_);
  or _45265_ (_26772_, _26761_, _25828_);
  and _45266_ (_26783_, _26772_, _26750_);
  nor _45267_ (_26794_, _26783_, _25719_);
  and _45268_ (_26805_, _26783_, _25719_);
  nor _45269_ (_26816_, _26805_, _26794_);
  nor _45270_ (_26827_, _25051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _45271_ (_26838_, _25051_, _23175_);
  nor _45272_ (_26849_, _26838_, _26827_);
  nor _45273_ (_26860_, _26849_, _25796_);
  not _45274_ (_26871_, _26860_);
  and _45275_ (_26882_, _26871_, _26816_);
  nor _45276_ (_26892_, _26882_, _26794_);
  nor _45277_ (_26903_, _26706_, _25631_);
  nor _45278_ (_26914_, _26903_, _26717_);
  not _45279_ (_26925_, _26914_);
  nor _45280_ (_26936_, _26925_, _26892_);
  nor _45281_ (_26947_, _26936_, _26717_);
  nor _45282_ (_26958_, _26947_, _26640_);
  nor _45283_ (_26969_, _26958_, _26607_);
  nor _45284_ (_26980_, _26520_, _26465_);
  nor _45285_ (_26991_, _26980_, _26530_);
  not _45286_ (_27002_, _26991_);
  nor _45287_ (_27013_, _27002_, _26969_);
  nor _45288_ (_27024_, _27013_, _26530_);
  nor _45289_ (_27035_, _27024_, _26454_);
  nor _45290_ (_27046_, _27035_, _26443_);
  nor _45291_ (_27057_, _27046_, _26344_);
  or _45292_ (_27068_, _27057_, _26311_);
  or _45293_ (_27079_, _27068_, _26234_);
  and _45294_ (_27090_, _27079_, _26136_);
  nor _45295_ (_27101_, _27090_, _26223_);
  and _45296_ (_27112_, _26234_, _26136_);
  and _45297_ (_27123_, _27112_, _27068_);
  or _45298_ (_27134_, _27123_, _27101_);
  and _45299_ (_00976_, _27134_, _43634_);
  or _45300_ (_27155_, _26212_, _25040_);
  and _45301_ (_27166_, _27155_, _27090_);
  and _45302_ (_02847_, _27166_, _43634_);
  and _45303_ (_02859_, _26158_, _43634_);
  and _45304_ (_02881_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _43634_);
  and _45305_ (_02906_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _43634_);
  and _45306_ (_02931_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _43634_);
  or _45307_ (_27227_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _45308_ (_27237_, _24879_, rst);
  and _45309_ (_02942_, _27237_, _27227_);
  and _45310_ (_27258_, _27166_, _25785_);
  or _45311_ (_27269_, _27258_, _26849_);
  nand _45312_ (_27280_, _27258_, _26849_);
  and _45313_ (_27291_, _27280_, _27269_);
  and _45314_ (_02955_, _27291_, _43634_);
  nor _45315_ (_27312_, _27166_, _26783_);
  nor _45316_ (_27323_, _26871_, _26816_);
  nor _45317_ (_27334_, _27323_, _26882_);
  and _45318_ (_27345_, _27334_, _27166_);
  or _45319_ (_27356_, _27345_, _27312_);
  and _45320_ (_02968_, _27356_, _43634_);
  and _45321_ (_27377_, _26925_, _26892_);
  or _45322_ (_27388_, _27377_, _26936_);
  nand _45323_ (_27399_, _27388_, _27166_);
  or _45324_ (_27410_, _27166_, _26706_);
  and _45325_ (_27421_, _27410_, _27399_);
  and _45326_ (_02980_, _27421_, _43634_);
  and _45327_ (_27442_, _26947_, _26640_);
  or _45328_ (_27453_, _27442_, _26958_);
  nand _45329_ (_27464_, _27453_, _27166_);
  or _45330_ (_27475_, _27166_, _26596_);
  and _45331_ (_27486_, _27475_, _27464_);
  and _45332_ (_02992_, _27486_, _43634_);
  and _45333_ (_27507_, _27002_, _26969_);
  or _45334_ (_27518_, _27507_, _27013_);
  nand _45335_ (_27529_, _27518_, _27166_);
  or _45336_ (_27540_, _27166_, _26520_);
  and _45337_ (_27551_, _27540_, _27529_);
  and _45338_ (_03005_, _27551_, _43634_);
  or _45339_ (_27572_, _26454_, _26443_);
  and _45340_ (_27582_, _27572_, _27024_);
  nor _45341_ (_27593_, _27572_, _27024_);
  or _45342_ (_27604_, _27593_, _27582_);
  nand _45343_ (_27615_, _27604_, _27166_);
  or _45344_ (_27626_, _27166_, _26432_);
  and _45345_ (_27637_, _27626_, _27615_);
  and _45346_ (_03016_, _27637_, _43634_);
  and _45347_ (_27658_, _27046_, _26344_);
  or _45348_ (_27669_, _27658_, _27057_);
  nand _45349_ (_27680_, _27669_, _27166_);
  or _45350_ (_27691_, _27166_, _26300_);
  and _45351_ (_27702_, _27691_, _27680_);
  and _45352_ (_03029_, _27702_, _43634_);
  not _45353_ (_27723_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _45354_ (_27734_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _19459_);
  and _45355_ (_27745_, _27734_, _27723_);
  and _45356_ (_27756_, _27745_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _45357_ (_27767_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _45358_ (_27778_, _27767_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _45359_ (_27789_, _27767_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _45360_ (_27800_, _27789_, _27778_);
  and _45361_ (_27811_, _27800_, _27756_);
  not _45362_ (_27832_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _45363_ (_27833_, _27745_, _27832_);
  and _45364_ (_27844_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _45365_ (_27855_, _27844_, _27811_);
  not _45366_ (_27866_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _45367_ (_27877_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _19459_);
  and _45368_ (_27888_, _27877_, _27866_);
  and _45369_ (_27899_, _27888_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _45370_ (_27910_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _45371_ (_27921_, _27888_, _27723_);
  and _45372_ (_27932_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or _45373_ (_27942_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _45374_ (_27953_, _27942_, _19459_);
  nor _45375_ (_27964_, _27953_, _27877_);
  and _45376_ (_27975_, _27964_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _45377_ (_27986_, _27975_, _27932_);
  nor _45378_ (_27997_, _27986_, _27910_);
  and _45379_ (_28008_, _27997_, _27855_);
  nor _45380_ (_28019_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _45381_ (_28030_, _28019_, _27767_);
  and _45382_ (_28041_, _28030_, _27756_);
  and _45383_ (_28052_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _45384_ (_28063_, _28052_, _28041_);
  and _45385_ (_28074_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _45386_ (_28085_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _45387_ (_28096_, _27964_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _45388_ (_28107_, _28096_, _28085_);
  nor _45389_ (_28118_, _28107_, _28074_);
  and _45390_ (_28139_, _28118_, _28063_);
  and _45391_ (_28140_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and _45392_ (_28151_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _45393_ (_28162_, _28151_, _28140_);
  and _45394_ (_28173_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _45395_ (_28184_, _28173_);
  not _45396_ (_28195_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _45397_ (_28206_, _27756_, _28195_);
  and _45398_ (_28217_, _27964_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _45399_ (_28228_, _28217_, _28206_);
  and _45400_ (_28239_, _28228_, _28184_);
  and _45401_ (_28250_, _28239_, _28162_);
  and _45402_ (_28260_, _28250_, _28139_);
  and _45403_ (_28271_, _28260_, _28008_);
  and _45404_ (_28282_, _27778_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _45405_ (_28293_, _28282_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _45406_ (_28304_, _28293_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _45407_ (_28315_, _28304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _45408_ (_28326_, _28315_);
  not _45409_ (_28337_, _27756_);
  nor _45410_ (_28348_, _28304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _45411_ (_28359_, _28348_, _28337_);
  and _45412_ (_28370_, _28359_, _28326_);
  not _45413_ (_28381_, _28370_);
  and _45414_ (_28392_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _45415_ (_28403_, _28392_, _27734_);
  and _45416_ (_28414_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _45417_ (_28425_, _28414_, _28403_);
  and _45418_ (_28436_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _45419_ (_28447_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _45420_ (_28458_, _28447_, _28436_);
  and _45421_ (_28469_, _28458_, _28425_);
  and _45422_ (_28490_, _28469_, _28381_);
  nor _45423_ (_28491_, _28293_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _45424_ (_28502_, _28491_);
  nor _45425_ (_28513_, _28304_, _28337_);
  and _45426_ (_28524_, _28513_, _28502_);
  not _45427_ (_28535_, _28524_);
  and _45428_ (_28546_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _45429_ (_28557_, _28546_, _28403_);
  and _45430_ (_28568_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _45431_ (_28579_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _45432_ (_28589_, _28579_, _28568_);
  and _45433_ (_28600_, _28589_, _28557_);
  and _45434_ (_28611_, _28600_, _28535_);
  nor _45435_ (_28622_, _28611_, _28490_);
  not _45436_ (_28633_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _45437_ (_28644_, _28315_, _28633_);
  and _45438_ (_28655_, _28315_, _28633_);
  nor _45439_ (_28666_, _28655_, _28644_);
  nor _45440_ (_28677_, _28666_, _28337_);
  not _45441_ (_28688_, _28677_);
  and _45442_ (_28699_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _45443_ (_28710_, _28699_, _28403_);
  and _45444_ (_28721_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _45445_ (_28732_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _45446_ (_28743_, _28732_, _28721_);
  and _45447_ (_28754_, _28743_, _28710_);
  and _45448_ (_28765_, _28754_, _28688_);
  not _45449_ (_28776_, _28765_);
  and _45450_ (_28787_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _45451_ (_28798_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _45452_ (_28809_, _28798_, _28787_);
  not _45453_ (_28820_, _28282_);
  nor _45454_ (_28831_, _27778_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _45455_ (_28842_, _28831_, _28337_);
  and _45456_ (_28863_, _28842_, _28820_);
  and _45457_ (_28864_, _27964_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _45458_ (_28875_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _45459_ (_28885_, _28875_, _28864_);
  not _45460_ (_28896_, _28885_);
  nor _45461_ (_28907_, _28896_, _28863_);
  and _45462_ (_28918_, _28907_, _28809_);
  not _45463_ (_28929_, _28918_);
  and _45464_ (_28940_, _27899_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor _45465_ (_28951_, _28940_, _28403_);
  nor _45466_ (_28962_, _28282_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _45467_ (_28973_, _28962_, _28337_);
  nor _45468_ (_28984_, _28973_, _28293_);
  and _45469_ (_28995_, _27921_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _45470_ (_29006_, _28995_, _28984_);
  and _45471_ (_29017_, _29006_, _28951_);
  and _45472_ (_29028_, _27964_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _45473_ (_29039_, _27833_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _45474_ (_29050_, _29039_, _29028_);
  and _45475_ (_29061_, _29050_, _29017_);
  nor _45476_ (_29072_, _29061_, _28929_);
  and _45477_ (_29083_, _29072_, _28776_);
  and _45478_ (_29094_, _29083_, _28622_);
  nand _45479_ (_29105_, _29094_, _28271_);
  and _45480_ (_29116_, _27134_, _24868_);
  not _45481_ (_29127_, _29116_);
  and _45482_ (_29138_, _24276_, _19525_);
  not _45483_ (_29149_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _45484_ (_29160_, _19470_, _29149_);
  and _45485_ (_29171_, _29160_, _19514_);
  not _45486_ (_29182_, _29171_);
  nor _45487_ (_29192_, _21576_, _21402_);
  and _45488_ (_29203_, _21576_, _21402_);
  nor _45489_ (_29214_, _29203_, _29192_);
  and _45490_ (_29225_, _20749_, _20422_);
  nor _45491_ (_29236_, _20738_, _20422_);
  and _45492_ (_29247_, _20738_, _20422_);
  nor _45493_ (_29258_, _29247_, _29236_);
  not _45494_ (_29269_, _21074_);
  nor _45495_ (_29280_, _21761_, _29269_);
  nor _45496_ (_29291_, _21761_, _21074_);
  and _45497_ (_29302_, _21761_, _21074_);
  nor _45498_ (_29313_, _29302_, _29291_);
  not _45499_ (_29324_, _20085_);
  and _45500_ (_29335_, _21946_, _29324_);
  nor _45501_ (_29346_, _29335_, _29313_);
  nor _45502_ (_29357_, _29346_, _29280_);
  nor _45503_ (_29368_, _29357_, _29258_);
  nor _45504_ (_29389_, _29368_, _29225_);
  and _45505_ (_29390_, _29357_, _29258_);
  nor _45506_ (_29401_, _29390_, _29368_);
  not _45507_ (_29412_, _29401_);
  and _45508_ (_29423_, _29335_, _29313_);
  nor _45509_ (_29434_, _29423_, _29346_);
  not _45510_ (_29445_, _29434_);
  nor _45511_ (_29456_, _21946_, _20085_);
  and _45512_ (_29467_, _21946_, _20085_);
  nor _45513_ (_29478_, _29467_, _29456_);
  not _45514_ (_29489_, _29478_);
  and _45515_ (_29499_, _22240_, _20912_);
  nor _45516_ (_29510_, _22240_, _20912_);
  nor _45517_ (_29521_, _29510_, _29499_);
  not _45518_ (_29532_, _29521_);
  nor _45519_ (_29543_, _22806_, _19922_);
  and _45520_ (_29554_, _22806_, _19922_);
  nor _45521_ (_29565_, _29554_, _29543_);
  nor _45522_ (_29576_, _22632_, _21227_);
  and _45523_ (_29587_, _22632_, _21227_);
  nor _45524_ (_29598_, _29587_, _29576_);
  not _45525_ (_29609_, _20248_);
  and _45526_ (_29620_, _23175_, _29609_);
  nor _45527_ (_29631_, _29620_, _29598_);
  not _45528_ (_29642_, _21227_);
  nor _45529_ (_29663_, _22632_, _29642_);
  nor _45530_ (_29664_, _29663_, _29631_);
  nor _45531_ (_29675_, _29664_, _29565_);
  not _45532_ (_29686_, _19922_);
  nor _45533_ (_29697_, _22806_, _29686_);
  nor _45534_ (_29708_, _29697_, _29675_);
  nor _45535_ (_29719_, _29708_, _29532_);
  and _45536_ (_29730_, _29708_, _29532_);
  nor _45537_ (_29741_, _29730_, _29719_);
  nor _45538_ (_29752_, _23175_, _20248_);
  and _45539_ (_29763_, _23175_, _20248_);
  nor _45540_ (_29774_, _29763_, _29752_);
  not _45541_ (_29785_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _45542_ (_29796_, _19743_, _29785_);
  not _45543_ (_29806_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _45544_ (_29817_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45545_ (_29828_, _29817_, _21293_);
  nor _45546_ (_29839_, _29828_, _29806_);
  nor _45547_ (_29850_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45548_ (_29861_, _29850_, _19977_);
  not _45549_ (_29872_, _29861_);
  not _45550_ (_29883_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45551_ (_29894_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _29883_);
  and _45552_ (_29905_, _29894_, _20955_);
  not _45553_ (_29916_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _45554_ (_29927_, _29916_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _45555_ (_29938_, _29927_, _20314_);
  nor _45556_ (_29949_, _29938_, _29905_);
  and _45557_ (_29960_, _29949_, _29872_);
  and _45558_ (_29971_, _29960_, _29839_);
  and _45559_ (_29982_, _29817_, _20803_);
  nor _45560_ (_29993_, _29982_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _45561_ (_30004_, _29927_, _19791_);
  not _45562_ (_30015_, _30004_);
  and _45563_ (_30026_, _29894_, _21119_);
  and _45564_ (_30037_, _29850_, _20140_);
  nor _45565_ (_30048_, _30037_, _30026_);
  and _45566_ (_30059_, _30048_, _30015_);
  and _45567_ (_30070_, _30059_, _29993_);
  nor _45568_ (_30081_, _30070_, _29971_);
  nor _45569_ (_30092_, _30081_, _19743_);
  nor _45570_ (_30102_, _30092_, _29796_);
  and _45571_ (_30113_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _45572_ (_30124_, _30113_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _45573_ (_30135_, _30124_);
  and _45574_ (_30146_, _30135_, _30102_);
  and _45575_ (_30157_, _30135_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _45576_ (_30168_, _30157_, _30146_);
  nor _45577_ (_30179_, _30168_, _29774_);
  and _45578_ (_30190_, _29664_, _29565_);
  nor _45579_ (_30201_, _30190_, _29675_);
  and _45580_ (_30212_, _29620_, _29598_);
  nor _45581_ (_30223_, _30212_, _29631_);
  nor _45582_ (_30234_, _30223_, _30201_);
  and _45583_ (_30244_, _30234_, _30179_);
  and _45584_ (_30255_, _30244_, _29741_);
  not _45585_ (_30266_, _20912_);
  or _45586_ (_30287_, _22240_, _30266_);
  and _45587_ (_30288_, _22240_, _30266_);
  or _45588_ (_30299_, _29708_, _30288_);
  and _45589_ (_30310_, _30299_, _30287_);
  or _45590_ (_30321_, _30310_, _30255_);
  and _45591_ (_30332_, _30321_, _29489_);
  and _45592_ (_30343_, _30332_, _29445_);
  and _45593_ (_30354_, _30343_, _29412_);
  nor _45594_ (_30365_, _30354_, _29389_);
  nor _45595_ (_30376_, _30365_, _29214_);
  and _45596_ (_30387_, _30365_, _29214_);
  nor _45597_ (_30397_, _30387_, _30376_);
  nor _45598_ (_30408_, _30397_, _29182_);
  not _45599_ (_30419_, _30408_);
  not _45600_ (_30430_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _45601_ (_30441_, _24825_, _30430_);
  and _45602_ (_30452_, _30441_, _19514_);
  not _45603_ (_30463_, _29214_);
  not _45604_ (_30474_, _29258_);
  and _45605_ (_30485_, _29456_, _29313_);
  nor _45606_ (_30496_, _30485_, _29291_);
  nor _45607_ (_30507_, _30496_, _30474_);
  not _45608_ (_30518_, _29565_);
  and _45609_ (_30529_, _29752_, _29598_);
  nor _45610_ (_30539_, _30529_, _29576_);
  nor _45611_ (_30550_, _30539_, _30518_);
  nor _45612_ (_30561_, _30550_, _29543_);
  nor _45613_ (_30572_, _30561_, _29521_);
  and _45614_ (_30583_, _30561_, _29521_);
  nor _45615_ (_30594_, _30583_, _30572_);
  not _45616_ (_30605_, _29774_);
  nor _45617_ (_30616_, _30168_, _30605_);
  and _45618_ (_30627_, _30616_, _29598_);
  and _45619_ (_30638_, _30539_, _30518_);
  nor _45620_ (_30649_, _30638_, _30550_);
  and _45621_ (_30660_, _30649_, _30627_);
  not _45622_ (_30671_, _30660_);
  nor _45623_ (_30682_, _30671_, _30594_);
  nor _45624_ (_30692_, _30561_, _29499_);
  or _45625_ (_30703_, _30692_, _29510_);
  or _45626_ (_30714_, _30703_, _30682_);
  and _45627_ (_30725_, _30714_, _29478_);
  nor _45628_ (_30736_, _29456_, _29313_);
  nor _45629_ (_30747_, _30736_, _30485_);
  and _45630_ (_30758_, _30747_, _30725_);
  and _45631_ (_30769_, _30496_, _30474_);
  nor _45632_ (_30780_, _30769_, _30507_);
  and _45633_ (_30791_, _30780_, _30758_);
  or _45634_ (_30802_, _30791_, _30507_);
  nor _45635_ (_30813_, _30802_, _29236_);
  nor _45636_ (_30824_, _30813_, _30463_);
  and _45637_ (_30835_, _30813_, _30463_);
  nor _45638_ (_30845_, _30835_, _30824_);
  and _45639_ (_30856_, _30845_, _30452_);
  and _45640_ (_30867_, _19503_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45641_ (_30878_, _30867_, _29160_);
  nor _45642_ (_30889_, _23175_, _22632_);
  and _45643_ (_30900_, _30889_, _22816_);
  and _45644_ (_30911_, _30900_, _22251_);
  and _45645_ (_30922_, _30911_, _21957_);
  and _45646_ (_30933_, _30922_, _21772_);
  and _45647_ (_30944_, _30933_, _20749_);
  and _45648_ (_30955_, _30944_, _30168_);
  not _45649_ (_30966_, _30168_);
  and _45650_ (_30977_, _20738_, _21761_);
  and _45651_ (_30998_, _23175_, _22632_);
  and _45652_ (_30999_, _30998_, _22806_);
  and _45653_ (_31021_, _30999_, _22240_);
  and _45654_ (_31022_, _31021_, _21946_);
  and _45655_ (_31044_, _31022_, _30977_);
  and _45656_ (_31045_, _31044_, _30966_);
  nor _45657_ (_31067_, _31045_, _30955_);
  and _45658_ (_31068_, _31067_, _21576_);
  nor _45659_ (_31079_, _31067_, _21576_);
  nor _45660_ (_31090_, _31079_, _31068_);
  and _45661_ (_31101_, _31090_, _30878_);
  not _45662_ (_31112_, _21402_);
  nor _45663_ (_31123_, _30168_, _31112_);
  not _45664_ (_31134_, _31123_);
  and _45665_ (_31144_, _30168_, _21576_);
  and _45666_ (_31155_, _30867_, _19481_);
  not _45667_ (_31166_, _31155_);
  nor _45668_ (_31177_, _31166_, _31144_);
  and _45669_ (_31188_, _31177_, _31134_);
  nor _45670_ (_31199_, _31188_, _31101_);
  and _45671_ (_31210_, _30441_, _24857_);
  not _45672_ (_31221_, _30977_);
  and _45673_ (_31232_, _22806_, _22632_);
  nor _45674_ (_31243_, _31232_, _22240_);
  and _45675_ (_31253_, _31243_, _31210_);
  and _45676_ (_31264_, _31253_, _21957_);
  nor _45677_ (_31275_, _31264_, _31221_);
  nor _45678_ (_31286_, _30977_, _21576_);
  nor _45679_ (_31297_, _31286_, _31253_);
  and _45680_ (_31308_, _31297_, _30168_);
  nor _45681_ (_31319_, _31308_, _31275_);
  nor _45682_ (_31330_, _31319_, _21587_);
  and _45683_ (_31341_, _31319_, _21587_);
  nor _45684_ (_31352_, _31341_, _31330_);
  and _45685_ (_31362_, _31352_, _31210_);
  and _45686_ (_31373_, _30867_, _30441_);
  not _45687_ (_31384_, _31373_);
  nor _45688_ (_31395_, _31384_, _30168_);
  not _45689_ (_31406_, _31395_);
  not _45690_ (_31417_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45691_ (_31428_, _19503_, _31417_);
  and _45692_ (_31439_, _31428_, _30441_);
  not _45693_ (_31450_, _31439_);
  nor _45694_ (_31461_, _31450_, _29203_);
  and _45695_ (_31471_, _31428_, _24835_);
  and _45696_ (_31482_, _31471_, _29214_);
  nor _45697_ (_31493_, _31482_, _31461_);
  and _45698_ (_31504_, _24857_, _19481_);
  and _45699_ (_31515_, _31504_, _29192_);
  and _45700_ (_31526_, _29160_, _24857_);
  and _45701_ (_31537_, _31526_, _21576_);
  nor _45702_ (_31548_, _31537_, _31515_);
  and _45703_ (_31559_, _31428_, _19470_);
  not _45704_ (_31570_, _31559_);
  nor _45705_ (_31580_, _31570_, _20738_);
  not _45706_ (_31591_, _31580_);
  and _45707_ (_31602_, _24835_, _19514_);
  not _45708_ (_31613_, _31602_);
  nor _45709_ (_31624_, _31613_, _21576_);
  and _45710_ (_31635_, _30867_, _24835_);
  not _45711_ (_31646_, _31635_);
  nor _45712_ (_31657_, _31646_, _23175_);
  nor _45713_ (_31668_, _31657_, _31624_);
  and _45714_ (_31679_, _31668_, _31591_);
  and _45715_ (_31690_, _31679_, _31548_);
  and _45716_ (_31700_, _31690_, _31493_);
  and _45717_ (_31711_, _31700_, _31406_);
  not _45718_ (_31722_, _31711_);
  nor _45719_ (_31733_, _31722_, _31362_);
  and _45720_ (_31744_, _31733_, _31199_);
  not _45721_ (_31755_, _31744_);
  nor _45722_ (_31766_, _31755_, _30856_);
  and _45723_ (_31777_, _31766_, _30419_);
  not _45724_ (_31788_, _31777_);
  nor _45725_ (_31799_, _31788_, _29138_);
  and _45726_ (_31809_, _31799_, _29127_);
  not _45727_ (_31820_, _31809_);
  or _45728_ (_31831_, _31820_, _29105_);
  not _45729_ (_31842_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45730_ (_31853_, \oc8051_top_1.oc8051_decoder1.wr , _19459_);
  not _45731_ (_31864_, _31853_);
  nor _45732_ (_31875_, _31864_, _27745_);
  and _45733_ (_31886_, _31875_, _31842_);
  not _45734_ (_31897_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _45735_ (_31908_, _29105_, _31897_);
  and _45736_ (_31918_, _31908_, _31886_);
  and _45737_ (_31929_, _31918_, _31831_);
  nor _45738_ (_31940_, _31875_, _31897_);
  not _45739_ (_31951_, _30452_);
  nor _45740_ (_31962_, _30824_, _29192_);
  nor _45741_ (_31973_, _31962_, _31951_);
  not _45742_ (_31984_, _31973_);
  and _45743_ (_31995_, _21576_, _31112_);
  nor _45744_ (_32006_, _31995_, _30376_);
  nor _45745_ (_32017_, _32006_, _29182_);
  not _45746_ (_32027_, _31210_);
  and _45747_ (_32038_, _31286_, _30168_);
  not _45748_ (_32049_, _32038_);
  nor _45749_ (_32060_, _31286_, _30168_);
  nor _45750_ (_32071_, _32060_, _31243_);
  and _45751_ (_32082_, _32071_, _32049_);
  nor _45752_ (_32093_, _32082_, _32027_);
  not _45753_ (_32104_, _32093_);
  nor _45754_ (_32115_, _30157_, _30102_);
  not _45755_ (_32126_, _31471_);
  nor _45756_ (_32136_, _32126_, _30146_);
  not _45757_ (_32147_, _32136_);
  nor _45758_ (_32158_, _31646_, _30102_);
  nor _45759_ (_32169_, _32158_, _31439_);
  and _45760_ (_32180_, _32169_, _32147_);
  nor _45761_ (_32191_, _32180_, _32115_);
  not _45762_ (_32202_, _32191_);
  and _45763_ (_32213_, _30124_, _30102_);
  and _45764_ (_32224_, _31428_, _29160_);
  and _45765_ (_32235_, _31504_, _30102_);
  nor _45766_ (_32245_, _32235_, _32224_);
  nor _45767_ (_32256_, _32245_, _32213_);
  nor _45768_ (_32267_, _31384_, _23175_);
  and _45769_ (_32278_, _31428_, _19481_);
  not _45770_ (_32289_, _32278_);
  nor _45771_ (_32300_, _32289_, _21576_);
  nor _45772_ (_32311_, _32300_, _32267_);
  not _45773_ (_32322_, _32311_);
  nor _45774_ (_32333_, _32322_, _32256_);
  nor _45775_ (_32344_, _31613_, _30168_);
  and _45776_ (_32354_, _31526_, _30168_);
  nor _45777_ (_32365_, _32354_, _32344_);
  and _45778_ (_32376_, _32365_, _32333_);
  and _45779_ (_32387_, _32376_, _32202_);
  and _45780_ (_32398_, _32387_, _32104_);
  not _45781_ (_32409_, _32398_);
  nor _45782_ (_32420_, _32409_, _32017_);
  and _45783_ (_32431_, _32420_, _31984_);
  not _45784_ (_32442_, _28008_);
  nor _45785_ (_32453_, _28250_, _28139_);
  and _45786_ (_32463_, _32453_, _32442_);
  and _45787_ (_32474_, _32463_, _29094_);
  nand _45788_ (_32485_, _32474_, _32431_);
  or _45789_ (_32496_, _32474_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _45790_ (_32507_, _31875_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45791_ (_32518_, _32507_, _32496_);
  and _45792_ (_32529_, _32518_, _32485_);
  or _45793_ (_32540_, _32529_, _31940_);
  or _45794_ (_32551_, _32540_, _31929_);
  and _45795_ (_06648_, _32551_, _43634_);
  and _45796_ (_32572_, _27291_, _24868_);
  not _45797_ (_32582_, _32572_);
  and _45798_ (_32593_, _24592_, _19525_);
  nor _45799_ (_32604_, _32126_, _29752_);
  nor _45800_ (_32615_, _32604_, _31439_);
  or _45801_ (_32626_, _32615_, _29763_);
  and _45802_ (_32637_, _30867_, _30430_);
  not _45803_ (_32648_, _32637_);
  nor _45804_ (_32659_, _32648_, _22632_);
  and _45805_ (_32670_, _32224_, _21587_);
  nor _45806_ (_32681_, _32670_, _32659_);
  and _45807_ (_32691_, _32681_, _32626_);
  nor _45808_ (_32702_, _32289_, _30168_);
  nor _45809_ (_32713_, _31166_, _20248_);
  and _45810_ (_32724_, _30878_, _23175_);
  nor _45811_ (_32735_, _32724_, _32713_);
  nor _45812_ (_32746_, _31602_, _31210_);
  nor _45813_ (_32757_, _32746_, _23175_);
  not _45814_ (_32768_, _32757_);
  nand _45815_ (_32779_, _32768_, _32735_);
  nor _45816_ (_32789_, _32779_, _32702_);
  and _45817_ (_32800_, _32789_, _32691_);
  and _45818_ (_32811_, _30168_, _30605_);
  nor _45819_ (_32822_, _32811_, _30616_);
  not _45820_ (_32833_, _32822_);
  nor _45821_ (_32844_, _30452_, _29171_);
  nor _45822_ (_32855_, _32844_, _32833_);
  not _45823_ (_32866_, _32855_);
  and _45824_ (_32877_, _31504_, _29752_);
  and _45825_ (_32888_, _31526_, _23175_);
  nor _45826_ (_32899_, _32888_, _32877_);
  and _45827_ (_32909_, _32899_, _32866_);
  and _45828_ (_32920_, _32909_, _32800_);
  not _45829_ (_32931_, _32920_);
  nor _45830_ (_32942_, _32931_, _32593_);
  and _45831_ (_32953_, _32942_, _32582_);
  not _45832_ (_32964_, _32953_);
  or _45833_ (_32975_, _32964_, _29105_);
  not _45834_ (_32986_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _45835_ (_32997_, _29105_, _32986_);
  and _45836_ (_33008_, _32997_, _31886_);
  and _45837_ (_33018_, _33008_, _32975_);
  nor _45838_ (_33029_, _31875_, _32986_);
  not _45839_ (_33040_, _32431_);
  or _45840_ (_33051_, _33040_, _29105_);
  and _45841_ (_33062_, _32997_, _32507_);
  and _45842_ (_33073_, _33062_, _33051_);
  or _45843_ (_33084_, _33073_, _33029_);
  or _45844_ (_33095_, _33084_, _33018_);
  and _45845_ (_08889_, _33095_, _43634_);
  and _45846_ (_33116_, _24624_, _19525_);
  not _45847_ (_33126_, _33116_);
  and _45848_ (_33137_, _27356_, _24868_);
  nor _45849_ (_33148_, _31166_, _21227_);
  nor _45850_ (_33159_, _30998_, _30889_);
  not _45851_ (_33170_, _33159_);
  nor _45852_ (_33181_, _33170_, _30168_);
  and _45853_ (_33192_, _33170_, _30168_);
  nor _45854_ (_33203_, _33192_, _33181_);
  and _45855_ (_33214_, _33203_, _30878_);
  nor _45856_ (_33225_, _33214_, _33148_);
  nor _45857_ (_33235_, _31243_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _45858_ (_33246_, _33235_, _22643_);
  nor _45859_ (_33257_, _33235_, _22643_);
  nor _45860_ (_33268_, _33257_, _33246_);
  nor _45861_ (_33279_, _33268_, _32027_);
  not _45862_ (_33290_, _33279_);
  and _45863_ (_33301_, _31471_, _29598_);
  and _45864_ (_33312_, _31504_, _29576_);
  nor _45865_ (_33323_, _31450_, _29587_);
  and _45866_ (_33334_, _31526_, _22632_);
  or _45867_ (_33345_, _33334_, _33323_);
  or _45868_ (_33355_, _33345_, _33312_);
  nor _45869_ (_33366_, _33355_, _33301_);
  nor _45870_ (_33377_, _31570_, _23175_);
  not _45871_ (_33388_, _33377_);
  nor _45872_ (_33399_, _31613_, _22632_);
  nor _45873_ (_33410_, _32648_, _22806_);
  nor _45874_ (_33421_, _33410_, _33399_);
  and _45875_ (_33432_, _33421_, _33388_);
  and _45876_ (_33443_, _33432_, _33366_);
  and _45877_ (_33454_, _33443_, _33290_);
  and _45878_ (_33464_, _33454_, _33225_);
  nor _45879_ (_33475_, _29752_, _29598_);
  or _45880_ (_33486_, _33475_, _30529_);
  and _45881_ (_33497_, _33486_, _30616_);
  nor _45882_ (_33508_, _33486_, _30616_);
  or _45883_ (_33519_, _33508_, _33497_);
  and _45884_ (_33530_, _33519_, _30452_);
  not _45885_ (_33541_, _30223_);
  and _45886_ (_33552_, _33541_, _30179_);
  nor _45887_ (_33562_, _33541_, _30179_);
  nor _45888_ (_33573_, _33562_, _33552_);
  nor _45889_ (_33584_, _33573_, _29182_);
  nor _45890_ (_33595_, _33584_, _33530_);
  and _45891_ (_33606_, _33595_, _33464_);
  not _45892_ (_33617_, _33606_);
  nor _45893_ (_33628_, _33617_, _33137_);
  and _45894_ (_33639_, _33628_, _33126_);
  not _45895_ (_33650_, _33639_);
  or _45896_ (_33661_, _33650_, _29105_);
  not _45897_ (_33672_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _45898_ (_33682_, _29105_, _33672_);
  and _45899_ (_33693_, _33682_, _31886_);
  and _45900_ (_33704_, _33693_, _33661_);
  nor _45901_ (_33715_, _31875_, _33672_);
  nand _45902_ (_33726_, _29094_, _28008_);
  not _45903_ (_33737_, _28250_);
  and _45904_ (_33748_, _33737_, _28139_);
  not _45905_ (_33759_, _33748_);
  nor _45906_ (_33770_, _33759_, _33726_);
  nand _45907_ (_33781_, _33770_, _32431_);
  or _45908_ (_33791_, _33770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _45909_ (_33802_, _33791_, _32507_);
  and _45910_ (_33813_, _33802_, _33781_);
  or _45911_ (_33824_, _33813_, _33715_);
  or _45912_ (_33835_, _33824_, _33704_);
  and _45913_ (_08900_, _33835_, _43634_);
  and _45914_ (_33856_, _27421_, _24868_);
  not _45915_ (_33867_, _33856_);
  not _45916_ (_33878_, _33552_);
  and _45917_ (_33889_, _33878_, _30201_);
  nor _45918_ (_33899_, _33889_, _30244_);
  nor _45919_ (_33910_, _33899_, _29182_);
  and _45920_ (_33921_, _31471_, _29565_);
  nor _45921_ (_33932_, _31450_, _29554_);
  not _45922_ (_33943_, _33932_);
  and _45923_ (_33954_, _31504_, _29543_);
  and _45924_ (_33965_, _31526_, _22806_);
  nor _45925_ (_33976_, _33965_, _33954_);
  nand _45926_ (_33987_, _33976_, _33943_);
  nor _45927_ (_33998_, _33987_, _33921_);
  nor _45928_ (_34008_, _31570_, _22632_);
  not _45929_ (_34019_, _34008_);
  nor _45930_ (_34030_, _31613_, _22806_);
  nor _45931_ (_34041_, _32648_, _22240_);
  nor _45932_ (_34052_, _34041_, _34030_);
  and _45933_ (_34063_, _34052_, _34019_);
  and _45934_ (_34074_, _34063_, _33998_);
  not _45935_ (_34085_, _34074_);
  nor _45936_ (_34096_, _34085_, _33910_);
  nor _45937_ (_34107_, _30649_, _30627_);
  nor _45938_ (_34117_, _34107_, _31951_);
  and _45939_ (_34128_, _34117_, _30671_);
  nor _45940_ (_34141_, _33257_, _22806_);
  and _45941_ (_34160_, _31232_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45942_ (_34171_, _34160_, _34141_);
  nor _45943_ (_34182_, _34171_, _32027_);
  nor _45944_ (_34193_, _34182_, _34128_);
  and _45945_ (_34204_, _34193_, _34096_);
  and _45946_ (_34215_, _24656_, _19525_);
  not _45947_ (_34226_, _34215_);
  nor _45948_ (_34237_, _31166_, _19922_);
  nor _45949_ (_34247_, _30998_, _30168_);
  nor _45950_ (_34258_, _30889_, _30966_);
  nor _45951_ (_34269_, _34258_, _34247_);
  and _45952_ (_34280_, _34269_, _22816_);
  not _45953_ (_34291_, _34280_);
  not _45954_ (_34302_, _30878_);
  nor _45955_ (_34313_, _34269_, _22816_);
  nor _45956_ (_34324_, _34313_, _34302_);
  and _45957_ (_34335_, _34324_, _34291_);
  nor _45958_ (_34345_, _34335_, _34237_);
  and _45959_ (_34356_, _34345_, _34226_);
  and _45960_ (_34367_, _34356_, _34204_);
  and _45961_ (_34378_, _34367_, _33867_);
  not _45962_ (_34389_, _34378_);
  or _45963_ (_34400_, _34389_, _29105_);
  not _45964_ (_34411_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _45965_ (_34422_, _29105_, _34411_);
  and _45966_ (_34433_, _34422_, _31886_);
  and _45967_ (_34444_, _34433_, _34400_);
  nor _45968_ (_34455_, _31875_, _34411_);
  or _45969_ (_34465_, _32453_, _33726_);
  and _45970_ (_34476_, _34465_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _45971_ (_34487_, _28139_);
  and _45972_ (_34498_, _28008_, _28250_);
  and _45973_ (_34509_, _34498_, _34487_);
  not _45974_ (_34520_, _34509_);
  nor _45975_ (_34531_, _34520_, _32431_);
  and _45976_ (_34542_, _28008_, _28139_);
  and _45977_ (_34553_, _34542_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _45978_ (_34564_, _34553_, _34531_);
  and _45979_ (_34574_, _34564_, _29094_);
  or _45980_ (_34585_, _34574_, _34476_);
  and _45981_ (_34596_, _34585_, _32507_);
  or _45982_ (_34607_, _34596_, _34455_);
  or _45983_ (_34618_, _34607_, _34444_);
  and _45984_ (_08911_, _34618_, _43634_);
  and _45985_ (_34639_, _24698_, _19525_);
  not _45986_ (_34650_, _34639_);
  and _45987_ (_34661_, _27486_, _24868_);
  nor _45988_ (_34672_, _31166_, _20912_);
  and _45989_ (_34682_, _30900_, _30168_);
  and _45990_ (_34693_, _30999_, _30966_);
  nor _45991_ (_34704_, _34693_, _34682_);
  nor _45992_ (_34715_, _34704_, _22240_);
  not _45993_ (_34726_, _34715_);
  and _45994_ (_34737_, _34704_, _22240_);
  nor _45995_ (_34748_, _34737_, _34302_);
  and _45996_ (_34759_, _34748_, _34726_);
  nor _45997_ (_34770_, _34759_, _34672_);
  not _45998_ (_34781_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45999_ (_34791_, _31232_, _34781_);
  nor _46000_ (_34802_, _34791_, _22251_);
  or _46001_ (_34813_, _34802_, _32027_);
  nor _46002_ (_34824_, _34813_, _31243_);
  not _46003_ (_34835_, _34824_);
  nor _46004_ (_34846_, _31450_, _29499_);
  and _46005_ (_34857_, _31471_, _29521_);
  nor _46006_ (_34868_, _34857_, _34846_);
  and _46007_ (_34879_, _31504_, _29510_);
  and _46008_ (_34890_, _31526_, _22240_);
  nor _46009_ (_34900_, _34890_, _34879_);
  nor _46010_ (_34911_, _31613_, _22240_);
  nor _46011_ (_34922_, _31570_, _22806_);
  nor _46012_ (_34933_, _32648_, _21946_);
  or _46013_ (_34944_, _34933_, _34922_);
  nor _46014_ (_34955_, _34944_, _34911_);
  and _46015_ (_34966_, _34955_, _34900_);
  and _46016_ (_34977_, _34966_, _34868_);
  and _46017_ (_34988_, _34977_, _34835_);
  and _46018_ (_34999_, _30671_, _30594_);
  or _46019_ (_35010_, _34999_, _31951_);
  nor _46020_ (_35020_, _35010_, _30682_);
  nor _46021_ (_35031_, _30244_, _29741_);
  nor _46022_ (_35042_, _35031_, _30255_);
  nor _46023_ (_35053_, _35042_, _29182_);
  nor _46024_ (_35064_, _35053_, _35020_);
  and _46025_ (_35075_, _35064_, _34988_);
  and _46026_ (_35086_, _35075_, _34770_);
  not _46027_ (_35097_, _35086_);
  nor _46028_ (_35108_, _35097_, _34661_);
  and _46029_ (_35118_, _35108_, _34650_);
  not _46030_ (_35129_, _35118_);
  or _46031_ (_35140_, _35129_, _29105_);
  not _46032_ (_35151_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _46033_ (_35162_, _29105_, _35151_);
  and _46034_ (_35173_, _35162_, _31886_);
  and _46035_ (_35184_, _35173_, _35140_);
  nor _46036_ (_35195_, _31875_, _35151_);
  and _46037_ (_35206_, _33726_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _46038_ (_35217_, _32453_, _28008_);
  and _46039_ (_35227_, _35217_, _33040_);
  nor _46040_ (_35238_, _34542_, _34498_);
  nor _46041_ (_35249_, _35238_, _35151_);
  or _46042_ (_35260_, _35249_, _35227_);
  and _46043_ (_35271_, _35260_, _29094_);
  or _46044_ (_35282_, _35271_, _35206_);
  and _46045_ (_35293_, _35282_, _32507_);
  or _46046_ (_35304_, _35293_, _35195_);
  or _46047_ (_35315_, _35304_, _35184_);
  and _46048_ (_08922_, _35315_, _43634_);
  and _46049_ (_35336_, _27551_, _24868_);
  not _46050_ (_35346_, _35336_);
  and _46051_ (_35357_, _24730_, _19525_);
  nor _46052_ (_35368_, _30321_, _29478_);
  and _46053_ (_35379_, _30321_, _29478_);
  nor _46054_ (_35390_, _35379_, _35368_);
  and _46055_ (_35401_, _35390_, _29171_);
  not _46056_ (_35412_, _35401_);
  nor _46057_ (_35423_, _30714_, _29478_);
  not _46058_ (_35434_, _35423_);
  nor _46059_ (_35445_, _31951_, _30725_);
  and _46060_ (_35455_, _35445_, _35434_);
  nor _46061_ (_35466_, _30168_, _20085_);
  and _46062_ (_35477_, _30168_, _21957_);
  nor _46063_ (_35488_, _35477_, _35466_);
  nor _46064_ (_35499_, _35488_, _31166_);
  and _46065_ (_35510_, _30911_, _30168_);
  and _46066_ (_35521_, _31021_, _30966_);
  nor _46067_ (_35532_, _35521_, _35510_);
  and _46068_ (_35543_, _35532_, _21946_);
  nor _46069_ (_35554_, _35532_, _21946_);
  nor _46070_ (_35564_, _35554_, _35543_);
  and _46071_ (_35575_, _35564_, _30878_);
  nor _46072_ (_35586_, _35575_, _35499_);
  nor _46073_ (_35597_, _31253_, _21957_);
  not _46074_ (_35608_, _35597_);
  nor _46075_ (_35619_, _31264_, _32027_);
  and _46076_ (_35630_, _35619_, _35608_);
  nor _46077_ (_35641_, _31450_, _29467_);
  and _46078_ (_35652_, _31471_, _29478_);
  nor _46079_ (_35663_, _35652_, _35641_);
  and _46080_ (_35673_, _31504_, _29456_);
  and _46081_ (_35684_, _31526_, _21946_);
  nor _46082_ (_35695_, _35684_, _35673_);
  nor _46083_ (_35706_, _32648_, _21761_);
  not _46084_ (_35717_, _35706_);
  nor _46085_ (_35728_, _31613_, _21946_);
  nor _46086_ (_35739_, _31570_, _22240_);
  nor _46087_ (_35750_, _35739_, _35728_);
  and _46088_ (_35761_, _35750_, _35717_);
  and _46089_ (_35772_, _35761_, _35695_);
  and _46090_ (_35782_, _35772_, _35663_);
  not _46091_ (_35793_, _35782_);
  nor _46092_ (_35804_, _35793_, _35630_);
  and _46093_ (_35815_, _35804_, _35586_);
  not _46094_ (_35826_, _35815_);
  nor _46095_ (_35837_, _35826_, _35455_);
  and _46096_ (_35848_, _35837_, _35412_);
  not _46097_ (_35859_, _35848_);
  nor _46098_ (_35869_, _35859_, _35357_);
  and _46099_ (_35880_, _35869_, _35346_);
  not _46100_ (_35891_, _35880_);
  or _46101_ (_35902_, _35891_, _29105_);
  not _46102_ (_35913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _46103_ (_35924_, _29105_, _35913_);
  and _46104_ (_35935_, _35924_, _31886_);
  and _46105_ (_35946_, _35935_, _35902_);
  nor _46106_ (_35957_, _31875_, _35913_);
  not _46107_ (_35968_, _29094_);
  and _46108_ (_35978_, _28260_, _32442_);
  nor _46109_ (_35989_, _28260_, _32442_);
  nor _46110_ (_36000_, _35989_, _35978_);
  or _46111_ (_36011_, _36000_, _35968_);
  and _46112_ (_36022_, _36011_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _46113_ (_36033_, _35978_, _33040_);
  and _46114_ (_36044_, _35989_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _46115_ (_36055_, _36044_, _36033_);
  and _46116_ (_36066_, _36055_, _29094_);
  or _46117_ (_36077_, _36066_, _36022_);
  and _46118_ (_36088_, _36077_, _32507_);
  or _46119_ (_36098_, _36088_, _35957_);
  or _46120_ (_36109_, _36098_, _35946_);
  and _46121_ (_08933_, _36109_, _43634_);
  and _46122_ (_36130_, _27637_, _24868_);
  not _46123_ (_36141_, _36130_);
  and _46124_ (_36152_, _24772_, _19525_);
  nor _46125_ (_36163_, _30747_, _30725_);
  nor _46126_ (_36174_, _36163_, _30758_);
  and _46127_ (_36185_, _36174_, _30452_);
  not _46128_ (_36196_, _36185_);
  nor _46129_ (_36207_, _30332_, _29445_);
  nor _46130_ (_36217_, _36207_, _30343_);
  nor _46131_ (_36228_, _36217_, _29182_);
  nor _46132_ (_36239_, _30168_, _21074_);
  and _46133_ (_36250_, _30168_, _21772_);
  nor _46134_ (_36261_, _36250_, _36239_);
  nor _46135_ (_36272_, _36261_, _31166_);
  and _46136_ (_36283_, _30922_, _30168_);
  and _46137_ (_36294_, _31022_, _30966_);
  nor _46138_ (_36305_, _36294_, _36283_);
  and _46139_ (_36316_, _36305_, _21761_);
  nor _46140_ (_36327_, _36305_, _21761_);
  or _46141_ (_36338_, _36327_, _34302_);
  nor _46142_ (_36348_, _36338_, _36316_);
  nor _46143_ (_36359_, _36348_, _36272_);
  nor _46144_ (_36370_, _31308_, _31264_);
  and _46145_ (_36381_, _36370_, _21761_);
  nor _46146_ (_36392_, _36370_, _21761_);
  nor _46147_ (_36403_, _36392_, _36381_);
  nor _46148_ (_36414_, _36403_, _32027_);
  nor _46149_ (_36425_, _31613_, _21761_);
  not _46150_ (_36436_, _36425_);
  nor _46151_ (_36447_, _32648_, _20738_);
  nor _46152_ (_36458_, _31570_, _21946_);
  nor _46153_ (_36468_, _36458_, _36447_);
  and _46154_ (_36479_, _36468_, _36436_);
  and _46155_ (_36490_, _31471_, _29313_);
  nor _46156_ (_36501_, _31450_, _29302_);
  not _46157_ (_36512_, _36501_);
  and _46158_ (_36523_, _31504_, _29291_);
  and _46159_ (_36534_, _31526_, _21761_);
  nor _46160_ (_36545_, _36534_, _36523_);
  nand _46161_ (_36556_, _36545_, _36512_);
  nor _46162_ (_36567_, _36556_, _36490_);
  and _46163_ (_36578_, _36567_, _36479_);
  not _46164_ (_36589_, _36578_);
  nor _46165_ (_36599_, _36589_, _36414_);
  and _46166_ (_36610_, _36599_, _36359_);
  not _46167_ (_36621_, _36610_);
  nor _46168_ (_36632_, _36621_, _36228_);
  and _46169_ (_36643_, _36632_, _36196_);
  not _46170_ (_36654_, _36643_);
  nor _46171_ (_36665_, _36654_, _36152_);
  and _46172_ (_36675_, _36665_, _36141_);
  not _46173_ (_36686_, _36675_);
  or _46174_ (_36697_, _36686_, _29105_);
  not _46175_ (_36708_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _46176_ (_36719_, _29105_, _36708_);
  and _46177_ (_36730_, _36719_, _31886_);
  and _46178_ (_36741_, _36730_, _36697_);
  nor _46179_ (_36752_, _31875_, _36708_);
  and _46180_ (_36762_, _33748_, _32442_);
  and _46181_ (_36773_, _36762_, _29094_);
  nand _46182_ (_36784_, _36773_, _32431_);
  or _46183_ (_36795_, _36773_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _46184_ (_36806_, _36795_, _32507_);
  and _46185_ (_36817_, _36806_, _36784_);
  or _46186_ (_36828_, _36817_, _36752_);
  or _46187_ (_36839_, _36828_, _36741_);
  and _46188_ (_08944_, _36839_, _43634_);
  and _46189_ (_36859_, _27702_, _24868_);
  not _46190_ (_36870_, _36859_);
  and _46191_ (_36881_, _24804_, _19525_);
  nor _46192_ (_36892_, _30343_, _29412_);
  nor _46193_ (_36903_, _36892_, _30354_);
  nor _46194_ (_36914_, _36903_, _29182_);
  not _46195_ (_36925_, _36914_);
  nor _46196_ (_36935_, _30168_, _20422_);
  and _46197_ (_36946_, _30168_, _20749_);
  nor _46198_ (_36957_, _36946_, _36935_);
  nor _46199_ (_36968_, _36957_, _31166_);
  or _46200_ (_36979_, _30168_, _21761_);
  or _46201_ (_36990_, _36294_, _30933_);
  and _46202_ (_37001_, _36990_, _36979_);
  nor _46203_ (_37011_, _37001_, _20749_);
  and _46204_ (_37022_, _37001_, _20749_);
  or _46205_ (_37033_, _37022_, _34302_);
  nor _46206_ (_37044_, _37033_, _37011_);
  nor _46207_ (_37055_, _37044_, _36968_);
  nor _46208_ (_37066_, _36381_, _20738_);
  and _46209_ (_37077_, _36381_, _20738_);
  nor _46210_ (_37088_, _37077_, _37066_);
  nor _46211_ (_37098_, _37088_, _32027_);
  nor _46212_ (_37109_, _31613_, _20738_);
  not _46213_ (_37120_, _37109_);
  nor _46214_ (_37131_, _32648_, _21576_);
  nor _46215_ (_37142_, _31570_, _21761_);
  nor _46216_ (_37153_, _37142_, _37131_);
  and _46217_ (_37164_, _37153_, _37120_);
  and _46218_ (_37175_, _31471_, _29258_);
  nor _46219_ (_37185_, _31450_, _29247_);
  not _46220_ (_37196_, _37185_);
  and _46221_ (_37207_, _31504_, _29236_);
  and _46222_ (_37218_, _31526_, _20738_);
  nor _46223_ (_37229_, _37218_, _37207_);
  nand _46224_ (_37240_, _37229_, _37196_);
  nor _46225_ (_37251_, _37240_, _37175_);
  and _46226_ (_37262_, _37251_, _37164_);
  not _46227_ (_37273_, _37262_);
  nor _46228_ (_37284_, _37273_, _37098_);
  and _46229_ (_37294_, _37284_, _37055_);
  not _46230_ (_37305_, _37294_);
  nor _46231_ (_37316_, _30780_, _30758_);
  not _46232_ (_37327_, _37316_);
  nor _46233_ (_37338_, _31951_, _30791_);
  and _46234_ (_37349_, _37338_, _37327_);
  nor _46235_ (_37360_, _37349_, _37305_);
  and _46236_ (_37371_, _37360_, _36925_);
  not _46237_ (_37382_, _37371_);
  nor _46238_ (_37393_, _37382_, _36881_);
  and _46239_ (_37403_, _37393_, _36870_);
  not _46240_ (_37414_, _37403_);
  or _46241_ (_37425_, _37414_, _29105_);
  not _46242_ (_37436_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _46243_ (_37447_, _29105_, _37436_);
  and _46244_ (_37458_, _37447_, _31886_);
  and _46245_ (_37469_, _37458_, _37425_);
  nor _46246_ (_37480_, _31875_, _37436_);
  nor _46247_ (_37491_, _28008_, _28139_);
  and _46248_ (_37502_, _37491_, _28250_);
  and _46249_ (_37513_, _37502_, _29094_);
  nand _46250_ (_37524_, _37513_, _32431_);
  or _46251_ (_37535_, _37513_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _46252_ (_37546_, _37535_, _32507_);
  and _46253_ (_37557_, _37546_, _37524_);
  or _46254_ (_37568_, _37557_, _37480_);
  or _46255_ (_37579_, _37568_, _37469_);
  and _46256_ (_08955_, _37579_, _43634_);
  and _46257_ (_37600_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46258_ (_37611_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _46259_ (_37622_, _37611_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _46260_ (_37633_, _37622_);
  not _46261_ (_37644_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _46262_ (_37654_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _46263_ (_37665_, _37654_, _37644_);
  and _46264_ (_37676_, _37611_, _19459_);
  and _46265_ (_37687_, _37676_, _37665_);
  and _46266_ (_37698_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _46267_ (_37709_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _46268_ (_37720_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _46269_ (_37731_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _46270_ (_37742_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _46271_ (_37753_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _46272_ (_37764_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _46273_ (_37774_, _37764_, _37753_);
  and _46274_ (_37785_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _46275_ (_37796_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _46276_ (_37807_, _37796_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _46277_ (_37818_, _37807_, _37753_);
  and _46278_ (_37829_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _46279_ (_37840_, _37829_, _37785_);
  nor _46280_ (_37851_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _46281_ (_37862_, _37851_, _37753_);
  and _46282_ (_37873_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _46283_ (_37883_, _37851_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _46284_ (_37894_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _46285_ (_37905_, _37894_, _37873_);
  and _46286_ (_37916_, _37851_, _37753_);
  and _46287_ (_37927_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _46288_ (_37938_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _46289_ (_37949_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _37938_);
  and _46290_ (_37960_, _37949_, _37753_);
  and _46291_ (_37971_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _46292_ (_37982_, _37971_, _37927_);
  and _46293_ (_37992_, _37982_, _37905_);
  and _46294_ (_38003_, _37992_, _37840_);
  nor _46295_ (_38014_, _38003_, _37742_);
  and _46296_ (_38025_, _38014_, _37731_);
  or _46297_ (_38036_, _38025_, _37720_);
  and _46298_ (_38047_, _38036_, _37709_);
  nor _46299_ (_38058_, _38047_, _37698_);
  and _46300_ (_38069_, _38058_, _37687_);
  not _46301_ (_38080_, _38069_);
  not _46302_ (_38091_, _37665_);
  nor _46303_ (_38102_, _37676_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _46304_ (_38113_, _38102_, _38091_);
  and _46305_ (_38124_, _38113_, _38080_);
  not _46306_ (_38135_, _37687_);
  and _46307_ (_38146_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _46308_ (_38157_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _46309_ (_38166_, _38157_, _38146_);
  and _46310_ (_38173_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not _46311_ (_38181_, _38173_);
  and _46312_ (_38189_, _38181_, _38166_);
  and _46313_ (_38196_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _46314_ (_38204_, _38196_, _37742_);
  and _46315_ (_38212_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _46316_ (_38219_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _46317_ (_38226_, _38219_, _38212_);
  and _46318_ (_38227_, _38226_, _38204_);
  and _46319_ (_38228_, _38227_, _38189_);
  and _46320_ (_38231_, _38228_, _37731_);
  nor _46321_ (_38238_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _37731_);
  nor _46322_ (_38249_, _38238_, _38231_);
  nor _46323_ (_38260_, _38249_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _46324_ (_38271_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _37709_);
  nor _46325_ (_38282_, _38271_, _38260_);
  nor _46326_ (_38293_, _38282_, _38135_);
  not _46327_ (_38304_, _38293_);
  nor _46328_ (_38315_, _37676_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _46329_ (_38326_, _38315_, _38091_);
  and _46330_ (_38337_, _38326_, _38304_);
  and _46331_ (_38348_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _46332_ (_38359_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _46333_ (_38370_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and _46334_ (_38381_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _46335_ (_38392_, _38381_, _38370_);
  and _46336_ (_38403_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _46337_ (_38414_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _46338_ (_38425_, _38414_, _38403_);
  and _46339_ (_38436_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _46340_ (_38447_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _46341_ (_38458_, _38447_, _38436_);
  and _46342_ (_38469_, _38458_, _38425_);
  and _46343_ (_38480_, _38469_, _38392_);
  nor _46344_ (_38491_, _38480_, _37742_);
  and _46345_ (_38502_, _38491_, _37731_);
  or _46346_ (_38513_, _38502_, _38359_);
  and _46347_ (_38524_, _38513_, _37709_);
  nor _46348_ (_38535_, _38524_, _38348_);
  and _46349_ (_38546_, _38535_, _37687_);
  not _46350_ (_38557_, _38546_);
  nor _46351_ (_38568_, _37676_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _46352_ (_38579_, _38568_, _38091_);
  and _46353_ (_38590_, _38579_, _38557_);
  and _46354_ (_38601_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _46355_ (_38612_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _46356_ (_38623_, _37742_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _46357_ (_38634_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _46358_ (_38645_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _46359_ (_38656_, _38645_, _38634_);
  and _46360_ (_38667_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _46361_ (_38678_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _46362_ (_38689_, _38678_, _38667_);
  and _46363_ (_38700_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _46364_ (_38711_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _46365_ (_38722_, _38711_, _38700_);
  and _46366_ (_38733_, _38722_, _38689_);
  and _46367_ (_38744_, _38733_, _38656_);
  nor _46368_ (_38755_, _38744_, _38623_);
  nor _46369_ (_38766_, _38755_, _38612_);
  nor _46370_ (_38777_, _38766_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _46371_ (_38788_, _38777_, _38601_);
  nor _46372_ (_38799_, _38788_, _38135_);
  and _46373_ (_38810_, _38135_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or _46374_ (_38821_, _38810_, _38799_);
  and _46375_ (_38832_, _38821_, _37665_);
  nor _46376_ (_38843_, _38832_, _38590_);
  and _46377_ (_38854_, _38843_, _38337_);
  and _46378_ (_38865_, _38854_, _38124_);
  and _46379_ (_38876_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _46380_ (_38886_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _46381_ (_38897_, _38886_, _38876_);
  and _46382_ (_38908_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _46383_ (_38918_, _38908_, _37742_);
  and _46384_ (_38929_, _38918_, _38897_);
  and _46385_ (_38940_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _46386_ (_38951_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _46387_ (_38962_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _46388_ (_38973_, _38962_, _38951_);
  nor _46389_ (_38984_, _38973_, _38940_);
  and _46390_ (_38988_, _38984_, _38929_);
  and _46391_ (_38989_, _38988_, _37731_);
  nor _46392_ (_38990_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _37731_);
  or _46393_ (_38991_, _38990_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _46394_ (_38992_, _38991_, _38989_);
  and _46395_ (_38993_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or _46396_ (_38994_, _38993_, _38992_);
  nor _46397_ (_38995_, _38994_, _38135_);
  not _46398_ (_38996_, _38995_);
  nor _46399_ (_38997_, _37676_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _46400_ (_38998_, _38997_, _38091_);
  and _46401_ (_38999_, _38998_, _38996_);
  not _46402_ (_39000_, _38999_);
  and _46403_ (_39001_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _46404_ (_39002_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _46405_ (_39003_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _46406_ (_39004_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _46407_ (_39005_, _39004_, _39003_);
  and _46408_ (_39006_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _46409_ (_39007_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _46410_ (_39008_, _39007_, _39006_);
  and _46411_ (_39009_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _46412_ (_39010_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _46413_ (_39011_, _39010_, _39009_);
  and _46414_ (_39012_, _39011_, _39008_);
  and _46415_ (_39013_, _39012_, _39005_);
  nor _46416_ (_39014_, _39013_, _37742_);
  and _46417_ (_39015_, _39014_, _37731_);
  or _46418_ (_39016_, _39015_, _39002_);
  and _46419_ (_39017_, _39016_, _37709_);
  nor _46420_ (_39018_, _39017_, _39001_);
  and _46421_ (_39019_, _39018_, _37687_);
  not _46422_ (_39020_, _39019_);
  nor _46423_ (_39021_, _37676_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _46424_ (_39022_, _39021_, _38091_);
  and _46425_ (_39023_, _39022_, _39020_);
  and _46426_ (_39024_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and _46427_ (_39025_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _46428_ (_39026_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _46429_ (_39027_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _46430_ (_39028_, _39027_, _39026_);
  and _46431_ (_39029_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _46432_ (_39030_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _46433_ (_39031_, _39030_, _39029_);
  and _46434_ (_39032_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _46435_ (_39033_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _46436_ (_39034_, _39033_, _39032_);
  and _46437_ (_39035_, _39034_, _39031_);
  and _46438_ (_39036_, _39035_, _39028_);
  nor _46439_ (_39037_, _39036_, _37742_);
  and _46440_ (_39038_, _39037_, _37731_);
  or _46441_ (_39039_, _39038_, _39025_);
  and _46442_ (_39040_, _39039_, _37709_);
  nor _46443_ (_39041_, _39040_, _39024_);
  and _46444_ (_39042_, _39041_, _37687_);
  not _46445_ (_39043_, _39042_);
  nor _46446_ (_39044_, _37676_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _46447_ (_39045_, _39044_, _38091_);
  and _46448_ (_39046_, _39045_, _39043_);
  not _46449_ (_39047_, _39046_);
  and _46450_ (_39048_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _46451_ (_39049_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _46452_ (_39050_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _46453_ (_39051_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _46454_ (_39052_, _39051_, _39050_);
  and _46455_ (_39053_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _46456_ (_39054_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _46457_ (_39055_, _39054_, _39053_);
  and _46458_ (_39056_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _46459_ (_39057_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _46460_ (_39058_, _39057_, _39056_);
  and _46461_ (_39059_, _39058_, _39055_);
  and _46462_ (_39060_, _39059_, _39052_);
  nor _46463_ (_39061_, _39060_, _38623_);
  nor _46464_ (_39062_, _39061_, _39049_);
  nor _46465_ (_39063_, _39062_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _46466_ (_39064_, _39063_, _39048_);
  nor _46467_ (_39065_, _39064_, _38135_);
  and _46468_ (_39066_, _38135_, \oc8051_top_1.oc8051_decoder1.op [6]);
  or _46469_ (_39067_, _39066_, _39065_);
  and _46470_ (_39068_, _39067_, _37665_);
  nor _46471_ (_39069_, _39068_, _39047_);
  and _46472_ (_39070_, _39069_, _39023_);
  and _46473_ (_39071_, _39070_, _39000_);
  and _46474_ (_39072_, _39071_, _38865_);
  not _46475_ (_39073_, _39072_);
  not _46476_ (_39074_, _39023_);
  and _46477_ (_39075_, _39069_, _39074_);
  and _46478_ (_39076_, _39075_, _38999_);
  and _46479_ (_39077_, _39076_, _38865_);
  and _46480_ (_39078_, _39068_, _39023_);
  and _46481_ (_39079_, _39078_, _39047_);
  and _46482_ (_39080_, _39079_, _38999_);
  and _46483_ (_39081_, _39080_, _38865_);
  nor _46484_ (_39082_, _39081_, _39077_);
  and _46485_ (_39083_, _39082_, _39073_);
  nor _46486_ (_39084_, _39083_, _37633_);
  not _46487_ (_39085_, _39084_);
  and _46488_ (_39086_, _39068_, _39047_);
  nor _46489_ (_39087_, _38124_, _38337_);
  and _46490_ (_39088_, _39087_, _38843_);
  not _46491_ (_39089_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _46492_ (_39090_, _19459_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _46493_ (_39091_, _39090_, _39089_);
  and _46494_ (_39092_, _39091_, _39088_);
  and _46495_ (_39093_, _39092_, _39086_);
  and _46496_ (_39094_, _39075_, _39000_);
  not _46497_ (_39095_, _38590_);
  and _46498_ (_39096_, _38832_, _39095_);
  and _46499_ (_39097_, _39087_, _39096_);
  and _46500_ (_39098_, _39097_, _39094_);
  and _46501_ (_39099_, _39097_, _39071_);
  nor _46502_ (_39100_, _39099_, _39098_);
  not _46503_ (_39101_, _39100_);
  nor _46504_ (_39102_, _39101_, _39093_);
  and _46505_ (_39103_, _39102_, _39085_);
  nor _46506_ (_39104_, _39103_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46507_ (_39105_, _39104_, _37600_);
  and _46508_ (_39106_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _46509_ (_39107_, _38337_);
  and _46510_ (_39108_, _38124_, _39107_);
  and _46511_ (_39109_, _39108_, _39096_);
  and _46512_ (_39110_, _39068_, _39074_);
  and _46513_ (_39111_, _39110_, _39046_);
  and _46514_ (_39112_, _39111_, _38999_);
  and _46515_ (_39113_, _39112_, _39109_);
  not _46516_ (_39114_, _39113_);
  and _46517_ (_39115_, _39086_, _39074_);
  and _46518_ (_39116_, _39115_, _39000_);
  and _46519_ (_39117_, _39116_, _38854_);
  not _46520_ (_39118_, _38124_);
  and _46521_ (_39119_, _38854_, _39118_);
  and _46522_ (_39120_, _39080_, _39119_);
  nor _46523_ (_39121_, _39120_, _39117_);
  and _46524_ (_39122_, _39121_, _39114_);
  and _46525_ (_39123_, _39111_, _39000_);
  and _46526_ (_39124_, _39123_, _39119_);
  and _46527_ (_39125_, _39070_, _38999_);
  and _46528_ (_39126_, _39125_, _39119_);
  nor _46529_ (_39127_, _39126_, _39124_);
  and _46530_ (_39128_, _39071_, _39088_);
  and _46531_ (_39129_, _39116_, _39109_);
  nor _46532_ (_39130_, _39129_, _39128_);
  nor _46533_ (_39131_, _39068_, _39046_);
  and _46534_ (_39132_, _39131_, _39074_);
  and _46535_ (_39133_, _39132_, _38999_);
  and _46536_ (_39134_, _39133_, _39109_);
  and _46537_ (_39135_, _39088_, _39125_);
  nor _46538_ (_39136_, _39135_, _39134_);
  and _46539_ (_39137_, _39136_, _39130_);
  and _46540_ (_39138_, _39137_, _39127_);
  and _46541_ (_39139_, _39138_, _39122_);
  and _46542_ (_39140_, _39076_, _39119_);
  and _46543_ (_39141_, _39094_, _39109_);
  nor _46544_ (_39142_, _39141_, _39140_);
  and _46545_ (_39143_, _39088_, _39111_);
  and _46546_ (_39144_, _39079_, _39000_);
  and _46547_ (_39145_, _39144_, _38854_);
  nor _46548_ (_39146_, _39145_, _39143_);
  and _46549_ (_39147_, _39146_, _39142_);
  and _46550_ (_39148_, _39094_, _39119_);
  and _46551_ (_39149_, _39115_, _38999_);
  and _46552_ (_39150_, _39149_, _38854_);
  nor _46553_ (_39151_, _39150_, _39148_);
  not _46554_ (_39152_, _39151_);
  not _46555_ (_39153_, _39109_);
  nor _46556_ (_39154_, _39076_, _39125_);
  nor _46557_ (_39155_, _39154_, _39153_);
  nor _46558_ (_39156_, _39155_, _39152_);
  and _46559_ (_39157_, _39156_, _39147_);
  and _46560_ (_39158_, _39131_, _39023_);
  nor _46561_ (_39159_, _39158_, _39149_);
  nor _46562_ (_39160_, _39159_, _39153_);
  not _46563_ (_39161_, _39160_);
  and _46564_ (_39162_, _39132_, _39000_);
  and _46565_ (_39163_, _39162_, _39109_);
  and _46566_ (_39164_, _39158_, _39119_);
  nor _46567_ (_39165_, _39164_, _39163_);
  and _46568_ (_39166_, _39165_, _39161_);
  and _46569_ (_39167_, _39144_, _39109_);
  and _46570_ (_39168_, _39123_, _39109_);
  nor _46571_ (_39169_, _39168_, _39167_);
  and _46572_ (_39170_, _39119_, _39112_);
  and _46573_ (_39171_, _39071_, _39119_);
  nor _46574_ (_39172_, _39171_, _39170_);
  and _46575_ (_39173_, _39172_, _39169_);
  and _46576_ (_39174_, _39173_, _39166_);
  and _46577_ (_39175_, _39158_, _38999_);
  and _46578_ (_39176_, _39175_, _39088_);
  not _46579_ (_39177_, _39176_);
  and _46580_ (_39178_, _39158_, _39000_);
  and _46581_ (_39179_, _39178_, _39088_);
  and _46582_ (_39180_, _39133_, _39088_);
  nor _46583_ (_39181_, _39180_, _39179_);
  and _46584_ (_39182_, _39181_, _39177_);
  and _46585_ (_39183_, _38337_, _38832_);
  and _46586_ (_39184_, _39183_, _39095_);
  and _46587_ (_39185_, _39184_, _39000_);
  and _46588_ (_39186_, _39185_, _39070_);
  not _46589_ (_39187_, _39186_);
  and _46590_ (_39188_, _39078_, _39046_);
  and _46591_ (_39189_, _39188_, _39000_);
  and _46592_ (_39190_, _39189_, _39109_);
  and _46593_ (_39191_, _39071_, _38590_);
  nor _46594_ (_39192_, _39191_, _39190_);
  and _46595_ (_39193_, _39192_, _39187_);
  and _46596_ (_39194_, _39193_, _39182_);
  and _46597_ (_39195_, _39194_, _39174_);
  and _46598_ (_39196_, _39195_, _39157_);
  and _46599_ (_39197_, _39196_, _39139_);
  nor _46600_ (_39198_, _39197_, _37633_);
  and _46601_ (_39199_, \oc8051_top_1.oc8051_decoder1.state [0], _19459_);
  and _46602_ (_39200_, _39199_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _46603_ (_39201_, _39200_, _39164_);
  or _46604_ (_39202_, _39093_, _39201_);
  nor _46605_ (_39203_, _39202_, _39198_);
  nor _46606_ (_39204_, _39203_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46607_ (_39205_, _39204_, _39106_);
  and _46608_ (_39206_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _46609_ (_39207_, _39184_);
  nor _46610_ (_39208_, _39207_, _39159_);
  and _46611_ (_39209_, _39184_, _39111_);
  nor _46612_ (_39210_, _39000_, _38590_);
  and _46613_ (_39211_, _39210_, _39183_);
  and _46614_ (_39212_, _39211_, _39075_);
  or _46615_ (_39213_, _39212_, _39209_);
  and _46616_ (_39214_, _39184_, _39132_);
  and _46617_ (_39215_, _39211_, _39070_);
  or _46618_ (_39216_, _39215_, _39214_);
  or _46619_ (_39217_, _39216_, _39213_);
  or _46620_ (_39218_, _39217_, _39208_);
  and _46621_ (_39219_, _39188_, _39185_);
  and _46622_ (_39220_, _39185_, _39110_);
  and _46623_ (_39221_, _39220_, _39047_);
  or _46624_ (_39222_, _39221_, _39219_);
  and _46625_ (_39223_, _39088_, _39112_);
  and _46626_ (_39224_, _39185_, _39075_);
  or _46627_ (_39225_, _39224_, _39223_);
  and _46628_ (_39226_, _39184_, _39144_);
  or _46629_ (_39227_, _39226_, _39164_);
  or _46630_ (_39228_, _39227_, _39225_);
  or _46631_ (_39229_, _39228_, _39222_);
  or _46632_ (_39230_, _39229_, _39218_);
  and _46633_ (_39231_, _39230_, _37622_);
  and _46634_ (_39232_, _39093_, _39023_);
  or _46635_ (_39233_, _39232_, _39201_);
  or _46636_ (_39234_, _39233_, _39084_);
  or _46637_ (_39235_, _39234_, _39231_);
  and _46638_ (_39236_, _39235_, _19459_);
  nor _46639_ (_39237_, _39236_, _39206_);
  nor _46640_ (_39238_, _39237_, _39205_);
  and _46641_ (_39239_, _39238_, _39105_);
  and _46642_ (_09506_, _39239_, _43634_);
  and _46643_ (_39240_, _29061_, _28611_);
  and _46644_ (_39241_, _28490_, _28776_);
  and _46645_ (_39242_, _39241_, _39240_);
  and _46646_ (_39243_, _39242_, _33748_);
  and _46647_ (_39244_, _31886_, _28918_);
  and _46648_ (_39245_, _39244_, _28008_);
  and _46649_ (_39246_, _39245_, _39243_);
  not _46650_ (_39247_, _39246_);
  and _46651_ (_39248_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _46652_ (_39249_, _39243_, _28008_);
  and _46653_ (_39250_, _39249_, _39244_);
  not _46654_ (_39251_, _39250_);
  nor _46655_ (_39252_, _24868_, _19525_);
  and _46656_ (_39253_, _30441_, _24846_);
  nor _46657_ (_39254_, _31602_, _39253_);
  and _46658_ (_39255_, _39254_, _39252_);
  nor _46659_ (_39256_, _32637_, _31559_);
  and _46660_ (_39257_, _39256_, _39255_);
  nor _46661_ (_39258_, _39257_, _20738_);
  not _46662_ (_39259_, _39258_);
  and _46663_ (_39260_, _39259_, _37251_);
  and _46664_ (_39261_, _39260_, _37055_);
  nor _46665_ (_39262_, _39261_, _39251_);
  nor _46666_ (_39263_, _39262_, _39248_);
  and _46667_ (_39264_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _46668_ (_39265_, _39257_, _21761_);
  not _46669_ (_39266_, _39265_);
  and _46670_ (_39267_, _39266_, _36567_);
  and _46671_ (_39268_, _39267_, _36359_);
  nor _46672_ (_39269_, _39268_, _39251_);
  nor _46673_ (_39270_, _39269_, _39264_);
  and _46674_ (_39271_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _46675_ (_39272_, _39257_, _21946_);
  not _46676_ (_39273_, _39272_);
  and _46677_ (_39274_, _39273_, _35695_);
  and _46678_ (_39275_, _39274_, _35663_);
  and _46679_ (_39276_, _39275_, _35586_);
  nor _46680_ (_39277_, _39276_, _39251_);
  nor _46681_ (_39278_, _39277_, _39271_);
  and _46682_ (_39279_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _46683_ (_39280_, _39257_, _22240_);
  not _46684_ (_39281_, _39280_);
  and _46685_ (_39282_, _39281_, _34900_);
  and _46686_ (_39283_, _39282_, _34868_);
  and _46687_ (_39284_, _39283_, _34770_);
  nor _46688_ (_39285_, _39284_, _39251_);
  nor _46689_ (_39286_, _39285_, _39279_);
  and _46690_ (_39287_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _46691_ (_39288_, _39257_, _22806_);
  not _46692_ (_39289_, _39288_);
  and _46693_ (_39290_, _39289_, _33998_);
  and _46694_ (_39291_, _39290_, _34345_);
  nor _46695_ (_39292_, _39291_, _39251_);
  nor _46696_ (_39293_, _39292_, _39287_);
  and _46697_ (_39294_, _39247_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _46698_ (_39295_, _39257_, _22632_);
  not _46699_ (_39296_, _39295_);
  and _46700_ (_39297_, _39296_, _33366_);
  and _46701_ (_39298_, _39297_, _33225_);
  nor _46702_ (_39299_, _39298_, _39247_);
  nor _46703_ (_39300_, _39299_, _39294_);
  nor _46704_ (_39301_, _39246_, _28195_);
  nor _46705_ (_39302_, _39257_, _23175_);
  not _46706_ (_39303_, _39302_);
  and _46707_ (_39304_, _39303_, _32735_);
  and _46708_ (_39305_, _39304_, _32899_);
  and _46709_ (_39306_, _39305_, _32626_);
  not _46710_ (_39307_, _39306_);
  and _46711_ (_39308_, _39307_, _39250_);
  nor _46712_ (_39309_, _39308_, _39301_);
  and _46713_ (_39310_, _39309_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46714_ (_39311_, _39310_, _39300_);
  and _46715_ (_39312_, _39311_, _39293_);
  and _46716_ (_39313_, _39312_, _39286_);
  and _46717_ (_39314_, _39313_, _39278_);
  and _46718_ (_39315_, _39314_, _39270_);
  and _46719_ (_39316_, _39315_, _39263_);
  nor _46720_ (_39317_, _39246_, _28633_);
  nand _46721_ (_39318_, _39317_, _39316_);
  or _46722_ (_39319_, _39317_, _39316_);
  and _46723_ (_39320_, _39319_, _28337_);
  and _46724_ (_39321_, _39320_, _39318_);
  or _46725_ (_39322_, _39246_, _28677_);
  or _46726_ (_39323_, _39322_, _39321_);
  or _46727_ (_39324_, _39257_, _21576_);
  and _46728_ (_39325_, _39324_, _31548_);
  and _46729_ (_39326_, _39325_, _31493_);
  and _46730_ (_39327_, _39326_, _31199_);
  nand _46731_ (_39328_, _39327_, _39246_);
  and _46732_ (_39329_, _39328_, _39323_);
  and _46733_ (_09527_, _39329_, _43634_);
  not _46734_ (_39330_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46735_ (_39331_, _39309_, _39330_);
  nor _46736_ (_39332_, _39309_, _39330_);
  nor _46737_ (_39333_, _39332_, _39331_);
  and _46738_ (_39334_, _39333_, _28337_);
  nor _46739_ (_39335_, _39334_, _28206_);
  nor _46740_ (_39336_, _39335_, _39250_);
  nor _46741_ (_39337_, _39336_, _39308_);
  nand _46742_ (_10682_, _39337_, _43634_);
  nor _46743_ (_39338_, _39310_, _39300_);
  nor _46744_ (_39339_, _39338_, _39311_);
  nor _46745_ (_39340_, _39339_, _27756_);
  nor _46746_ (_39341_, _39340_, _28041_);
  nor _46747_ (_39342_, _39341_, _39250_);
  nor _46748_ (_39343_, _39342_, _39299_);
  nand _46749_ (_10693_, _39343_, _43634_);
  nor _46750_ (_39344_, _39311_, _39293_);
  nor _46751_ (_39345_, _39344_, _39312_);
  nor _46752_ (_39346_, _39345_, _27756_);
  nor _46753_ (_39347_, _39346_, _27811_);
  nor _46754_ (_39348_, _39347_, _39250_);
  nor _46755_ (_39349_, _39348_, _39292_);
  nand _46756_ (_10704_, _39349_, _43634_);
  nor _46757_ (_39350_, _39312_, _39286_);
  nor _46758_ (_39351_, _39350_, _39313_);
  nor _46759_ (_39352_, _39351_, _27756_);
  nor _46760_ (_39353_, _39352_, _28863_);
  nor _46761_ (_39354_, _39353_, _39250_);
  nor _46762_ (_39355_, _39354_, _39285_);
  nor _46763_ (_10715_, _39355_, rst);
  nor _46764_ (_39356_, _39313_, _39278_);
  nor _46765_ (_39357_, _39356_, _39314_);
  nor _46766_ (_39358_, _39357_, _27756_);
  nor _46767_ (_39359_, _39358_, _28984_);
  nor _46768_ (_39360_, _39359_, _39250_);
  nor _46769_ (_39361_, _39360_, _39277_);
  nor _46770_ (_10726_, _39361_, rst);
  nor _46771_ (_39362_, _39314_, _39270_);
  nor _46772_ (_39363_, _39362_, _39315_);
  nor _46773_ (_39364_, _39363_, _27756_);
  nor _46774_ (_39365_, _39364_, _28524_);
  nor _46775_ (_39366_, _39365_, _39250_);
  nor _46776_ (_39367_, _39366_, _39269_);
  nor _46777_ (_10737_, _39367_, rst);
  nor _46778_ (_39368_, _39315_, _39263_);
  nor _46779_ (_39369_, _39368_, _39316_);
  nor _46780_ (_39370_, _39369_, _27756_);
  nor _46781_ (_39371_, _39370_, _28370_);
  nor _46782_ (_39372_, _39371_, _39250_);
  nor _46783_ (_39373_, _39372_, _39262_);
  nor _46784_ (_10748_, _39373_, rst);
  and _46785_ (_39374_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _19459_);
  and _46786_ (_39375_, _39374_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not _46787_ (_39376_, _39375_);
  nor _46788_ (_39377_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _46789_ (_39378_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46790_ (_39379_, _39378_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46791_ (_39380_, _39379_, _39377_);
  nor _46792_ (_39381_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _46793_ (_39382_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46794_ (_39383_, _39382_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46795_ (_39384_, _39383_, _39381_);
  nor _46796_ (_39385_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _46797_ (_39386_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46798_ (_39387_, _39386_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46799_ (_39388_, _39387_, _39385_);
  not _46800_ (_39389_, _39388_);
  nor _46801_ (_39390_, _39389_, _31962_);
  nor _46802_ (_39391_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _46803_ (_39392_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46804_ (_39393_, _39392_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46805_ (_39394_, _39393_, _39391_);
  and _46806_ (_39395_, _39394_, _39390_);
  nor _46807_ (_39396_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _46808_ (_39397_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46809_ (_39398_, _39397_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46810_ (_39399_, _39398_, _39396_);
  and _46811_ (_39400_, _39399_, _39395_);
  and _46812_ (_39401_, _39400_, _39384_);
  nor _46813_ (_39402_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _46814_ (_39403_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46815_ (_39404_, _39403_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46816_ (_39405_, _39404_, _39402_);
  and _46817_ (_39406_, _39405_, _39401_);
  and _46818_ (_39407_, _39406_, _39380_);
  nor _46819_ (_39408_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _46820_ (_39409_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46821_ (_39410_, _39409_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46822_ (_39411_, _39410_, _39408_);
  and _46823_ (_39412_, _39411_, _39407_);
  nor _46824_ (_39413_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _46825_ (_39414_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _46826_ (_39415_, _39414_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46827_ (_39416_, _39415_, _39413_);
  nor _46828_ (_39417_, _39416_, _39412_);
  and _46829_ (_39418_, _39416_, _39412_);
  or _46830_ (_39419_, _39418_, _39417_);
  nor _46831_ (_39420_, _39419_, _31951_);
  not _46832_ (_39421_, _39420_);
  and _46833_ (_39422_, _24561_, _19525_);
  and _46834_ (_39423_, _30944_, _21587_);
  and _46835_ (_39424_, _39423_, _29609_);
  and _46836_ (_39425_, _39424_, _29642_);
  and _46837_ (_39426_, _39425_, _29686_);
  and _46838_ (_39427_, _39426_, _30266_);
  nor _46839_ (_39428_, _39427_, _30966_);
  and _46840_ (_39429_, _30168_, _20085_);
  nor _46841_ (_39430_, _39429_, _39428_);
  and _46842_ (_39431_, _31044_, _21576_);
  and _46843_ (_39432_, _20912_, _19922_);
  and _46844_ (_39433_, _21227_, _20248_);
  and _46845_ (_39434_, _39433_, _39432_);
  and _46846_ (_39435_, _39434_, _39431_);
  and _46847_ (_39436_, _39435_, _20085_);
  and _46848_ (_39437_, _39436_, _21074_);
  nor _46849_ (_39438_, _39437_, _30168_);
  and _46850_ (_39439_, _30168_, _21074_);
  nor _46851_ (_39440_, _39439_, _39438_);
  and _46852_ (_39441_, _39440_, _39430_);
  and _46853_ (_39442_, _30168_, _20422_);
  nor _46854_ (_39443_, _39442_, _36935_);
  and _46855_ (_39444_, _39443_, _39441_);
  nor _46856_ (_39445_, _39444_, _31112_);
  and _46857_ (_39446_, _39444_, _31112_);
  nor _46858_ (_39447_, _39446_, _39445_);
  and _46859_ (_39448_, _39447_, _30878_);
  and _46860_ (_39449_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _46861_ (_39450_, _30168_, _21576_);
  and _46862_ (_39451_, _30168_, _31112_);
  nor _46863_ (_39452_, _39451_, _39450_);
  nor _46864_ (_39453_, _39452_, _31166_);
  nor _46865_ (_39454_, _32289_, _22240_);
  nor _46866_ (_39455_, _31613_, _21402_);
  or _46867_ (_39456_, _39455_, _39454_);
  or _46868_ (_39457_, _39456_, _39453_);
  nor _46869_ (_39458_, _39457_, _39449_);
  not _46870_ (_39459_, _39458_);
  nor _46871_ (_39460_, _39459_, _39448_);
  not _46872_ (_39461_, _39460_);
  nor _46873_ (_39462_, _39461_, _39422_);
  and _46874_ (_39463_, _39462_, _39421_);
  nor _46875_ (_39464_, _39463_, _39376_);
  and _46876_ (_39465_, _39242_, _35217_);
  and _46877_ (_39466_, _39465_, _39244_);
  nand _46878_ (_39467_, _39466_, _31809_);
  or _46879_ (_39468_, _39466_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _46880_ (_39469_, _39468_, _39376_);
  and _46881_ (_39470_, _39469_, _39467_);
  or _46882_ (_39471_, _39470_, _39464_);
  and _46883_ (_12699_, _39471_, _43634_);
  and _46884_ (_39472_, _39242_, _34509_);
  and _46885_ (_39473_, _39472_, _39244_);
  nor _46886_ (_39474_, _39473_, _39375_);
  not _46887_ (_39475_, _39474_);
  nand _46888_ (_39476_, _39475_, _31809_);
  or _46889_ (_39477_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _46890_ (_39478_, _39477_, _43634_);
  and _46891_ (_12720_, _39478_, _39476_);
  not _46892_ (_39479_, _39466_);
  nor _46893_ (_39480_, _39479_, _32953_);
  and _46894_ (_39481_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _46895_ (_39482_, _39481_, _39375_);
  or _46896_ (_39483_, _39482_, _39480_);
  and _46897_ (_39484_, _27166_, _24868_);
  not _46898_ (_39485_, _39484_);
  and _46899_ (_39486_, _39389_, _31962_);
  nor _46900_ (_39487_, _39486_, _39390_);
  and _46901_ (_39488_, _39487_, _30452_);
  nor _46902_ (_39489_, _39450_, _31144_);
  not _46903_ (_39490_, _39489_);
  nor _46904_ (_39491_, _39490_, _31067_);
  nor _46905_ (_39492_, _39491_, _29609_);
  and _46906_ (_39493_, _39491_, _29609_);
  nor _46907_ (_39494_, _39493_, _39492_);
  and _46908_ (_39495_, _39494_, _30878_);
  nor _46909_ (_39496_, _31613_, _20248_);
  and _46910_ (_39497_, _24340_, _19525_);
  nor _46911_ (_39498_, _32289_, _21946_);
  nor _46912_ (_39499_, _31166_, _23175_);
  or _46913_ (_39500_, _39499_, _39498_);
  or _46914_ (_39501_, _39500_, _39497_);
  nor _46915_ (_39502_, _39501_, _39496_);
  not _46916_ (_39503_, _39502_);
  nor _46917_ (_39504_, _39503_, _39495_);
  not _46918_ (_39505_, _39504_);
  nor _46919_ (_39506_, _39505_, _39488_);
  and _46920_ (_39507_, _39506_, _39485_);
  nand _46921_ (_39508_, _39507_, _39375_);
  and _46922_ (_39509_, _39508_, _43634_);
  and _46923_ (_13637_, _39509_, _39483_);
  nor _46924_ (_39510_, _39479_, _33639_);
  and _46925_ (_39511_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _46926_ (_39512_, _39511_, _39375_);
  or _46927_ (_39513_, _39512_, _39510_);
  nor _46928_ (_39514_, _39394_, _39390_);
  not _46929_ (_39515_, _39514_);
  nor _46930_ (_39516_, _39395_, _31951_);
  and _46931_ (_39517_, _39516_, _39515_);
  not _46932_ (_39518_, _39517_);
  and _46933_ (_39519_, _26158_, _24868_);
  nor _46934_ (_39520_, _39424_, _30966_);
  and _46935_ (_39521_, _39431_, _20248_);
  nor _46936_ (_39522_, _39521_, _30168_);
  or _46937_ (_39523_, _39522_, _39520_);
  nor _46938_ (_39524_, _39523_, _29642_);
  and _46939_ (_39525_, _39523_, _29642_);
  or _46940_ (_39526_, _39525_, _39524_);
  and _46941_ (_39527_, _39526_, _30878_);
  nor _46942_ (_39528_, _31613_, _21227_);
  and _46943_ (_39529_, _24371_, _19525_);
  nor _46944_ (_39530_, _32289_, _21761_);
  nor _46945_ (_39531_, _31166_, _22632_);
  or _46946_ (_39532_, _39531_, _39530_);
  or _46947_ (_39533_, _39532_, _39529_);
  nor _46948_ (_39534_, _39533_, _39528_);
  not _46949_ (_39535_, _39534_);
  nor _46950_ (_39536_, _39535_, _39527_);
  not _46951_ (_39537_, _39536_);
  nor _46952_ (_39538_, _39537_, _39519_);
  and _46953_ (_39539_, _39538_, _39518_);
  nand _46954_ (_39540_, _39539_, _39375_);
  and _46955_ (_39541_, _39540_, _43634_);
  and _46956_ (_13648_, _39541_, _39513_);
  nor _46957_ (_39542_, _39479_, _34378_);
  and _46958_ (_39543_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _46959_ (_39544_, _39543_, _39375_);
  or _46960_ (_39545_, _39544_, _39542_);
  nor _46961_ (_39546_, _39399_, _39395_);
  nor _46962_ (_39547_, _39546_, _39400_);
  and _46963_ (_39548_, _39547_, _30452_);
  not _46964_ (_39549_, _39548_);
  and _46965_ (_39550_, _39521_, _21227_);
  and _46966_ (_39551_, _39550_, _30966_);
  and _46967_ (_39552_, _39425_, _30168_);
  nor _46968_ (_39553_, _39552_, _39551_);
  and _46969_ (_39554_, _39553_, _19922_);
  nor _46970_ (_39555_, _39553_, _19922_);
  nor _46971_ (_39556_, _39555_, _39554_);
  and _46972_ (_39557_, _39556_, _30878_);
  not _46973_ (_39558_, _39557_);
  nor _46974_ (_39559_, _31166_, _22806_);
  and _46975_ (_39560_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _46976_ (_39561_, _39560_, _39559_);
  and _46977_ (_39562_, _24403_, _19525_);
  nor _46978_ (_39563_, _32289_, _20738_);
  nor _46979_ (_39564_, _31613_, _19922_);
  or _46980_ (_39565_, _39564_, _39563_);
  nor _46981_ (_39566_, _39565_, _39562_);
  and _46982_ (_39567_, _39566_, _39561_);
  and _46983_ (_39568_, _39567_, _39558_);
  and _46984_ (_39569_, _39568_, _39549_);
  nand _46985_ (_39570_, _39569_, _39375_);
  and _46986_ (_39571_, _39570_, _43634_);
  and _46987_ (_13659_, _39571_, _39545_);
  nor _46988_ (_39572_, _39479_, _35118_);
  and _46989_ (_39573_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _46990_ (_39574_, _39573_, _39375_);
  or _46991_ (_39575_, _39574_, _39572_);
  nor _46992_ (_39576_, _39400_, _39384_);
  nor _46993_ (_39577_, _39576_, _39401_);
  and _46994_ (_39578_, _39577_, _30452_);
  not _46995_ (_39579_, _39578_);
  and _46996_ (_39580_, _24434_, _19525_);
  not _46997_ (_39581_, _39580_);
  nor _46998_ (_39582_, _39426_, _30266_);
  not _46999_ (_39583_, _39582_);
  and _47000_ (_39584_, _39583_, _39428_);
  and _47001_ (_39585_, _39550_, _19922_);
  nor _47002_ (_39586_, _39585_, _20912_);
  nor _47003_ (_39587_, _39586_, _39435_);
  nor _47004_ (_39588_, _39587_, _30168_);
  nor _47005_ (_39589_, _39588_, _39584_);
  nor _47006_ (_39590_, _39589_, _34302_);
  nor _47007_ (_39591_, _31613_, _20912_);
  nor _47008_ (_39592_, _31166_, _22240_);
  and _47009_ (_39593_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _47010_ (_39594_, _39593_, _39592_);
  or _47011_ (_39595_, _39594_, _32300_);
  nor _47012_ (_39596_, _39595_, _39591_);
  not _47013_ (_39597_, _39596_);
  nor _47014_ (_39598_, _39597_, _39590_);
  and _47015_ (_39599_, _39598_, _39581_);
  and _47016_ (_39600_, _39599_, _39579_);
  nand _47017_ (_39601_, _39600_, _39375_);
  and _47018_ (_39602_, _39601_, _43634_);
  and _47019_ (_13670_, _39602_, _39575_);
  nor _47020_ (_39603_, _39479_, _35880_);
  and _47021_ (_39604_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _47022_ (_39605_, _39604_, _39375_);
  or _47023_ (_39606_, _39605_, _39603_);
  nor _47024_ (_39607_, _39405_, _39401_);
  nor _47025_ (_39608_, _39607_, _39406_);
  and _47026_ (_39609_, _39608_, _30452_);
  not _47027_ (_39610_, _39609_);
  and _47028_ (_39611_, _24466_, _19525_);
  nor _47029_ (_39612_, _39435_, _30168_);
  nor _47030_ (_39613_, _39612_, _39428_);
  nor _47031_ (_39614_, _39613_, _29324_);
  and _47032_ (_39615_, _39613_, _29324_);
  nor _47033_ (_39616_, _39615_, _39614_);
  and _47034_ (_39617_, _39616_, _30878_);
  and _47035_ (_39618_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _47036_ (_39619_, _30168_, _21957_);
  or _47037_ (_39620_, _39619_, _31166_);
  nor _47038_ (_39621_, _39620_, _39429_);
  nor _47039_ (_39622_, _32289_, _23175_);
  nor _47040_ (_39623_, _31613_, _20085_);
  or _47041_ (_39624_, _39623_, _39622_);
  or _47042_ (_39625_, _39624_, _39621_);
  nor _47043_ (_39626_, _39625_, _39618_);
  not _47044_ (_39627_, _39626_);
  nor _47045_ (_39628_, _39627_, _39617_);
  not _47046_ (_39629_, _39628_);
  nor _47047_ (_39630_, _39629_, _39611_);
  and _47048_ (_39631_, _39630_, _39610_);
  nand _47049_ (_39632_, _39631_, _39375_);
  and _47050_ (_39633_, _39632_, _43634_);
  and _47051_ (_13681_, _39633_, _39606_);
  nor _47052_ (_39634_, _39479_, _36675_);
  and _47053_ (_39635_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _47054_ (_39636_, _39635_, _39375_);
  or _47055_ (_39637_, _39636_, _39634_);
  nor _47056_ (_39638_, _39406_, _39380_);
  not _47057_ (_39639_, _39638_);
  nor _47058_ (_39640_, _39407_, _31951_);
  and _47059_ (_39641_, _39640_, _39639_);
  not _47060_ (_39642_, _39641_);
  and _47061_ (_39643_, _24498_, _19525_);
  nor _47062_ (_39644_, _39436_, _30168_);
  not _47063_ (_39645_, _39644_);
  and _47064_ (_39646_, _39645_, _39430_);
  and _47065_ (_39647_, _39646_, _21074_);
  nor _47066_ (_39648_, _39646_, _21074_);
  nor _47067_ (_39649_, _39648_, _39647_);
  nor _47068_ (_39650_, _39649_, _34302_);
  and _47069_ (_39651_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _47070_ (_39652_, _30168_, _21772_);
  or _47071_ (_39653_, _39652_, _31166_);
  nor _47072_ (_39654_, _39653_, _39439_);
  nor _47073_ (_39655_, _32289_, _22632_);
  nor _47074_ (_39656_, _31613_, _21074_);
  or _47075_ (_39657_, _39656_, _39655_);
  or _47076_ (_39658_, _39657_, _39654_);
  nor _47077_ (_39659_, _39658_, _39651_);
  not _47078_ (_39660_, _39659_);
  nor _47079_ (_39661_, _39660_, _39650_);
  not _47080_ (_39662_, _39661_);
  nor _47081_ (_39663_, _39662_, _39643_);
  and _47082_ (_39664_, _39663_, _39642_);
  nand _47083_ (_39665_, _39664_, _39375_);
  and _47084_ (_39666_, _39665_, _43634_);
  and _47085_ (_13691_, _39666_, _39637_);
  nor _47086_ (_39667_, _39479_, _37403_);
  and _47087_ (_39668_, _39479_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _47088_ (_39669_, _39668_, _39375_);
  or _47089_ (_39670_, _39669_, _39667_);
  nor _47090_ (_39671_, _39411_, _39407_);
  nor _47091_ (_39672_, _39671_, _39412_);
  and _47092_ (_39673_, _39672_, _30452_);
  not _47093_ (_39674_, _39673_);
  and _47094_ (_39675_, _24529_, _19525_);
  and _47095_ (_39676_, _39441_, _20422_);
  nor _47096_ (_39677_, _39441_, _20422_);
  nor _47097_ (_39678_, _39677_, _39676_);
  nor _47098_ (_39679_, _39678_, _34302_);
  and _47099_ (_39680_, _24868_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _47100_ (_39681_, _30168_, _20749_);
  or _47101_ (_39682_, _39681_, _31166_);
  nor _47102_ (_39683_, _39682_, _39442_);
  nor _47103_ (_39684_, _32289_, _22806_);
  nor _47104_ (_39685_, _31613_, _20422_);
  or _47105_ (_39686_, _39685_, _39684_);
  or _47106_ (_39687_, _39686_, _39683_);
  nor _47107_ (_39688_, _39687_, _39680_);
  not _47108_ (_39689_, _39688_);
  nor _47109_ (_39690_, _39689_, _39679_);
  not _47110_ (_39691_, _39690_);
  nor _47111_ (_39692_, _39691_, _39675_);
  and _47112_ (_39693_, _39692_, _39674_);
  nand _47113_ (_39694_, _39693_, _39375_);
  and _47114_ (_39697_, _39694_, _43634_);
  and _47115_ (_13702_, _39697_, _39670_);
  nand _47116_ (_39699_, _39475_, _32953_);
  or _47117_ (_39700_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _47118_ (_39701_, _39700_, _43634_);
  and _47119_ (_13713_, _39701_, _39699_);
  nand _47120_ (_39702_, _39475_, _33639_);
  or _47121_ (_39703_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _47122_ (_39704_, _39703_, _43634_);
  and _47123_ (_13724_, _39704_, _39702_);
  nand _47124_ (_39705_, _39475_, _34378_);
  or _47125_ (_39707_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _47126_ (_39716_, _39707_, _43634_);
  and _47127_ (_13735_, _39716_, _39705_);
  nand _47128_ (_39727_, _39475_, _35118_);
  or _47129_ (_39730_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _47130_ (_39731_, _39730_, _43634_);
  and _47131_ (_13746_, _39731_, _39727_);
  nand _47132_ (_39732_, _39475_, _35880_);
  or _47133_ (_39733_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _47134_ (_39734_, _39733_, _43634_);
  and _47135_ (_13757_, _39734_, _39732_);
  nand _47136_ (_39735_, _39475_, _36675_);
  or _47137_ (_39736_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _47138_ (_39737_, _39736_, _43634_);
  and _47139_ (_13768_, _39737_, _39735_);
  nand _47140_ (_39738_, _39475_, _37403_);
  or _47141_ (_39739_, _39475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _47142_ (_39740_, _39739_, _43634_);
  and _47143_ (_13779_, _39740_, _39738_);
  not _47144_ (_39741_, _28611_);
  nor _47145_ (_39742_, _39741_, _28490_);
  and _47146_ (_39743_, _39742_, _32507_);
  and _47147_ (_39744_, _39743_, _29083_);
  not _47148_ (_39745_, _32463_);
  nor _47149_ (_39746_, _39745_, _32431_);
  not _47150_ (_39747_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _47151_ (_39748_, _32463_, _39747_);
  or _47152_ (_39749_, _39748_, _39746_);
  and _47153_ (_39750_, _39749_, _39744_);
  nor _47154_ (_39753_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _47155_ (_39754_, _39753_);
  nand _47156_ (_39755_, _39754_, _32431_);
  and _47157_ (_39756_, _39753_, _39747_);
  nor _47158_ (_39757_, _39756_, _39744_);
  and _47159_ (_39758_, _39757_, _39755_);
  nor _47160_ (_39759_, _29061_, _39741_);
  nor _47161_ (_39760_, _28490_, _28765_);
  and _47162_ (_39761_, _39244_, _28271_);
  and _47163_ (_39762_, _39761_, _39760_);
  and _47164_ (_39763_, _39762_, _39759_);
  or _47165_ (_39764_, _39763_, _39758_);
  or _47166_ (_39765_, _39764_, _39750_);
  nand _47167_ (_39766_, _39763_, _39327_);
  and _47168_ (_39767_, _39766_, _43634_);
  and _47169_ (_15177_, _39767_, _39765_);
  and _47170_ (_39768_, _33748_, _28008_);
  and _47171_ (_39769_, _39744_, _39768_);
  nand _47172_ (_39770_, _39769_, _32431_);
  not _47173_ (_39771_, _39763_);
  or _47174_ (_39772_, _39769_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _47175_ (_39773_, _39772_, _39771_);
  and _47176_ (_39774_, _39773_, _39770_);
  nor _47177_ (_39775_, _39771_, _39298_);
  or _47178_ (_39776_, _39775_, _39774_);
  and _47179_ (_17358_, _39776_, _43634_);
  or _47180_ (_39777_, _24624_, _24592_);
  or _47181_ (_39778_, _39777_, _24656_);
  or _47182_ (_39779_, _39778_, _24698_);
  or _47183_ (_39780_, _39779_, _24772_);
  or _47184_ (_39781_, _39780_, _24804_);
  and _47185_ (_39782_, _39781_, _19525_);
  or _47186_ (_39783_, _32006_, _30365_);
  not _47187_ (_39784_, _31995_);
  nand _47188_ (_39785_, _39784_, _30365_);
  and _47189_ (_39786_, _39785_, _29171_);
  and _47190_ (_39787_, _39786_, _39783_);
  not _47191_ (_39788_, _29192_);
  nand _47192_ (_39790_, _30813_, _39788_);
  or _47193_ (_39794_, _30813_, _29203_);
  and _47194_ (_39800_, _30452_, _39794_);
  and _47195_ (_39805_, _39800_, _39790_);
  and _47196_ (_39812_, _24868_, _21074_);
  and _47197_ (_39820_, _39812_, _20085_);
  and _47198_ (_39828_, _39820_, _26059_);
  nand _47199_ (_39829_, _39828_, _39434_);
  nand _47200_ (_39830_, _39829_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _47201_ (_39831_, _39830_, _39805_);
  or _47202_ (_39832_, _39831_, _39787_);
  or _47203_ (_39833_, _39832_, _35357_);
  or _47204_ (_39834_, _39833_, _29138_);
  or _47205_ (_39835_, _39834_, _39782_);
  nor _47206_ (_39836_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _47207_ (_39837_, _39836_, _39744_);
  and _47208_ (_39838_, _39837_, _39835_);
  and _47209_ (_39839_, _34520_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _47210_ (_39840_, _39839_, _34531_);
  and _47211_ (_39841_, _39840_, _39744_);
  or _47212_ (_39842_, _39841_, _39763_);
  or _47213_ (_39843_, _39842_, _39838_);
  nand _47214_ (_39844_, _39763_, _39291_);
  and _47215_ (_39845_, _39844_, _43634_);
  and _47216_ (_17369_, _39845_, _39843_);
  and _47217_ (_39846_, _39744_, _35217_);
  nand _47218_ (_39847_, _39846_, _32431_);
  or _47219_ (_39848_, _39846_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _47220_ (_39849_, _39848_, _39771_);
  and _47221_ (_39850_, _39849_, _39847_);
  nor _47222_ (_39851_, _39771_, _39284_);
  or _47223_ (_39852_, _39851_, _39850_);
  and _47224_ (_17380_, _39852_, _43634_);
  not _47225_ (_39853_, _39744_);
  or _47226_ (_39854_, _39853_, _36000_);
  and _47227_ (_39855_, _39854_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _47228_ (_39856_, _35989_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _47229_ (_39857_, _39856_, _36033_);
  and _47230_ (_39858_, _39857_, _39744_);
  or _47231_ (_39859_, _39858_, _39855_);
  and _47232_ (_39860_, _39859_, _39771_);
  nor _47233_ (_39861_, _39771_, _39276_);
  or _47234_ (_39862_, _39861_, _39860_);
  and _47235_ (_17391_, _39862_, _43634_);
  and _47236_ (_39868_, _39744_, _36762_);
  nand _47237_ (_39879_, _39868_, _32431_);
  or _47238_ (_39880_, _39868_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _47239_ (_39881_, _39880_, _39771_);
  and _47240_ (_39882_, _39881_, _39879_);
  nor _47241_ (_39893_, _39771_, _39268_);
  or _47242_ (_39899_, _39893_, _39882_);
  and _47243_ (_17402_, _39899_, _43634_);
  and _47244_ (_39900_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _47245_ (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _47246_ (_39902_, _30321_, _29171_);
  and _47247_ (_39903_, _30452_, _30714_);
  nand _47248_ (_39904_, _31602_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _47249_ (_39905_, _39904_, _39900_);
  or _47250_ (_39906_, _39905_, _39903_);
  or _47251_ (_39907_, _39906_, _39902_);
  and _47252_ (_39908_, _39907_, _39901_);
  or _47253_ (_39909_, _39908_, _39744_);
  not _47254_ (_39910_, _37502_);
  nor _47255_ (_39911_, _39910_, _32431_);
  or _47256_ (_39912_, _37502_, _34781_);
  nand _47257_ (_39913_, _39912_, _39744_);
  or _47258_ (_39914_, _39913_, _39911_);
  and _47259_ (_39915_, _39914_, _39909_);
  or _47260_ (_39916_, _39915_, _39763_);
  nand _47261_ (_39917_, _39763_, _39261_);
  and _47262_ (_39918_, _39917_, _43634_);
  and _47263_ (_17413_, _39918_, _39916_);
  not _47264_ (_39919_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _47265_ (_39920_, _39374_, _39919_);
  not _47266_ (_39921_, _39920_);
  nor _47267_ (_39922_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _47268_ (_39923_, _39922_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _47269_ (_39924_, _28271_, _28918_);
  and _47270_ (_39925_, _29061_, _39741_);
  and _47271_ (_39926_, _39925_, _39760_);
  and _47272_ (_39927_, _39926_, _39924_);
  and _47273_ (_39928_, _39927_, _31886_);
  nor _47274_ (_39929_, _39928_, _39923_);
  nor _47275_ (_39930_, _39929_, _31809_);
  and _47276_ (_39931_, _29061_, _28918_);
  and _47277_ (_39932_, _39931_, _28622_);
  not _47278_ (_39933_, _32507_);
  nor _47279_ (_39934_, _39933_, _28765_);
  and _47280_ (_39935_, _39934_, _39932_);
  and _47281_ (_39936_, _39935_, _32463_);
  and _47282_ (_39937_, _39936_, _32431_);
  nor _47283_ (_39938_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _47284_ (_39939_, _39929_, _39921_);
  not _47285_ (_39940_, _39939_);
  nor _47286_ (_39941_, _39940_, _39938_);
  not _47287_ (_39942_, _39941_);
  nor _47288_ (_39943_, _39942_, _39937_);
  or _47289_ (_39944_, _39943_, _39930_);
  and _47290_ (_39945_, _39944_, _39921_);
  nor _47291_ (_39946_, _39921_, _39463_);
  or _47292_ (_39947_, _39946_, _39945_);
  and _47293_ (_17982_, _39947_, _43634_);
  nor _47294_ (_39948_, _39921_, _39507_);
  not _47295_ (_39949_, _39929_);
  and _47296_ (_39950_, _39949_, _32953_);
  not _47297_ (_39951_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _47298_ (_39952_, _39935_, _39951_);
  nor _47299_ (_39953_, _39952_, _39949_);
  and _47300_ (_39954_, _39931_, _28776_);
  and _47301_ (_39955_, _32507_, _28622_);
  and _47302_ (_39956_, _39955_, _39954_);
  not _47303_ (_39957_, _28271_);
  nor _47304_ (_39958_, _32431_, _39957_);
  nor _47305_ (_39959_, _28271_, _39951_);
  nor _47306_ (_39960_, _39959_, _39958_);
  not _47307_ (_39961_, _39960_);
  nand _47308_ (_39962_, _39961_, _39956_);
  and _47309_ (_39963_, _39962_, _39953_);
  nor _47310_ (_39964_, _39963_, _39920_);
  not _47311_ (_39965_, _39964_);
  nor _47312_ (_39966_, _39965_, _39950_);
  nor _47313_ (_39967_, _39966_, _39948_);
  nor _47314_ (_19709_, _39967_, rst);
  nor _47315_ (_39968_, _39921_, _39539_);
  and _47316_ (_39969_, _39949_, _33639_);
  not _47317_ (_39970_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _47318_ (_39971_, _39935_, _39970_);
  nor _47319_ (_39972_, _39971_, _39949_);
  not _47320_ (_39973_, _39972_);
  not _47321_ (_39974_, _39768_);
  nor _47322_ (_39975_, _39974_, _32431_);
  nor _47323_ (_39976_, _39768_, _39970_);
  nor _47324_ (_39977_, _39976_, _39975_);
  and _47325_ (_39978_, _39939_, _39956_);
  not _47326_ (_39979_, _39978_);
  nor _47327_ (_39980_, _39979_, _39977_);
  nor _47328_ (_39981_, _39980_, _39973_);
  nor _47329_ (_39982_, _39981_, _39920_);
  not _47330_ (_39983_, _39982_);
  nor _47331_ (_39984_, _39983_, _39969_);
  nor _47332_ (_39985_, _39984_, _39968_);
  nor _47333_ (_19721_, _39985_, rst);
  nor _47334_ (_39986_, _39929_, _34378_);
  not _47335_ (_39987_, _39935_);
  and _47336_ (_39988_, _39939_, _39987_);
  and _47337_ (_39989_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _47338_ (_39990_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _47339_ (_39991_, _34509_, _39990_);
  nor _47340_ (_39992_, _39991_, _34531_);
  nor _47341_ (_39993_, _39992_, _39979_);
  nor _47342_ (_39994_, _39993_, _39989_);
  not _47343_ (_39995_, _39994_);
  nor _47344_ (_39996_, _39995_, _39986_);
  nor _47345_ (_39997_, _39996_, _39920_);
  nor _47346_ (_39998_, _39921_, _39569_);
  nor _47347_ (_39999_, _39998_, _39997_);
  nor _47348_ (_19733_, _39999_, rst);
  nor _47349_ (_40000_, _39929_, _35118_);
  and _47350_ (_40001_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not _47351_ (_40002_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _47352_ (_40003_, _35217_, _40002_);
  nor _47353_ (_40004_, _40003_, _35227_);
  nor _47354_ (_40005_, _40004_, _39979_);
  nor _47355_ (_40006_, _40005_, _40001_);
  not _47356_ (_40007_, _40006_);
  nor _47357_ (_40008_, _40007_, _40000_);
  nor _47358_ (_40009_, _40008_, _39920_);
  nor _47359_ (_40010_, _39921_, _39600_);
  nor _47360_ (_40011_, _40010_, _40009_);
  nor _47361_ (_19744_, _40011_, rst);
  nor _47362_ (_40012_, _39929_, _35880_);
  and _47363_ (_40013_, _39935_, _35978_);
  nor _47364_ (_40014_, _40013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _47365_ (_40015_, _40014_);
  and _47366_ (_40016_, _40013_, _32431_);
  nor _47367_ (_40017_, _40016_, _39940_);
  and _47368_ (_40018_, _40017_, _40015_);
  or _47369_ (_40019_, _40018_, _40012_);
  and _47370_ (_40020_, _40019_, _39921_);
  nor _47371_ (_40021_, _39921_, _39631_);
  or _47372_ (_40022_, _40021_, _40020_);
  and _47373_ (_19756_, _40022_, _43634_);
  nor _47374_ (_40023_, _39929_, _36675_);
  and _47375_ (_40024_, _39935_, _36762_);
  and _47376_ (_40025_, _40024_, _32431_);
  nor _47377_ (_40026_, _40024_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _47378_ (_40027_, _40026_, _39940_);
  not _47379_ (_40028_, _40027_);
  nor _47380_ (_40029_, _40028_, _40025_);
  or _47381_ (_40030_, _40029_, _40023_);
  and _47382_ (_40031_, _40030_, _39921_);
  nor _47383_ (_40032_, _39921_, _39664_);
  or _47384_ (_40033_, _40032_, _40031_);
  and _47385_ (_19768_, _40033_, _43634_);
  nor _47386_ (_40034_, _39929_, _37403_);
  and _47387_ (_40035_, _39935_, _37502_);
  and _47388_ (_40036_, _40035_, _32431_);
  nor _47389_ (_40037_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _47390_ (_40038_, _40037_, _39940_);
  not _47391_ (_40039_, _40038_);
  nor _47392_ (_40040_, _40039_, _40036_);
  or _47393_ (_40041_, _40040_, _40034_);
  and _47394_ (_40042_, _40041_, _39921_);
  nor _47395_ (_40043_, _39921_, _39693_);
  or _47396_ (_40044_, _40043_, _40042_);
  and _47397_ (_19780_, _40044_, _43634_);
  and _47398_ (_40045_, _28611_, _28490_);
  and _47399_ (_40046_, _39954_, _40045_);
  and _47400_ (_40047_, _40046_, _32463_);
  nand _47401_ (_40048_, _40047_, _32431_);
  or _47402_ (_40049_, _40047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _47403_ (_40050_, _40049_, _32507_);
  and _47404_ (_40051_, _40050_, _40048_);
  and _47405_ (_40052_, _39242_, _39924_);
  nand _47406_ (_40053_, _40052_, _39327_);
  or _47407_ (_40054_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _47408_ (_40055_, _40054_, _31886_);
  and _47409_ (_40056_, _40055_, _40053_);
  not _47410_ (_40057_, _31875_);
  and _47411_ (_40058_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _47412_ (_40059_, _40058_, rst);
  or _47413_ (_40060_, _40059_, _40056_);
  or _47414_ (_30987_, _40060_, _40051_);
  and _47415_ (_40061_, _40045_, _29083_);
  and _47416_ (_40062_, _40061_, _32463_);
  nand _47417_ (_40063_, _40062_, _32431_);
  or _47418_ (_40064_, _40062_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _47419_ (_40065_, _40064_, _32507_);
  and _47420_ (_40066_, _40065_, _40063_);
  and _47421_ (_40067_, _39759_, _39241_);
  and _47422_ (_40068_, _40067_, _39924_);
  nand _47423_ (_40069_, _40068_, _39327_);
  or _47424_ (_40070_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _47425_ (_40071_, _40070_, _31886_);
  and _47426_ (_40072_, _40071_, _40069_);
  and _47427_ (_40073_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _47428_ (_40074_, _40073_, rst);
  or _47429_ (_40075_, _40074_, _40072_);
  or _47430_ (_31010_, _40075_, _40066_);
  and _47431_ (_40094_, _39741_, _28490_);
  and _47432_ (_40105_, _40094_, _39954_);
  and _47433_ (_40114_, _40105_, _32463_);
  nand _47434_ (_40120_, _40114_, _32431_);
  or _47435_ (_40131_, _40114_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _47436_ (_40142_, _40131_, _32507_);
  and _47437_ (_40153_, _40142_, _40120_);
  and _47438_ (_40164_, _39925_, _39241_);
  and _47439_ (_40175_, _40164_, _39924_);
  not _47440_ (_40186_, _40175_);
  nor _47441_ (_40197_, _40186_, _39327_);
  and _47442_ (_40208_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _47443_ (_40219_, _40208_, _40197_);
  and _47444_ (_40230_, _40219_, _31886_);
  and _47445_ (_40241_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _47446_ (_40252_, _40241_, rst);
  or _47447_ (_40263_, _40252_, _40230_);
  or _47448_ (_31033_, _40263_, _40153_);
  and _47449_ (_40284_, _40094_, _29083_);
  and _47450_ (_40288_, _40284_, _32463_);
  nand _47451_ (_40289_, _40288_, _32431_);
  or _47452_ (_40290_, _40288_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _47453_ (_40291_, _40290_, _32507_);
  and _47454_ (_40292_, _40291_, _40289_);
  nor _47455_ (_40293_, _29061_, _28611_);
  and _47456_ (_40294_, _39241_, _40293_);
  and _47457_ (_40295_, _40294_, _39924_);
  not _47458_ (_40296_, _40295_);
  nor _47459_ (_40297_, _40296_, _39327_);
  and _47460_ (_40298_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _47461_ (_40299_, _40298_, _40297_);
  and _47462_ (_40300_, _40299_, _31886_);
  and _47463_ (_40301_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _47464_ (_40302_, _40301_, rst);
  or _47465_ (_40303_, _40302_, _40300_);
  or _47466_ (_31056_, _40303_, _40292_);
  or _47467_ (_40304_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _47468_ (_40305_, _40304_, _32507_);
  and _47469_ (_40306_, _40046_, _28271_);
  nand _47470_ (_40307_, _40306_, _32431_);
  and _47471_ (_40308_, _40307_, _40305_);
  nand _47472_ (_40309_, _40052_, _39306_);
  and _47473_ (_40310_, _40309_, _31886_);
  and _47474_ (_40311_, _40310_, _40304_);
  and _47475_ (_40312_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _47476_ (_40313_, _40312_, rst);
  or _47477_ (_40314_, _40313_, _40311_);
  or _47478_ (_41329_, _40314_, _40308_);
  and _47479_ (_40315_, _39768_, _28918_);
  and _47480_ (_40316_, _40315_, _39242_);
  nand _47481_ (_40317_, _40316_, _32431_);
  or _47482_ (_40318_, _40316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _47483_ (_40319_, _40318_, _32507_);
  and _47484_ (_40320_, _40319_, _40317_);
  nand _47485_ (_40321_, _40052_, _39298_);
  or _47486_ (_40322_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _47487_ (_40323_, _40322_, _31886_);
  and _47488_ (_40324_, _40323_, _40321_);
  and _47489_ (_40325_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _47490_ (_40326_, _40325_, rst);
  or _47491_ (_40327_, _40326_, _40324_);
  or _47492_ (_41331_, _40327_, _40320_);
  not _47493_ (_40328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  not _47494_ (_40329_, _35238_);
  and _47495_ (_40330_, _40046_, _40329_);
  nor _47496_ (_40331_, _40330_, _40328_);
  and _47497_ (_40332_, _34542_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _47498_ (_40333_, _40332_, _34531_);
  and _47499_ (_40334_, _40333_, _40046_);
  or _47500_ (_40335_, _40334_, _40331_);
  and _47501_ (_40336_, _40335_, _32507_);
  nand _47502_ (_40337_, _40052_, _39291_);
  or _47503_ (_40338_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _47504_ (_40339_, _40338_, _31886_);
  and _47505_ (_40340_, _40339_, _40337_);
  nor _47506_ (_40341_, _31875_, _40328_);
  or _47507_ (_40342_, _40341_, rst);
  or _47508_ (_40343_, _40342_, _40340_);
  or _47509_ (_41333_, _40343_, _40336_);
  and _47510_ (_40344_, _40046_, _35217_);
  nand _47511_ (_40345_, _40344_, _32431_);
  or _47512_ (_40346_, _40344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47513_ (_40347_, _40346_, _32507_);
  and _47514_ (_40348_, _40347_, _40345_);
  nand _47515_ (_40349_, _40052_, _39284_);
  or _47516_ (_40350_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _47517_ (_40351_, _40350_, _31886_);
  and _47518_ (_40352_, _40351_, _40349_);
  and _47519_ (_40353_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _47520_ (_40354_, _40353_, rst);
  or _47521_ (_40355_, _40354_, _40352_);
  or _47522_ (_41335_, _40355_, _40348_);
  not _47523_ (_40356_, _40046_);
  or _47524_ (_40357_, _40356_, _36000_);
  and _47525_ (_40358_, _40357_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _47526_ (_40359_, _35989_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _47527_ (_40360_, _40359_, _36033_);
  and _47528_ (_40361_, _40360_, _40046_);
  or _47529_ (_40362_, _40361_, _40358_);
  and _47530_ (_40363_, _40362_, _32507_);
  nand _47531_ (_40364_, _40052_, _39276_);
  or _47532_ (_40365_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _47533_ (_40366_, _40365_, _31886_);
  and _47534_ (_40367_, _40366_, _40364_);
  and _47535_ (_40368_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _47536_ (_40369_, _40368_, rst);
  or _47537_ (_40370_, _40369_, _40367_);
  or _47538_ (_41337_, _40370_, _40363_);
  and _47539_ (_40371_, _40046_, _36762_);
  nand _47540_ (_40372_, _40371_, _32431_);
  or _47541_ (_40373_, _40371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _47542_ (_40374_, _40373_, _32507_);
  and _47543_ (_40375_, _40374_, _40372_);
  nand _47544_ (_40376_, _40052_, _39268_);
  or _47545_ (_40377_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _47546_ (_40378_, _40377_, _31886_);
  and _47547_ (_40379_, _40378_, _40376_);
  and _47548_ (_40380_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _47549_ (_40381_, _40380_, rst);
  or _47550_ (_40382_, _40381_, _40379_);
  or _47551_ (_41339_, _40382_, _40375_);
  and _47552_ (_40383_, _40046_, _37502_);
  nand _47553_ (_40384_, _40383_, _32431_);
  or _47554_ (_40385_, _40383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47555_ (_40386_, _40385_, _32507_);
  and _47556_ (_40387_, _40386_, _40384_);
  nand _47557_ (_40388_, _40052_, _39261_);
  or _47558_ (_40389_, _40052_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _47559_ (_40390_, _40389_, _31886_);
  and _47560_ (_40391_, _40390_, _40388_);
  and _47561_ (_40392_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _47562_ (_40393_, _40392_, rst);
  or _47563_ (_40394_, _40393_, _40391_);
  or _47564_ (_41341_, _40394_, _40387_);
  and _47565_ (_40395_, _40061_, _28271_);
  nand _47566_ (_40396_, _40395_, _32431_);
  or _47567_ (_40397_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _47568_ (_40398_, _40397_, _32507_);
  and _47569_ (_40399_, _40398_, _40396_);
  nand _47570_ (_40400_, _40068_, _39306_);
  and _47571_ (_40401_, _40400_, _31886_);
  and _47572_ (_40402_, _40401_, _40397_);
  and _47573_ (_40403_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _47574_ (_40404_, _40403_, rst);
  or _47575_ (_40405_, _40404_, _40402_);
  or _47576_ (_41343_, _40405_, _40399_);
  and _47577_ (_40406_, _40061_, _39768_);
  nand _47578_ (_40407_, _40406_, _32431_);
  or _47579_ (_40408_, _40406_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _47580_ (_40409_, _40408_, _32507_);
  and _47581_ (_40410_, _40409_, _40407_);
  nand _47582_ (_40411_, _40068_, _39298_);
  or _47583_ (_40412_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _47584_ (_40413_, _40412_, _31886_);
  and _47585_ (_40414_, _40413_, _40411_);
  and _47586_ (_40415_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _47587_ (_40416_, _40415_, rst);
  or _47588_ (_40417_, _40416_, _40414_);
  or _47589_ (_41345_, _40417_, _40410_);
  and _47590_ (_40418_, _40061_, _34509_);
  nand _47591_ (_40419_, _40418_, _32431_);
  or _47592_ (_40420_, _40418_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47593_ (_40421_, _40420_, _32507_);
  and _47594_ (_40422_, _40421_, _40419_);
  nand _47595_ (_40423_, _40068_, _39291_);
  or _47596_ (_40424_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _47597_ (_40425_, _40424_, _31886_);
  and _47598_ (_40426_, _40425_, _40423_);
  and _47599_ (_40427_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _47600_ (_40428_, _40427_, rst);
  or _47601_ (_40429_, _40428_, _40426_);
  or _47602_ (_41347_, _40429_, _40422_);
  and _47603_ (_40430_, _40061_, _35217_);
  nand _47604_ (_40431_, _40430_, _32431_);
  or _47605_ (_40432_, _40430_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47606_ (_40433_, _40432_, _32507_);
  and _47607_ (_40434_, _40433_, _40431_);
  nand _47608_ (_40435_, _40068_, _39284_);
  or _47609_ (_40436_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47610_ (_40437_, _40436_, _31886_);
  and _47611_ (_40438_, _40437_, _40435_);
  and _47612_ (_40439_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _47613_ (_40440_, _40439_, rst);
  or _47614_ (_40441_, _40440_, _40438_);
  or _47615_ (_41348_, _40441_, _40434_);
  and _47616_ (_40442_, _40061_, _35978_);
  nand _47617_ (_40443_, _40442_, _32431_);
  or _47618_ (_40444_, _40442_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47619_ (_40445_, _40444_, _32507_);
  and _47620_ (_40446_, _40445_, _40443_);
  nand _47621_ (_40447_, _40068_, _39276_);
  or _47622_ (_40448_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47623_ (_40449_, _40448_, _31886_);
  and _47624_ (_40450_, _40449_, _40447_);
  and _47625_ (_40451_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _47626_ (_40452_, _40451_, rst);
  or _47627_ (_40453_, _40452_, _40450_);
  or _47628_ (_41350_, _40453_, _40446_);
  and _47629_ (_40454_, _40061_, _36762_);
  nand _47630_ (_40455_, _40454_, _32431_);
  or _47631_ (_40456_, _40454_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47632_ (_40457_, _40456_, _32507_);
  and _47633_ (_40458_, _40457_, _40455_);
  nand _47634_ (_40459_, _40068_, _39268_);
  or _47635_ (_40460_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47636_ (_40461_, _40460_, _31886_);
  and _47637_ (_40462_, _40461_, _40459_);
  and _47638_ (_40463_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _47639_ (_40464_, _40463_, rst);
  or _47640_ (_40465_, _40464_, _40462_);
  or _47641_ (_41352_, _40465_, _40458_);
  and _47642_ (_40466_, _40061_, _37502_);
  nand _47643_ (_40467_, _40466_, _32431_);
  or _47644_ (_40468_, _40466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47645_ (_40469_, _40468_, _32507_);
  and _47646_ (_40470_, _40469_, _40467_);
  nand _47647_ (_40471_, _40068_, _39261_);
  or _47648_ (_40472_, _40068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47649_ (_40473_, _40472_, _31886_);
  and _47650_ (_40474_, _40473_, _40471_);
  and _47651_ (_40475_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _47652_ (_40476_, _40475_, rst);
  or _47653_ (_40477_, _40476_, _40474_);
  or _47654_ (_41354_, _40477_, _40470_);
  and _47655_ (_40478_, _40105_, _28271_);
  nand _47656_ (_40479_, _40478_, _32431_);
  or _47657_ (_40480_, _40478_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _47658_ (_40481_, _40480_, _32507_);
  and _47659_ (_40482_, _40481_, _40479_);
  and _47660_ (_40483_, _40175_, _39307_);
  and _47661_ (_40484_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _47662_ (_40485_, _40484_, _40483_);
  and _47663_ (_40486_, _40485_, _31886_);
  and _47664_ (_40487_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _47665_ (_40488_, _40487_, rst);
  or _47666_ (_40489_, _40488_, _40486_);
  or _47667_ (_41356_, _40489_, _40482_);
  and _47668_ (_40490_, _40105_, _39768_);
  nand _47669_ (_40491_, _40490_, _32431_);
  or _47670_ (_40492_, _40490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _47671_ (_40493_, _40492_, _32507_);
  and _47672_ (_40494_, _40493_, _40491_);
  nor _47673_ (_40495_, _40186_, _39298_);
  and _47674_ (_40496_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47675_ (_40497_, _40496_, _40495_);
  and _47676_ (_40498_, _40497_, _31886_);
  and _47677_ (_40503_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47678_ (_40505_, _40503_, rst);
  or _47679_ (_40506_, _40505_, _40498_);
  or _47680_ (_41358_, _40506_, _40494_);
  and _47681_ (_40507_, _40105_, _34509_);
  nand _47682_ (_40508_, _40507_, _32431_);
  or _47683_ (_40509_, _40507_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _47684_ (_40510_, _40509_, _32507_);
  and _47685_ (_40511_, _40510_, _40508_);
  nor _47686_ (_40512_, _40186_, _39291_);
  and _47687_ (_40513_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47688_ (_40514_, _40513_, _40512_);
  and _47689_ (_40515_, _40514_, _31886_);
  and _47690_ (_40516_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47691_ (_40517_, _40516_, rst);
  or _47692_ (_40518_, _40517_, _40515_);
  or _47693_ (_41360_, _40518_, _40511_);
  and _47694_ (_40519_, _40105_, _35217_);
  nand _47695_ (_40520_, _40519_, _32431_);
  or _47696_ (_40521_, _40519_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _47697_ (_40522_, _40521_, _32507_);
  and _47698_ (_40523_, _40522_, _40520_);
  nor _47699_ (_40524_, _40186_, _39284_);
  and _47700_ (_40525_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47701_ (_40526_, _40525_, _40524_);
  and _47702_ (_40527_, _40526_, _31886_);
  and _47703_ (_40528_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47704_ (_40529_, _40528_, rst);
  or _47705_ (_40530_, _40529_, _40527_);
  or _47706_ (_41362_, _40530_, _40523_);
  and _47707_ (_40538_, _40105_, _35978_);
  nand _47708_ (_40549_, _40538_, _32431_);
  or _47709_ (_40560_, _40538_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _47710_ (_40562_, _40560_, _32507_);
  and _47711_ (_40563_, _40562_, _40549_);
  nor _47712_ (_40564_, _40186_, _39276_);
  and _47713_ (_40565_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47714_ (_40566_, _40565_, _40564_);
  and _47715_ (_40567_, _40566_, _31886_);
  and _47716_ (_40568_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47717_ (_40569_, _40568_, rst);
  or _47718_ (_40570_, _40569_, _40567_);
  or _47719_ (_41363_, _40570_, _40563_);
  and _47720_ (_40571_, _40105_, _36762_);
  nand _47721_ (_40572_, _40571_, _32431_);
  or _47722_ (_40573_, _40571_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _47723_ (_40574_, _40573_, _32507_);
  and _47724_ (_40575_, _40574_, _40572_);
  nor _47725_ (_40576_, _40186_, _39268_);
  and _47726_ (_40577_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47727_ (_40578_, _40577_, _40576_);
  and _47728_ (_40579_, _40578_, _31886_);
  and _47729_ (_40580_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47730_ (_40581_, _40580_, rst);
  or _47731_ (_40582_, _40581_, _40579_);
  or _47732_ (_41365_, _40582_, _40575_);
  and _47733_ (_40583_, _40105_, _37502_);
  nand _47734_ (_40584_, _40583_, _32431_);
  or _47735_ (_40585_, _40583_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47736_ (_40586_, _40585_, _32507_);
  and _47737_ (_40587_, _40586_, _40584_);
  nor _47738_ (_40588_, _40186_, _39261_);
  and _47739_ (_40589_, _40186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47740_ (_40591_, _40589_, _40588_);
  and _47741_ (_40597_, _40591_, _31886_);
  and _47742_ (_40598_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47743_ (_40599_, _40598_, rst);
  or _47744_ (_40600_, _40599_, _40597_);
  or _47745_ (_41367_, _40600_, _40587_);
  and _47746_ (_40601_, _40284_, _28271_);
  nand _47747_ (_40602_, _40601_, _32431_);
  or _47748_ (_40603_, _40601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _47749_ (_40604_, _40603_, _32507_);
  and _47750_ (_40605_, _40604_, _40602_);
  and _47751_ (_40606_, _40295_, _39307_);
  and _47752_ (_40607_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _47753_ (_40608_, _40607_, _40606_);
  and _47754_ (_40609_, _40608_, _31886_);
  and _47755_ (_40610_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _47756_ (_40611_, _40610_, rst);
  or _47757_ (_40612_, _40611_, _40609_);
  or _47758_ (_41369_, _40612_, _40605_);
  and _47759_ (_40613_, _40284_, _39768_);
  nand _47760_ (_40614_, _40613_, _32431_);
  or _47761_ (_40615_, _40613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _47762_ (_40616_, _40615_, _32507_);
  and _47763_ (_40617_, _40616_, _40614_);
  nor _47764_ (_40618_, _40296_, _39298_);
  and _47765_ (_40619_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47766_ (_40620_, _40619_, _40618_);
  and _47767_ (_40621_, _40620_, _31886_);
  and _47768_ (_40622_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47769_ (_40623_, _40622_, rst);
  or _47770_ (_40624_, _40623_, _40621_);
  or _47771_ (_41370_, _40624_, _40617_);
  and _47772_ (_40625_, _40284_, _34509_);
  nand _47773_ (_40626_, _40625_, _32431_);
  or _47774_ (_40627_, _40625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47775_ (_40628_, _40627_, _32507_);
  and _47776_ (_40629_, _40628_, _40626_);
  nor _47777_ (_40630_, _40296_, _39291_);
  and _47778_ (_40631_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47779_ (_40632_, _40631_, _40630_);
  and _47780_ (_40633_, _40632_, _31886_);
  and _47781_ (_40634_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47782_ (_40635_, _40634_, rst);
  or _47783_ (_40636_, _40635_, _40633_);
  or _47784_ (_41372_, _40636_, _40629_);
  and _47785_ (_40637_, _40284_, _35217_);
  nand _47786_ (_40638_, _40637_, _32431_);
  or _47787_ (_40639_, _40637_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47788_ (_40640_, _40639_, _32507_);
  and _47789_ (_40641_, _40640_, _40638_);
  nor _47790_ (_40642_, _40296_, _39284_);
  and _47791_ (_40643_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47792_ (_40644_, _40643_, _40642_);
  and _47793_ (_40645_, _40644_, _31886_);
  and _47794_ (_40646_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47795_ (_40647_, _40646_, rst);
  or _47796_ (_40648_, _40647_, _40645_);
  or _47797_ (_41374_, _40648_, _40641_);
  and _47798_ (_40649_, _40284_, _35978_);
  nand _47799_ (_40650_, _40649_, _32431_);
  or _47800_ (_40651_, _40649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47801_ (_40652_, _40651_, _32507_);
  and _47802_ (_40653_, _40652_, _40650_);
  nor _47803_ (_40654_, _40296_, _39276_);
  and _47804_ (_40655_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47805_ (_40656_, _40655_, _40654_);
  and _47806_ (_40657_, _40656_, _31886_);
  and _47807_ (_40658_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47808_ (_40659_, _40658_, rst);
  or _47809_ (_40660_, _40659_, _40657_);
  or _47810_ (_41376_, _40660_, _40653_);
  and _47811_ (_40661_, _40284_, _36762_);
  nand _47812_ (_40662_, _40661_, _32431_);
  or _47813_ (_40663_, _40661_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47814_ (_40664_, _40663_, _32507_);
  and _47815_ (_40665_, _40664_, _40662_);
  nor _47816_ (_40666_, _40296_, _39268_);
  and _47817_ (_40667_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47818_ (_40668_, _40667_, _40666_);
  and _47819_ (_40669_, _40668_, _31886_);
  and _47820_ (_40670_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47821_ (_40671_, _40670_, rst);
  or _47822_ (_40676_, _40671_, _40669_);
  or _47823_ (_41377_, _40676_, _40665_);
  and _47824_ (_40683_, _40284_, _37502_);
  nand _47825_ (_40684_, _40683_, _32431_);
  or _47826_ (_40685_, _40683_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _47827_ (_40686_, _40685_, _32507_);
  and _47828_ (_40687_, _40686_, _40684_);
  nor _47829_ (_40688_, _40296_, _39261_);
  and _47830_ (_40689_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47831_ (_40690_, _40689_, _40688_);
  and _47832_ (_40691_, _40690_, _31886_);
  and _47833_ (_40692_, _40057_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47834_ (_40693_, _40692_, rst);
  or _47835_ (_40694_, _40693_, _40691_);
  or _47836_ (_41379_, _40694_, _40687_);
  and _47837_ (_41828_, t0_i, _43634_);
  and _47838_ (_41831_, t1_i, _43634_);
  not _47839_ (_40695_, _31886_);
  nor _47840_ (_40696_, _40695_, _28918_);
  and _47841_ (_40697_, _40696_, _35217_);
  and _47842_ (_40698_, _40697_, _39242_);
  nand _47843_ (_40699_, _40698_, _39327_);
  not _47844_ (_40700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47845_ (_40701_, _40700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47846_ (_40702_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47847_ (_40703_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _40702_);
  nor _47848_ (_40704_, _40703_, _40701_);
  nor _47849_ (_40705_, _28008_, _28918_);
  and _47850_ (_40706_, _40705_, _39243_);
  and _47851_ (_40707_, _40706_, _31886_);
  or _47852_ (_40708_, _40707_, _40704_);
  and _47853_ (_40709_, _40708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _47854_ (_40710_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _47855_ (_40711_, t1_i);
  and _47856_ (_40712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _40711_);
  nor _47857_ (_40713_, _40712_, _40710_);
  not _47858_ (_40714_, _40713_);
  not _47859_ (_40715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47860_ (_40716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _40715_);
  nor _47861_ (_40717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _47862_ (_40718_, _40717_);
  and _47863_ (_40719_, _40718_, _40716_);
  and _47864_ (_40720_, _40719_, _40714_);
  and _47865_ (_40721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _47866_ (_40722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47867_ (_40723_, _40722_, _40721_);
  and _47868_ (_40724_, _40723_, _40720_);
  and _47869_ (_40725_, _40724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _47870_ (_40726_, _40725_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47871_ (_40727_, _40726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _47872_ (_40728_, _40727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47873_ (_40729_, _40723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _47874_ (_40730_, _40729_, _40720_);
  and _47875_ (_40731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47876_ (_40732_, _40731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47877_ (_40733_, _40732_, _40730_);
  nor _47878_ (_40734_, _40733_, _40704_);
  and _47879_ (_40735_, _40734_, _40728_);
  and _47880_ (_40736_, _40733_, _40701_);
  and _47881_ (_40737_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47882_ (_40738_, _40737_, _40735_);
  nor _47883_ (_40739_, _40738_, _40707_);
  or _47884_ (_40740_, _40739_, _40709_);
  or _47885_ (_40741_, _40698_, _40740_);
  and _47886_ (_40742_, _40741_, _43634_);
  and _47887_ (_41834_, _40742_, _40699_);
  not _47888_ (_40743_, _40707_);
  nor _47889_ (_40744_, _40743_, _39327_);
  and _47890_ (_40745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47891_ (_40746_, _40745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47892_ (_40747_, _40732_, _40729_);
  and _47893_ (_40748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47894_ (_40749_, _40748_, _40747_);
  and _47895_ (_40751_, _40749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47896_ (_40755_, _40751_, _40720_);
  and _47897_ (_40756_, _40755_, _40746_);
  and _47898_ (_40757_, _40756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47899_ (_40758_, _40757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47900_ (_40759_, _40757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47901_ (_40760_, _40759_, _40758_);
  and _47902_ (_40761_, _40760_, _40703_);
  and _47903_ (_40762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not _47904_ (_40763_, _40746_);
  and _47905_ (_40764_, _40748_, _40729_);
  and _47906_ (_40765_, _40764_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _47907_ (_40766_, _40765_, _40720_);
  nor _47908_ (_40767_, _40766_, _40763_);
  and _47909_ (_40768_, _40767_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47910_ (_40769_, _40768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47911_ (_40770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _47912_ (_40771_, _40768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _47913_ (_40781_, _40771_, _40770_);
  nor _47914_ (_40782_, _40781_, _40769_);
  or _47915_ (_40783_, _40782_, _40762_);
  or _47916_ (_40784_, _40783_, _40761_);
  nand _47917_ (_40785_, _40696_, _39465_);
  and _47918_ (_40786_, _40785_, _40743_);
  and _47919_ (_40787_, _40786_, _40784_);
  not _47920_ (_40788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47921_ (_40789_, _40785_, _40788_);
  or _47922_ (_40790_, _40789_, _40787_);
  or _47923_ (_40791_, _40790_, _40744_);
  and _47924_ (_41837_, _40791_, _43634_);
  not _47925_ (_40792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _47926_ (_40793_, _40720_, _40792_);
  or _47927_ (_40794_, _40793_, _40758_);
  and _47928_ (_40795_, _40794_, _40703_);
  or _47929_ (_40796_, _40793_, _40769_);
  and _47930_ (_40797_, _40796_, _40770_);
  nand _47931_ (_40798_, _40720_, _40700_);
  and _47932_ (_40799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _47933_ (_40800_, _40799_, _40798_);
  or _47934_ (_40801_, _40800_, _40736_);
  or _47935_ (_40802_, _40801_, _40797_);
  or _47936_ (_40803_, _40802_, _40795_);
  and _47937_ (_40804_, _40803_, _43634_);
  and _47938_ (_41840_, _40804_, _40786_);
  and _47939_ (_40805_, _40696_, _35978_);
  and _47940_ (_40806_, _40805_, _39242_);
  nor _47941_ (_40807_, _40806_, rst);
  and _47942_ (_40808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47943_ (_40809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _47944_ (_40810_, _40809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47945_ (_40811_, _40810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47946_ (_40812_, _40811_, _40808_);
  and _47947_ (_40813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47948_ (_40814_, _40813_, _40812_);
  or _47949_ (_40815_, _40814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _47950_ (_40816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _47951_ (_40817_, t0_i);
  and _47952_ (_40818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _40817_);
  nor _47953_ (_40819_, _40818_, _40816_);
  not _47954_ (_40820_, _40819_);
  not _47955_ (_40821_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _47956_ (_40822_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _47957_ (_40823_, _40822_, _40821_);
  and _47958_ (_40824_, _40823_, _40820_);
  and _47959_ (_40825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47960_ (_40826_, _40825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _47961_ (_40827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47962_ (_40828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47963_ (_40829_, _40828_, _40827_);
  and _47964_ (_40830_, _40829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _47965_ (_40831_, _40830_, _40826_);
  and _47966_ (_40832_, _40831_, _40824_);
  nor _47967_ (_40833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _47968_ (_40834_, _40833_);
  and _47969_ (_40835_, _40834_, _40832_);
  and _47970_ (_40836_, _40835_, _40815_);
  not _47971_ (_40837_, _40824_);
  and _47972_ (_40838_, _40837_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _47973_ (_40839_, _40830_, _40824_);
  and _47974_ (_40840_, _40839_, _40812_);
  and _47975_ (_40841_, _40840_, _40813_);
  and _47976_ (_40842_, _40841_, _40833_);
  or _47977_ (_40843_, _40842_, _40838_);
  nor _47978_ (_40844_, _40843_, _40836_);
  and _47979_ (_40845_, _40696_, _34509_);
  and _47980_ (_40846_, _40845_, _39242_);
  nor _47981_ (_40847_, _40846_, _40844_);
  and _47982_ (_41843_, _40847_, _40807_);
  and _47983_ (_40848_, _40833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47984_ (_40849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47985_ (_40850_, _40849_, _40839_);
  or _47986_ (_40851_, _40850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _47987_ (_40852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47988_ (_40853_, _40852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47989_ (_40854_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _47990_ (_40855_, _40833_, _40832_);
  or _47991_ (_40856_, _40855_, _40854_);
  or _47992_ (_40857_, _40856_, _40806_);
  and _47993_ (_40858_, _40857_, _40851_);
  or _47994_ (_40859_, _40858_, _40848_);
  and _47995_ (_40860_, _40696_, _39472_);
  not _47996_ (_40861_, _40860_);
  not _47997_ (_40862_, _40806_);
  or _47998_ (_40863_, _40862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47999_ (_40864_, _40863_, _40861_);
  and _48000_ (_40865_, _40864_, _40859_);
  nor _48001_ (_40866_, _40861_, _39327_);
  or _48002_ (_40867_, _40866_, _40865_);
  and _48003_ (_41846_, _40867_, _43634_);
  nand _48004_ (_40868_, _40806_, _39327_);
  not _48005_ (_40869_, _40846_);
  not _48006_ (_40870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _48007_ (_40871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40870_);
  or _48008_ (_40872_, _40853_, _40871_);
  not _48009_ (_40873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _48010_ (_40874_, _40832_, _40870_);
  and _48011_ (_40875_, _40874_, _40812_);
  and _48012_ (_40876_, _40875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _48013_ (_40877_, _40876_, _40873_);
  and _48014_ (_40878_, _40876_, _40873_);
  or _48015_ (_40879_, _40878_, _40877_);
  and _48016_ (_40880_, _40879_, _40872_);
  and _48017_ (_40881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _48018_ (_40882_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _48019_ (_40883_, _40882_, _40811_);
  and _48020_ (_40884_, _40883_, _40808_);
  and _48021_ (_40885_, _40884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _48022_ (_40886_, _40885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _48023_ (_40887_, _40885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _48024_ (_40888_, _40887_, _40886_);
  and _48025_ (_40889_, _40888_, _40881_);
  and _48026_ (_40890_, _40840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _48027_ (_40891_, _40890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _48028_ (_40892_, _40841_, _40834_);
  and _48029_ (_40893_, _40892_, _40891_);
  or _48030_ (_40894_, _40893_, _40889_);
  or _48031_ (_40895_, _40894_, _40880_);
  or _48032_ (_40896_, _40895_, _40806_);
  and _48033_ (_40897_, _40896_, _40869_);
  and _48034_ (_40898_, _40897_, _40868_);
  and _48035_ (_40899_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _48036_ (_40900_, _40899_, _40898_);
  and _48037_ (_41849_, _40900_, _43634_);
  or _48038_ (_40901_, _40882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and _48039_ (_40902_, _40881_, _43634_);
  nand _48040_ (_40903_, _40902_, _40901_);
  nor _48041_ (_40904_, _40903_, _40806_);
  not _48042_ (_40905_, _40882_);
  nor _48043_ (_40906_, _40905_, _40814_);
  nor _48044_ (_40907_, _40906_, _40846_);
  and _48045_ (_41852_, _40907_, _40904_);
  and _48046_ (_40908_, _40696_, _39249_);
  or _48047_ (_40909_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _48048_ (_40910_, _40909_, _43634_);
  nand _48049_ (_40911_, _40908_, _39327_);
  and _48050_ (_41855_, _40911_, _40910_);
  and _48051_ (_40912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _48052_ (_40913_, _40912_, _40707_);
  and _48053_ (_40914_, _40913_, _40720_);
  not _48054_ (_40915_, _40914_);
  nor _48055_ (_40916_, _40915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _48056_ (_40917_, _40915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _48057_ (_40918_, _40917_, _40916_);
  and _48058_ (_40919_, _40918_, _40785_);
  and _48059_ (_40920_, _40747_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _48060_ (_40921_, _40920_, _40701_);
  and _48061_ (_40922_, _40921_, _40786_);
  and _48062_ (_40923_, _40698_, _39307_);
  or _48063_ (_40924_, _40923_, _40922_);
  or _48064_ (_40925_, _40924_, _40919_);
  and _48065_ (_42352_, _40925_, _43634_);
  nand _48066_ (_40926_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _48067_ (_40927_, _40926_, _40785_);
  nor _48068_ (_40928_, _40927_, _40707_);
  and _48069_ (_40929_, _40720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _48070_ (_40930_, _40913_, _40929_);
  nand _48071_ (_40931_, _40930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _48072_ (_40932_, _40930_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _48073_ (_40933_, _40932_, _40931_);
  or _48074_ (_40934_, _40933_, _40928_);
  nand _48075_ (_40935_, _40698_, _39298_);
  and _48076_ (_40936_, _40935_, _43634_);
  and _48077_ (_42354_, _40936_, _40934_);
  and _48078_ (_40937_, _40929_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _48079_ (_40938_, _40937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _48080_ (_40939_, _40929_, _40721_);
  nor _48081_ (_40940_, _40912_, _40939_);
  and _48082_ (_40941_, _40940_, _40938_);
  and _48083_ (_40942_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _48084_ (_40943_, _40942_, _40941_);
  and _48085_ (_40944_, _40943_, _40786_);
  nand _48086_ (_40945_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _48087_ (_40946_, _40945_, _40913_);
  or _48088_ (_40947_, _40946_, _40944_);
  and _48089_ (_40948_, _35217_, _28929_);
  and _48090_ (_40949_, _40948_, _39242_);
  and _48091_ (_40950_, _40949_, _31886_);
  not _48092_ (_40951_, _40950_);
  nor _48093_ (_40952_, _40951_, _39291_);
  or _48094_ (_40953_, _40952_, _40947_);
  and _48095_ (_42355_, _40953_, _43634_);
  or _48096_ (_40954_, _40939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _48097_ (_40955_, _40912_, _40724_);
  and _48098_ (_40956_, _40955_, _40954_);
  and _48099_ (_40957_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _48100_ (_40958_, _40957_, _40956_);
  and _48101_ (_40959_, _40958_, _40786_);
  nand _48102_ (_40960_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _48103_ (_40961_, _40960_, _40913_);
  or _48104_ (_40962_, _40961_, _40959_);
  nor _48105_ (_40963_, _40951_, _39284_);
  or _48106_ (_40964_, _40963_, _40962_);
  and _48107_ (_42357_, _40964_, _43634_);
  or _48108_ (_40965_, _40724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _48109_ (_40966_, _40912_, _40730_);
  and _48110_ (_40967_, _40966_, _40965_);
  and _48111_ (_40968_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _48112_ (_40969_, _40968_, _40967_);
  and _48113_ (_40970_, _40969_, _40786_);
  nand _48114_ (_40971_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _48115_ (_40972_, _40971_, _40913_);
  or _48116_ (_40973_, _40972_, _40970_);
  nor _48117_ (_40974_, _40951_, _39276_);
  or _48118_ (_40975_, _40974_, _40973_);
  and _48119_ (_42359_, _40975_, _43634_);
  or _48120_ (_40976_, _40730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _48121_ (_40977_, _40730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _48122_ (_40978_, _40977_, _40704_);
  and _48123_ (_40979_, _40978_, _40976_);
  and _48124_ (_40980_, _40736_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _48125_ (_40981_, _40980_, _40979_);
  and _48126_ (_40982_, _40981_, _40786_);
  and _48127_ (_40983_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _48128_ (_40984_, _40983_, _40708_);
  or _48129_ (_40985_, _40984_, _40982_);
  nor _48130_ (_40986_, _40951_, _39268_);
  or _48131_ (_40987_, _40986_, _40985_);
  and _48132_ (_42361_, _40987_, _43634_);
  and _48133_ (_40988_, _40785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _48134_ (_40989_, _40988_, _40708_);
  and _48135_ (_40990_, _40701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _48136_ (_40991_, _40990_, _40720_);
  and _48137_ (_40992_, _40991_, _40747_);
  nor _48138_ (_40993_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _48139_ (_40994_, _40993_, _40704_);
  nor _48140_ (_40995_, _40994_, _40727_);
  or _48141_ (_40996_, _40995_, _40992_);
  and _48142_ (_40997_, _40996_, _40786_);
  or _48143_ (_40998_, _40997_, _40989_);
  nor _48144_ (_40999_, _40951_, _39261_);
  or _48145_ (_41000_, _40999_, _40998_);
  and _48146_ (_42363_, _41000_, _43634_);
  and _48147_ (_41001_, _40730_, _40702_);
  nor _48148_ (_41002_, _40732_, _40700_);
  not _48149_ (_41003_, _41002_);
  and _48150_ (_41004_, _41003_, _41001_);
  and _48151_ (_41005_, _41004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _48152_ (_41006_, _41004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _48153_ (_41007_, _41006_, _41005_);
  and _48154_ (_41008_, _41007_, _40786_);
  and _48155_ (_41009_, _40707_, _39307_);
  not _48156_ (_41010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _48157_ (_41011_, _40785_, _41010_);
  or _48158_ (_41012_, _41011_, _41009_);
  or _48159_ (_41013_, _41012_, _41008_);
  and _48160_ (_42364_, _41013_, _43634_);
  nor _48161_ (_41014_, _40743_, _39298_);
  not _48162_ (_41015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _48163_ (_41016_, _41005_, _41015_);
  and _48164_ (_41017_, _41005_, _41015_);
  or _48165_ (_41018_, _41017_, _41016_);
  and _48166_ (_41019_, _41018_, _40786_);
  nor _48167_ (_41020_, _40785_, _41015_);
  or _48168_ (_41021_, _41020_, _41019_);
  or _48169_ (_41022_, _41021_, _41014_);
  and _48170_ (_42366_, _41022_, _43634_);
  nor _48171_ (_41023_, _40743_, _39291_);
  and _48172_ (_41024_, _40748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _48173_ (_41025_, _41024_, _40730_);
  and _48174_ (_41026_, _41025_, _40702_);
  nand _48175_ (_41027_, _41026_, _41003_);
  and _48176_ (_41028_, _41027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _48177_ (_41029_, _40747_, _40703_);
  and _48178_ (_41030_, _40770_, _40729_);
  or _48179_ (_41031_, _41030_, _41029_);
  not _48180_ (_41032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _48181_ (_41033_, _40748_, _41032_);
  and _48182_ (_41034_, _41033_, _40720_);
  and _48183_ (_41035_, _41034_, _41031_);
  or _48184_ (_41036_, _41035_, _41028_);
  and _48185_ (_41037_, _41036_, _40786_);
  nor _48186_ (_41038_, _40785_, _41032_);
  or _48187_ (_41039_, _41038_, _41037_);
  or _48188_ (_41040_, _41039_, _41023_);
  and _48189_ (_42368_, _41040_, _43634_);
  nor _48190_ (_41041_, _40743_, _39284_);
  and _48191_ (_41042_, _40755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _48192_ (_41043_, _40755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _48193_ (_41044_, _41043_, _40703_);
  nor _48194_ (_41045_, _41044_, _41042_);
  not _48195_ (_41046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _48196_ (_41047_, _41026_, _41046_);
  and _48197_ (_41048_, _41026_, _41046_);
  nor _48198_ (_41049_, _41048_, _41047_);
  nor _48199_ (_41050_, _41049_, _40703_);
  or _48200_ (_41051_, _41050_, _41045_);
  and _48201_ (_41052_, _41051_, _40786_);
  nor _48202_ (_41053_, _40785_, _41046_);
  or _48203_ (_41054_, _41053_, _41052_);
  or _48204_ (_41055_, _41054_, _41041_);
  and _48205_ (_42370_, _41055_, _43634_);
  nor _48206_ (_41056_, _40743_, _39276_);
  not _48207_ (_41057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _48208_ (_41058_, _40785_, _41057_);
  or _48209_ (_41059_, _41042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _48210_ (_41060_, _41059_, _40703_);
  and _48211_ (_41061_, _41042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _48212_ (_41062_, _41061_, _41060_);
  and _48213_ (_41063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _48214_ (_41064_, _40766_, _41046_);
  or _48215_ (_41065_, _41064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _48216_ (_41066_, _41064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _48217_ (_41067_, _41066_, _41065_);
  and _48218_ (_41068_, _41067_, _40770_);
  or _48219_ (_41069_, _41068_, _41063_);
  or _48220_ (_41070_, _41069_, _41062_);
  and _48221_ (_41071_, _41070_, _40786_);
  or _48222_ (_41072_, _41071_, _41058_);
  or _48223_ (_41073_, _41072_, _41056_);
  and _48224_ (_42371_, _41073_, _43634_);
  nand _48225_ (_41074_, _40707_, _39268_);
  and _48226_ (_41075_, _41025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _48227_ (_41076_, _41075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _48228_ (_41077_, _41076_, _40770_);
  and _48229_ (_41078_, _41061_, _40703_);
  nor _48230_ (_41079_, _41078_, _41077_);
  not _48231_ (_41080_, _41079_);
  and _48232_ (_41081_, _41080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _48233_ (_41082_, _41080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _48234_ (_41083_, _41082_, _41081_);
  and _48235_ (_41084_, _41083_, _40785_);
  or _48236_ (_41085_, _41084_, _40707_);
  and _48237_ (_41086_, _41085_, _41074_);
  and _48238_ (_41087_, _40698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _48239_ (_41088_, _41087_, _41086_);
  and _48240_ (_42373_, _41088_, _43634_);
  nand _48241_ (_41089_, _40707_, _39261_);
  not _48242_ (_41090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _48243_ (_41091_, _41076_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _48244_ (_41092_, _41002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand _48245_ (_41093_, _41092_, _41091_);
  nand _48246_ (_41094_, _41093_, _41090_);
  or _48247_ (_41095_, _41093_, _41090_);
  and _48248_ (_41096_, _41095_, _41094_);
  and _48249_ (_41097_, _41096_, _40785_);
  or _48250_ (_41098_, _41097_, _40707_);
  and _48251_ (_41099_, _41098_, _41089_);
  and _48252_ (_41100_, _40698_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _48253_ (_41101_, _41100_, _41099_);
  and _48254_ (_42375_, _41101_, _43634_);
  nor _48255_ (_41102_, _40837_, _40806_);
  or _48256_ (_41103_, _41102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _48257_ (_41104_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _48258_ (_41105_, _41104_, _40831_);
  and _48259_ (_41106_, _40824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _48260_ (_41107_, _41106_, _41105_);
  or _48261_ (_41108_, _41107_, _40806_);
  and _48262_ (_41109_, _41108_, _41103_);
  or _48263_ (_41110_, _41109_, _40846_);
  nand _48264_ (_41111_, _40846_, _39306_);
  and _48265_ (_41112_, _41111_, _43634_);
  and _48266_ (_42377_, _41112_, _41110_);
  nor _48267_ (_41113_, _41106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _48268_ (_41114_, _41106_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _48269_ (_41115_, _41114_, _41113_);
  and _48270_ (_41116_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _48271_ (_41117_, _41116_, _40832_);
  nor _48272_ (_41118_, _41117_, _41115_);
  nor _48273_ (_41119_, _41118_, _40806_);
  and _48274_ (_41120_, _40806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _48275_ (_41121_, _41120_, _41119_);
  and _48276_ (_41122_, _41121_, _40861_);
  nor _48277_ (_41123_, _40869_, _39298_);
  or _48278_ (_41124_, _41123_, _41122_);
  and _48279_ (_42378_, _41124_, _43634_);
  nor _48280_ (_41125_, _41114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _48281_ (_41126_, _41106_, _40827_);
  nor _48282_ (_41127_, _41126_, _41125_);
  and _48283_ (_41128_, _40853_, _40832_);
  and _48284_ (_41129_, _41128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _48285_ (_41130_, _41129_, _41127_);
  nor _48286_ (_41131_, _41130_, _40806_);
  and _48287_ (_41132_, _40806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _48288_ (_41133_, _41132_, _41131_);
  and _48289_ (_41134_, _41133_, _40861_);
  nor _48290_ (_41135_, _40869_, _39291_);
  or _48291_ (_41136_, _41135_, _41134_);
  and _48292_ (_42380_, _41136_, _43634_);
  and _48293_ (_41137_, _40829_, _40824_);
  nor _48294_ (_41138_, _41126_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _48295_ (_41139_, _41138_, _41137_);
  and _48296_ (_41140_, _41128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _48297_ (_41141_, _41140_, _41139_);
  nor _48298_ (_41142_, _41141_, _40806_);
  and _48299_ (_41143_, _40806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _48300_ (_41144_, _41143_, _41142_);
  and _48301_ (_41145_, _41144_, _40861_);
  nor _48302_ (_41146_, _40869_, _39284_);
  or _48303_ (_41147_, _41146_, _41145_);
  and _48304_ (_42382_, _41147_, _43634_);
  nand _48305_ (_41148_, _40846_, _39276_);
  or _48306_ (_41149_, _40862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _48307_ (_41150_, _41137_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _48308_ (_41151_, _41150_, _40839_);
  and _48309_ (_41152_, _41128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _48310_ (_41153_, _41152_, _41151_);
  or _48311_ (_41154_, _41153_, _40806_);
  and _48312_ (_41155_, _41154_, _41149_);
  or _48313_ (_41156_, _41155_, _40846_);
  and _48314_ (_41157_, _41156_, _43634_);
  and _48315_ (_42384_, _41157_, _41148_);
  nand _48316_ (_41158_, _40846_, _39268_);
  and _48317_ (_41159_, _41128_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not _48318_ (_41160_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _48319_ (_41161_, _40834_, _40839_);
  and _48320_ (_41162_, _41161_, _41160_);
  nor _48321_ (_41163_, _41162_, _41159_);
  nor _48322_ (_41164_, _41163_, _40806_);
  and _48323_ (_41165_, _41161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _48324_ (_41166_, _41165_);
  or _48325_ (_41167_, _41166_, _40806_);
  and _48326_ (_41168_, _41167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _48327_ (_41169_, _41168_, _41164_);
  or _48328_ (_41170_, _41169_, _40846_);
  and _48329_ (_41171_, _41170_, _43634_);
  and _48330_ (_42385_, _41171_, _41158_);
  nor _48331_ (_41172_, _41166_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _48332_ (_41173_, _40853_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _48333_ (_41174_, _41173_, _40824_);
  and _48334_ (_41175_, _41174_, _40831_);
  nor _48335_ (_41176_, _41175_, _41172_);
  nor _48336_ (_41177_, _41176_, _40806_);
  and _48337_ (_41178_, _41167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _48338_ (_41179_, _41178_, _41177_);
  and _48339_ (_41180_, _41179_, _40861_);
  nor _48340_ (_41181_, _40869_, _39261_);
  or _48341_ (_41182_, _41181_, _41180_);
  and _48342_ (_42387_, _41182_, _43634_);
  and _48343_ (_41183_, _40874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _48344_ (_41184_, _40874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _48345_ (_41185_, _41184_, _40872_);
  nor _48346_ (_41186_, _41185_, _41183_);
  and _48347_ (_41187_, _40882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _48348_ (_41188_, _40882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _48349_ (_41189_, _41188_, _40881_);
  nor _48350_ (_41190_, _41189_, _41187_);
  and _48351_ (_41191_, _40839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _48352_ (_41192_, _40839_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _48353_ (_41193_, _41192_, _40833_);
  nor _48354_ (_41194_, _41193_, _41191_);
  or _48355_ (_41195_, _41194_, _41190_);
  or _48356_ (_41196_, _41195_, _41186_);
  or _48357_ (_41197_, _41196_, _40806_);
  nand _48358_ (_41198_, _40806_, _39306_);
  and _48359_ (_41199_, _41198_, _40869_);
  and _48360_ (_41200_, _41199_, _41197_);
  and _48361_ (_41201_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _48362_ (_41202_, _41201_, _41200_);
  and _48363_ (_42389_, _41202_, _43634_);
  nand _48364_ (_41203_, _40806_, _39298_);
  or _48365_ (_41204_, _41183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _48366_ (_41205_, _40832_, _40809_);
  not _48367_ (_41206_, _41205_);
  or _48368_ (_41207_, _41206_, _40853_);
  and _48369_ (_41208_, _41207_, _40872_);
  and _48370_ (_41209_, _41208_, _41204_);
  and _48371_ (_41210_, _40882_, _40809_);
  or _48372_ (_41211_, _41187_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _48373_ (_41212_, _41211_, _40881_);
  nor _48374_ (_41213_, _41212_, _41210_);
  and _48375_ (_41214_, _41191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _48376_ (_41215_, _41191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _48377_ (_41216_, _41215_, _40833_);
  nor _48378_ (_41217_, _41216_, _41214_);
  or _48379_ (_41218_, _41217_, _41213_);
  or _48380_ (_41219_, _41218_, _41209_);
  or _48381_ (_41220_, _41219_, _40806_);
  and _48382_ (_41221_, _41220_, _40869_);
  and _48383_ (_41222_, _41221_, _41203_);
  and _48384_ (_41223_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _48385_ (_41224_, _41223_, _41222_);
  and _48386_ (_42391_, _41224_, _43634_);
  nor _48387_ (_41225_, _40862_, _39291_);
  or _48388_ (_41226_, _41205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48389_ (_41227_, _40832_, _40810_);
  not _48390_ (_41228_, _41227_);
  and _48391_ (_41229_, _41228_, _40871_);
  and _48392_ (_41230_, _41229_, _41226_);
  and _48393_ (_41231_, _40824_, _40809_);
  and _48394_ (_41232_, _41231_, _40830_);
  or _48395_ (_41233_, _41232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48396_ (_41234_, _40839_, _40810_);
  nor _48397_ (_41235_, _41234_, _40834_);
  and _48398_ (_41236_, _41235_, _41233_);
  and _48399_ (_41237_, _41210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _48400_ (_41238_, _41237_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48401_ (_41239_, _40882_, _40810_);
  nand _48402_ (_41240_, _41239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _48403_ (_41241_, _41240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _48404_ (_41242_, _41241_, _41238_);
  or _48405_ (_41243_, _41242_, _41236_);
  nor _48406_ (_41244_, _41243_, _41230_);
  nor _48407_ (_41245_, _41244_, _40806_);
  or _48408_ (_41246_, _41245_, _40860_);
  or _48409_ (_41247_, _41246_, _41225_);
  or _48410_ (_41248_, _40861_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48411_ (_41249_, _41248_, _43634_);
  and _48412_ (_42392_, _41249_, _41247_);
  nor _48413_ (_41250_, _40862_, _39284_);
  not _48414_ (_41251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _48415_ (_41252_, _41227_, _40870_);
  nor _48416_ (_41253_, _41252_, _41251_);
  and _48417_ (_41254_, _41252_, _41251_);
  or _48418_ (_41255_, _41254_, _41253_);
  and _48419_ (_41256_, _41255_, _40872_);
  or _48420_ (_41257_, _41239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _48421_ (_41258_, _40883_);
  and _48422_ (_41259_, _41258_, _40881_);
  and _48423_ (_41260_, _41259_, _41257_);
  or _48424_ (_41261_, _41234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _48425_ (_41262_, _40839_, _40811_);
  nor _48426_ (_41263_, _41262_, _40834_);
  and _48427_ (_41264_, _41263_, _41261_);
  or _48428_ (_41265_, _41264_, _41260_);
  nor _48429_ (_41266_, _41265_, _41256_);
  nor _48430_ (_41267_, _41266_, _40806_);
  or _48431_ (_41268_, _41267_, _40860_);
  or _48432_ (_41269_, _41268_, _41250_);
  nand _48433_ (_41270_, _40860_, _41251_);
  and _48434_ (_41271_, _41270_, _43634_);
  and _48435_ (_42394_, _41271_, _41269_);
  nand _48436_ (_41272_, _40806_, _39276_);
  or _48437_ (_41273_, _41262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _48438_ (_41274_, _41232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _48439_ (_41275_, _41274_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _48440_ (_41276_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _48441_ (_41277_, _41276_, _40834_);
  and _48442_ (_41278_, _41277_, _41273_);
  and _48443_ (_41279_, _40832_, _40811_);
  or _48444_ (_41280_, _41279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _48445_ (_41281_, _41279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _48446_ (_41282_, _41281_, _40871_);
  and _48447_ (_41283_, _41282_, _41280_);
  and _48448_ (_41284_, _40883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _48449_ (_41285_, _41284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _48450_ (_41286_, _40883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _48451_ (_41287_, _41286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _48452_ (_41288_, _41287_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _48453_ (_41289_, _41288_, _41285_);
  or _48454_ (_41290_, _41289_, _41283_);
  or _48455_ (_41291_, _41290_, _41278_);
  or _48456_ (_41292_, _41291_, _40806_);
  and _48457_ (_41293_, _41292_, _40869_);
  and _48458_ (_41294_, _41293_, _41272_);
  and _48459_ (_41295_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _48460_ (_41296_, _41295_, _41294_);
  and _48461_ (_42396_, _41296_, _43634_);
  nand _48462_ (_41297_, _40806_, _39268_);
  not _48463_ (_41298_, _41276_);
  nor _48464_ (_41299_, _41298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _48465_ (_41300_, _41298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _48466_ (_41301_, _41300_, _41299_);
  and _48467_ (_41302_, _41301_, _40833_);
  nor _48468_ (_41303_, _41281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _48469_ (_41304_, _41303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _48470_ (_41305_, _41303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _48471_ (_41306_, _41305_, _40872_);
  and _48472_ (_41307_, _41306_, _41304_);
  not _48473_ (_41308_, _40884_);
  and _48474_ (_41309_, _41308_, _40881_);
  or _48475_ (_41310_, _41284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _48476_ (_41311_, _41310_, _41309_);
  or _48477_ (_41312_, _41311_, _41307_);
  or _48478_ (_41313_, _41312_, _41302_);
  or _48479_ (_41314_, _41313_, _40806_);
  and _48480_ (_41315_, _41314_, _40869_);
  and _48481_ (_41316_, _41315_, _41297_);
  and _48482_ (_41317_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _48483_ (_41318_, _41317_, _41316_);
  and _48484_ (_42398_, _41318_, _43634_);
  nand _48485_ (_41319_, _40806_, _39261_);
  or _48486_ (_41320_, _40875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _48487_ (_41321_, _40876_);
  and _48488_ (_41322_, _41321_, _40872_);
  and _48489_ (_41323_, _41322_, _41320_);
  or _48490_ (_41324_, _40884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _48491_ (_41325_, _40885_);
  and _48492_ (_41326_, _41325_, _40881_);
  and _48493_ (_41327_, _41326_, _41324_);
  or _48494_ (_41328_, _40840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _48495_ (_41330_, _40890_, _40834_);
  and _48496_ (_41332_, _41330_, _41328_);
  or _48497_ (_41334_, _41332_, _41327_);
  or _48498_ (_41336_, _41334_, _41323_);
  or _48499_ (_41338_, _41336_, _40806_);
  and _48500_ (_41340_, _41338_, _40869_);
  and _48501_ (_41342_, _41340_, _41319_);
  and _48502_ (_41344_, _40846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _48503_ (_41346_, _41344_, _41342_);
  and _48504_ (_42399_, _41346_, _43634_);
  nor _48505_ (_41349_, _32442_, _28918_);
  and _48506_ (_41351_, _41349_, _33748_);
  and _48507_ (_41353_, _41351_, _39242_);
  and _48508_ (_41355_, _41353_, _31886_);
  nor _48509_ (_41357_, _41355_, _40852_);
  and _48510_ (_41359_, _41355_, _39307_);
  or _48511_ (_41361_, _41359_, _41357_);
  and _48512_ (_42401_, _41361_, _43634_);
  or _48513_ (_41364_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _48514_ (_41366_, _41364_, _43634_);
  nand _48515_ (_41368_, _40908_, _39298_);
  and _48516_ (_42402_, _41368_, _41366_);
  or _48517_ (_41371_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _48518_ (_41373_, _41371_, _43634_);
  nand _48519_ (_41375_, _40908_, _39291_);
  and _48520_ (_42404_, _41375_, _41373_);
  or _48521_ (_41378_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _48522_ (_41380_, _41378_, _43634_);
  nand _48523_ (_41381_, _40908_, _39284_);
  and _48524_ (_42406_, _41381_, _41380_);
  or _48525_ (_41382_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _48526_ (_41383_, _41382_, _43634_);
  nand _48527_ (_41384_, _40908_, _39276_);
  and _48528_ (_42407_, _41384_, _41383_);
  or _48529_ (_41385_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _48530_ (_41386_, _41385_, _43634_);
  nand _48531_ (_41387_, _40908_, _39268_);
  and _48532_ (_42409_, _41387_, _41386_);
  or _48533_ (_41388_, _40908_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _48534_ (_41389_, _41388_, _43634_);
  nand _48535_ (_41390_, _40908_, _39261_);
  and _48536_ (_42411_, _41390_, _41389_);
  nor _48537_ (_41391_, _29061_, _28918_);
  and _48538_ (_41392_, _41391_, _39934_);
  and _48539_ (_41393_, _41392_, _40094_);
  and _48540_ (_41394_, _41393_, _32463_);
  nand _48541_ (_41395_, _41394_, _32431_);
  and _48542_ (_41396_, _39244_, _32463_);
  and _48543_ (_41397_, _41396_, _40294_);
  not _48544_ (_41398_, _41397_);
  or _48545_ (_41399_, _41394_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _48546_ (_41400_, _41399_, _41398_);
  and _48547_ (_41401_, _41400_, _41395_);
  nor _48548_ (_41402_, _41398_, _39327_);
  or _48549_ (_41403_, _41402_, _41401_);
  and _48550_ (_43572_, _41403_, _43634_);
  and _48551_ (_41404_, _40696_, _28271_);
  and _48552_ (_41405_, _41404_, _40164_);
  not _48553_ (_41406_, _41405_);
  and _48554_ (_41407_, _29061_, _28929_);
  and _48555_ (_41408_, _41407_, _39934_);
  and _48556_ (_41409_, _41408_, _40094_);
  and _48557_ (_41410_, _41409_, _32463_);
  or _48558_ (_41411_, _41410_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _48559_ (_41412_, _41411_, _41406_);
  nand _48560_ (_41413_, _41410_, _32431_);
  and _48561_ (_41414_, _41413_, _41412_);
  nor _48562_ (_41415_, _41406_, _39327_);
  or _48563_ (_41416_, _41415_, _41414_);
  and _48564_ (_43575_, _41416_, _43634_);
  and _48565_ (_41417_, _41404_, _39242_);
  nor _48566_ (_41418_, _39933_, _28918_);
  and _48567_ (_41419_, _41418_, _29061_);
  and _48568_ (_41420_, _41419_, _28776_);
  and _48569_ (_41421_, _41420_, _40045_);
  nand _48570_ (_41422_, _41421_, _28250_);
  and _48571_ (_41423_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _48572_ (_41424_, _41423_, _41417_);
  or _48573_ (_41425_, _28260_, _34498_);
  and _48574_ (_41426_, _41425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _48575_ (_41427_, _41426_, _39911_);
  and _48576_ (_41428_, _41427_, _41421_);
  or _48577_ (_41429_, _41428_, _41424_);
  nand _48578_ (_41430_, _41417_, _39261_);
  and _48579_ (_41431_, _41430_, _43634_);
  and _48580_ (_43577_, _41431_, _41429_);
  not _48581_ (_41432_, _41417_);
  nor _48582_ (_41433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _48583_ (_41434_, _41433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _48584_ (_41435_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _48585_ (_41436_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _48586_ (_41437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48587_ (_41438_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _41437_);
  and _48588_ (_41439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48589_ (_41440_, _41439_, _41438_);
  nor _48590_ (_41441_, _41440_, _41436_);
  or _48591_ (_41442_, _41441_, _41435_);
  and _48592_ (_41443_, _41437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _48593_ (_41444_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _48594_ (_41445_, _41444_, _41443_);
  nor _48595_ (_41446_, _41445_, _41436_);
  and _48596_ (_41447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _41437_);
  and _48597_ (_41448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48598_ (_41449_, _41448_, _41447_);
  nand _48599_ (_41450_, _41449_, _41446_);
  or _48600_ (_41451_, _41450_, _41442_);
  and _48601_ (_41452_, _41451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _48602_ (_41453_, _41452_, _41434_);
  and _48603_ (_41454_, _39242_, _32463_);
  and _48604_ (_41455_, _41454_, _41418_);
  or _48605_ (_41456_, _41455_, _41453_);
  and _48606_ (_41457_, _41456_, _41432_);
  nand _48607_ (_41458_, _41455_, _32431_);
  and _48608_ (_41459_, _41458_, _41457_);
  nor _48609_ (_41460_, _41432_, _39327_);
  or _48610_ (_41461_, _41460_, _41459_);
  and _48611_ (_43580_, _41461_, _43634_);
  and _48612_ (_41462_, _40706_, _32507_);
  nand _48613_ (_41463_, _41462_, _32431_);
  not _48614_ (_41464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _48615_ (_41465_, _41464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _48616_ (_41466_, _41449_, _41436_);
  not _48617_ (_41467_, _41466_);
  or _48618_ (_41468_, _41467_, _41446_);
  or _48619_ (_41469_, _41468_, _41442_);
  and _48620_ (_41470_, _41469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _48621_ (_41471_, _41470_, _41465_);
  or _48622_ (_41472_, _41471_, _41462_);
  and _48623_ (_41473_, _41472_, _41432_);
  and _48624_ (_41474_, _41473_, _41463_);
  nor _48625_ (_41475_, _41432_, _39268_);
  or _48626_ (_41476_, _41475_, _41474_);
  and _48627_ (_43582_, _41476_, _43634_);
  not _48628_ (_41477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _48629_ (_41478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _41477_);
  nand _48630_ (_41479_, _41441_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _48631_ (_41480_, _41466_, _41446_);
  or _48632_ (_41481_, _41480_, _41479_);
  and _48633_ (_41482_, _41481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _48634_ (_41483_, _41482_, _41478_);
  and _48635_ (_41484_, _41418_, _39249_);
  or _48636_ (_41485_, _41484_, _41483_);
  and _48637_ (_41486_, _41485_, _41432_);
  nand _48638_ (_41487_, _41484_, _32431_);
  and _48639_ (_41488_, _41487_, _41486_);
  nor _48640_ (_41489_, _41432_, _39298_);
  or _48641_ (_41490_, _41489_, _41488_);
  and _48642_ (_43584_, _41490_, _43634_);
  and _48643_ (_41491_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _48644_ (_41492_, _41479_, _41468_);
  and _48645_ (_41493_, _41492_, _41491_);
  and _48646_ (_41494_, _41418_, _39465_);
  or _48647_ (_41500_, _41494_, _41493_);
  and _48648_ (_41506_, _41500_, _41432_);
  nand _48649_ (_41512_, _41494_, _32431_);
  and _48650_ (_41518_, _41512_, _41506_);
  nor _48651_ (_41524_, _41432_, _39284_);
  or _48652_ (_41527_, _41524_, _41518_);
  and _48653_ (_43585_, _41527_, _43634_);
  nand _48654_ (_41528_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _48655_ (_41529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _41437_);
  and _48656_ (_41530_, _41529_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _48657_ (_41531_, _41530_, _41528_);
  or _48658_ (_41532_, _41531_, _41436_);
  and _48659_ (_41533_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _48660_ (_41534_, _41533_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _48661_ (_41535_, _41534_);
  and _48662_ (_41536_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _48663_ (_41537_, _41536_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _48664_ (_41538_, _41537_);
  and _48665_ (_41539_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _48666_ (_41540_, _41539_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48667_ (_41544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _48668_ (_41547_, _41544_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _48669_ (_41551_, _41547_, _41540_);
  and _48670_ (_41552_, _41551_, _41538_);
  and _48671_ (_41553_, _41552_, _41535_);
  not _48672_ (_41555_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _48673_ (_41561_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _48674_ (_41564_, _41561_, _41555_);
  nand _48675_ (_41565_, _41564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _48676_ (_41566_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _48677_ (_41569_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _48678_ (_41575_, _41569_, _41566_);
  and _48679_ (_41577_, _41575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _48680_ (_41578_, _41577_);
  and _48681_ (_41580_, _41578_, _41565_);
  nand _48682_ (_41586_, _41580_, _41553_);
  and _48683_ (_41589_, _41586_, _41532_);
  and _48684_ (_41590_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _48685_ (_41591_, _41590_, _41437_);
  and _48686_ (_41599_, _41591_, _41589_);
  not _48687_ (_41600_, _41599_);
  not _48688_ (_41602_, _41591_);
  and _48689_ (_41603_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41436_);
  not _48690_ (_41606_, _41603_);
  not _48691_ (_41612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _48692_ (_41614_, _41536_, _41612_);
  not _48693_ (_41615_, _41614_);
  not _48694_ (_41617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48695_ (_41623_, _41539_, _41617_);
  not _48696_ (_41626_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _48697_ (_41627_, _41544_, _41626_);
  nor _48698_ (_41629_, _41627_, _41623_);
  and _48699_ (_41635_, _41629_, _41615_);
  or _48700_ (_41638_, _41635_, _41606_);
  not _48701_ (_41639_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _48702_ (_41640_, _41564_, _41639_);
  not _48703_ (_41643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _48704_ (_41650_, _41575_, _41643_);
  nor _48705_ (_41651_, _41650_, _41640_);
  not _48706_ (_41654_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _48707_ (_41655_, _41533_, _41654_);
  not _48708_ (_41661_, _41655_);
  and _48709_ (_41663_, _41661_, _41651_);
  nor _48710_ (_41664_, _41663_, _41606_);
  not _48711_ (_41666_, _41664_);
  and _48712_ (_41672_, _41666_, _41638_);
  or _48713_ (_41675_, _41672_, _41602_);
  and _48714_ (_41676_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43634_);
  and _48715_ (_41678_, _41676_, _41675_);
  and _48716_ (_43620_, _41678_, _41600_);
  nor _48717_ (_41686_, _41590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _48718_ (_41687_, _41686_);
  not _48719_ (_41688_, _41589_);
  and _48720_ (_41693_, _41672_, _41688_);
  nor _48721_ (_41698_, _41693_, _41687_);
  nand _48722_ (_41699_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43634_);
  nor _48723_ (_43622_, _41699_, _41698_);
  and _48724_ (_41704_, _41580_, _41535_);
  nand _48725_ (_41709_, _41704_, _41589_);
  or _48726_ (_41710_, _41664_, _41589_);
  and _48727_ (_41711_, _41710_, _41591_);
  and _48728_ (_41715_, _41711_, _41709_);
  or _48729_ (_41721_, _41715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _48730_ (_41722_, _41600_, _41552_);
  nor _48731_ (_41723_, _41602_, _41589_);
  not _48732_ (_41727_, _41723_);
  or _48733_ (_41732_, _41727_, _41638_);
  and _48734_ (_41733_, _41732_, _43634_);
  and _48735_ (_41734_, _41733_, _41722_);
  and _48736_ (_43624_, _41734_, _41721_);
  and _48737_ (_41735_, _41709_, _41686_);
  or _48738_ (_41736_, _41735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _48739_ (_41737_, _41686_, _41589_);
  not _48740_ (_41738_, _41737_);
  or _48741_ (_41739_, _41738_, _41552_);
  or _48742_ (_41740_, _41664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _48743_ (_41741_, _41687_, _41638_);
  and _48744_ (_41742_, _41741_, _41740_);
  or _48745_ (_41743_, _41742_, _41589_);
  and _48746_ (_41744_, _41743_, _43634_);
  and _48747_ (_41745_, _41744_, _41739_);
  and _48748_ (_43626_, _41745_, _41736_);
  nand _48749_ (_41746_, _41693_, _41436_);
  nor _48750_ (_41747_, _41437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _48751_ (_41748_, _41747_, _41590_);
  and _48752_ (_41749_, _41748_, _43634_);
  and _48753_ (_43628_, _41749_, _41746_);
  and _48754_ (_41750_, _41693_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _48755_ (_41751_, _41437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _48756_ (_41752_, _41751_, _41747_);
  nor _48757_ (_41753_, _41752_, _41688_);
  or _48758_ (_41754_, _41753_, _41590_);
  or _48759_ (_41755_, _41754_, _41750_);
  not _48760_ (_41756_, _41590_);
  or _48761_ (_41757_, _41752_, _41756_);
  and _48762_ (_41758_, _41757_, _43634_);
  and _48763_ (_43630_, _41758_, _41755_);
  and _48764_ (_41759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43634_);
  and _48765_ (_43632_, _41759_, _41590_);
  nor _48766_ (_43637_, _41433_, rst);
  and _48767_ (_43638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _43634_);
  nor _48768_ (_41760_, _41693_, _41590_);
  and _48769_ (_41761_, _41590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _48770_ (_41762_, _41761_, _41760_);
  and _48771_ (_00137_, _41762_, _43634_);
  and _48772_ (_41763_, _41590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _48773_ (_41764_, _41763_, _41760_);
  and _48774_ (_00139_, _41764_, _43634_);
  and _48775_ (_41765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _43634_);
  and _48776_ (_00141_, _41765_, _41590_);
  not _48777_ (_41766_, _41627_);
  nor _48778_ (_41767_, _41650_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _48779_ (_41768_, _41767_, _41640_);
  or _48780_ (_41769_, _41768_, _41655_);
  and _48781_ (_41770_, _41769_, _41766_);
  or _48782_ (_41771_, _41770_, _41623_);
  nor _48783_ (_41772_, _41672_, _41589_);
  and _48784_ (_41773_, _41772_, _41615_);
  and _48785_ (_41774_, _41773_, _41771_);
  not _48786_ (_41775_, _41547_);
  or _48787_ (_41776_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48788_ (_41777_, _41776_, _41565_);
  or _48789_ (_41778_, _41777_, _41534_);
  and _48790_ (_41779_, _41778_, _41775_);
  or _48791_ (_41780_, _41779_, _41540_);
  and _48792_ (_41781_, _41589_, _41538_);
  and _48793_ (_41782_, _41781_, _41780_);
  or _48794_ (_41783_, _41782_, _41590_);
  or _48795_ (_41784_, _41783_, _41774_);
  or _48796_ (_41785_, _41756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48797_ (_41786_, _41785_, _43634_);
  and _48798_ (_00143_, _41786_, _41784_);
  nor _48799_ (_41787_, _41623_, _41614_);
  or _48800_ (_41788_, _41655_, _41627_);
  and _48801_ (_41789_, _41651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48802_ (_41790_, _41789_, _41788_);
  and _48803_ (_41791_, _41790_, _41787_);
  and _48804_ (_41792_, _41791_, _41772_);
  not _48805_ (_41793_, _41540_);
  or _48806_ (_41794_, _41547_, _41534_);
  and _48807_ (_41795_, _41580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48808_ (_41796_, _41795_, _41794_);
  and _48809_ (_41797_, _41796_, _41793_);
  and _48810_ (_41798_, _41797_, _41781_);
  or _48811_ (_41799_, _41798_, _41590_);
  or _48812_ (_41800_, _41799_, _41792_);
  or _48813_ (_41801_, _41756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _48814_ (_41802_, _41801_, _43634_);
  and _48815_ (_00145_, _41802_, _41800_);
  and _48816_ (_41803_, _41661_, _41603_);
  nand _48817_ (_41804_, _41803_, _41635_);
  or _48818_ (_41805_, _41804_, _41651_);
  nor _48819_ (_41806_, _41805_, _41589_);
  nand _48820_ (_41807_, _41553_, _41532_);
  nor _48821_ (_41808_, _41807_, _41580_);
  or _48822_ (_41809_, _41808_, _41590_);
  or _48823_ (_41810_, _41809_, _41806_);
  or _48824_ (_41811_, _41756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _48825_ (_41812_, _41811_, _43634_);
  and _48826_ (_00146_, _41812_, _41810_);
  and _48827_ (_41813_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _43634_);
  and _48828_ (_00148_, _41813_, _41590_);
  and _48829_ (_41814_, _41590_, _41437_);
  or _48830_ (_41815_, _41814_, _41698_);
  or _48831_ (_41816_, _41815_, _41723_);
  and _48832_ (_00150_, _41816_, _43634_);
  not _48833_ (_41817_, _41760_);
  and _48834_ (_41818_, _41817_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _48835_ (_41819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _48836_ (_41820_, _41577_, _41437_);
  or _48837_ (_41821_, _41820_, _41819_);
  nor _48838_ (_41822_, _41565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48839_ (_41823_, _41822_, _41534_);
  nand _48840_ (_41824_, _41823_, _41821_);
  or _48841_ (_41825_, _41535_, _41439_);
  and _48842_ (_41826_, _41825_, _41824_);
  or _48843_ (_41827_, _41826_, _41547_);
  or _48844_ (_41829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _41437_);
  or _48845_ (_41830_, _41829_, _41775_);
  and _48846_ (_41832_, _41830_, _41793_);
  and _48847_ (_41833_, _41832_, _41827_);
  and _48848_ (_41835_, _41540_, _41439_);
  or _48849_ (_41836_, _41835_, _41537_);
  or _48850_ (_41838_, _41836_, _41833_);
  or _48851_ (_41839_, _41829_, _41538_);
  and _48852_ (_41841_, _41839_, _41589_);
  and _48853_ (_41842_, _41841_, _41838_);
  and _48854_ (_41844_, _41650_, _41437_);
  or _48855_ (_41845_, _41844_, _41819_);
  and _48856_ (_41847_, _41640_, _41437_);
  nor _48857_ (_41848_, _41847_, _41655_);
  nand _48858_ (_41850_, _41848_, _41845_);
  or _48859_ (_41851_, _41661_, _41439_);
  and _48860_ (_41853_, _41851_, _41850_);
  or _48861_ (_41854_, _41853_, _41627_);
  not _48862_ (_41856_, _41623_);
  or _48863_ (_41857_, _41829_, _41766_);
  and _48864_ (_41858_, _41857_, _41856_);
  and _48865_ (_41859_, _41858_, _41854_);
  and _48866_ (_41860_, _41623_, _41439_);
  or _48867_ (_41861_, _41860_, _41614_);
  or _48868_ (_41862_, _41861_, _41859_);
  and _48869_ (_41863_, _41829_, _41772_);
  or _48870_ (_41864_, _41863_, _41773_);
  and _48871_ (_41865_, _41864_, _41862_);
  or _48872_ (_41866_, _41865_, _41842_);
  and _48873_ (_41867_, _41866_, _41756_);
  or _48874_ (_41868_, _41867_, _41818_);
  and _48875_ (_00152_, _41868_, _43634_);
  or _48876_ (_41869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _41437_);
  and _48877_ (_41870_, _41869_, _41538_);
  or _48878_ (_41871_, _41870_, _41552_);
  or _48879_ (_41872_, _41820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48880_ (_41873_, _41872_, _41823_);
  nand _48881_ (_41874_, _41534_, _41448_);
  nand _48882_ (_41875_, _41874_, _41551_);
  or _48883_ (_41876_, _41875_, _41873_);
  and _48884_ (_41877_, _41876_, _41871_);
  nand _48885_ (_41878_, _41537_, _41448_);
  nand _48886_ (_41879_, _41878_, _41589_);
  or _48887_ (_41880_, _41879_, _41877_);
  not _48888_ (_41881_, _41629_);
  and _48889_ (_41882_, _41869_, _41881_);
  or _48890_ (_41883_, _41844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48891_ (_41884_, _41848_, _41629_);
  and _48892_ (_41885_, _41884_, _41883_);
  or _48893_ (_41886_, _41885_, _41882_);
  and _48894_ (_41887_, _41886_, _41615_);
  and _48895_ (_41888_, _41655_, _41629_);
  or _48896_ (_41889_, _41888_, _41614_);
  and _48897_ (_41890_, _41889_, _41448_);
  or _48898_ (_41891_, _41890_, _41672_);
  or _48899_ (_41892_, _41891_, _41589_);
  or _48900_ (_41893_, _41892_, _41887_);
  and _48901_ (_41894_, _41893_, _41880_);
  or _48902_ (_41895_, _41894_, _41590_);
  or _48903_ (_41896_, _41760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48904_ (_41897_, _41896_, _43634_);
  and _48905_ (_00154_, _41897_, _41895_);
  and _48906_ (_41898_, _41817_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _48907_ (_41899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48908_ (_41900_, _41899_, _41538_);
  and _48909_ (_41901_, _41900_, _41589_);
  not _48910_ (_41902_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _48911_ (_41903_, _41577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48912_ (_41904_, _41903_, _41902_);
  nor _48913_ (_41905_, _41565_, _41437_);
  nor _48914_ (_41906_, _41905_, _41534_);
  nand _48915_ (_41907_, _41906_, _41904_);
  or _48916_ (_41908_, _41535_, _41438_);
  and _48917_ (_41909_, _41908_, _41907_);
  or _48918_ (_41910_, _41909_, _41547_);
  or _48919_ (_41911_, _41899_, _41775_);
  and _48920_ (_41912_, _41911_, _41793_);
  and _48921_ (_41913_, _41912_, _41910_);
  and _48922_ (_41914_, _41540_, _41438_);
  or _48923_ (_41915_, _41914_, _41537_);
  or _48924_ (_41916_, _41915_, _41913_);
  and _48925_ (_41917_, _41916_, _41901_);
  or _48926_ (_41918_, _41899_, _41615_);
  and _48927_ (_41919_, _41650_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48928_ (_41920_, _41919_, _41902_);
  and _48929_ (_41921_, _41640_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48930_ (_41922_, _41921_, _41655_);
  nand _48931_ (_41923_, _41922_, _41920_);
  or _48932_ (_41924_, _41661_, _41438_);
  and _48933_ (_41925_, _41924_, _41923_);
  or _48934_ (_41926_, _41925_, _41627_);
  or _48935_ (_41927_, _41899_, _41766_);
  and _48936_ (_41928_, _41927_, _41856_);
  and _48937_ (_41929_, _41928_, _41926_);
  and _48938_ (_41930_, _41623_, _41438_);
  or _48939_ (_41931_, _41930_, _41614_);
  or _48940_ (_41932_, _41931_, _41929_);
  and _48941_ (_41933_, _41932_, _41772_);
  and _48942_ (_41934_, _41933_, _41918_);
  or _48943_ (_41935_, _41934_, _41917_);
  and _48944_ (_41936_, _41935_, _41756_);
  or _48945_ (_41937_, _41936_, _41898_);
  and _48946_ (_00156_, _41937_, _43634_);
  or _48947_ (_41938_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48948_ (_41939_, _41938_, _41538_);
  or _48949_ (_41940_, _41939_, _41552_);
  or _48950_ (_41941_, _41903_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48951_ (_41942_, _41941_, _41906_);
  nand _48952_ (_41943_, _41534_, _41447_);
  nand _48953_ (_41944_, _41943_, _41551_);
  or _48954_ (_41945_, _41944_, _41942_);
  and _48955_ (_41946_, _41945_, _41940_);
  nand _48956_ (_41947_, _41537_, _41447_);
  nand _48957_ (_41948_, _41947_, _41589_);
  or _48958_ (_41949_, _41948_, _41946_);
  and _48959_ (_41950_, _41938_, _41881_);
  or _48960_ (_41951_, _41919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48961_ (_41952_, _41922_, _41629_);
  and _48962_ (_41953_, _41952_, _41951_);
  or _48963_ (_41954_, _41953_, _41950_);
  and _48964_ (_41955_, _41954_, _41615_);
  and _48965_ (_41956_, _41889_, _41447_);
  or _48966_ (_41957_, _41956_, _41672_);
  or _48967_ (_41958_, _41957_, _41589_);
  or _48968_ (_41959_, _41958_, _41955_);
  and _48969_ (_41960_, _41959_, _41949_);
  or _48970_ (_41961_, _41960_, _41590_);
  or _48971_ (_41962_, _41760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48972_ (_41963_, _41962_, _43634_);
  and _48973_ (_00157_, _41963_, _41961_);
  or _48974_ (_41964_, _41687_, _41672_);
  and _48975_ (_41965_, _41964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _48976_ (_41966_, _41965_, _41737_);
  and _48977_ (_00159_, _41966_, _43634_);
  and _48978_ (_41967_, _41675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _48979_ (_41968_, _41967_, _41599_);
  and _48980_ (_00161_, _41968_, _43634_);
  and _48981_ (_41969_, _41421_, _28271_);
  or _48982_ (_41970_, _41969_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _48983_ (_41971_, _41970_, _41432_);
  nand _48984_ (_41972_, _41969_, _32431_);
  and _48985_ (_41973_, _41972_, _41971_);
  and _48986_ (_41974_, _41417_, _39307_);
  or _48987_ (_41975_, _41974_, _41973_);
  and _48988_ (_00163_, _41975_, _43634_);
  and _48989_ (_41976_, _41421_, _34509_);
  or _48990_ (_41977_, _41976_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _48991_ (_41978_, _41977_, _41432_);
  nand _48992_ (_41979_, _41976_, _32431_);
  and _48993_ (_41980_, _41979_, _41978_);
  nor _48994_ (_41981_, _41432_, _39291_);
  or _48995_ (_41982_, _41981_, _41980_);
  and _48996_ (_00165_, _41982_, _43634_);
  and _48997_ (_41983_, _41421_, _35978_);
  or _48998_ (_41984_, _41983_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _48999_ (_41985_, _41984_, _41432_);
  nand _49000_ (_41986_, _41983_, _32431_);
  and _49001_ (_41987_, _41986_, _41985_);
  nor _49002_ (_41988_, _41432_, _39276_);
  or _49003_ (_41989_, _41988_, _41987_);
  and _49004_ (_00167_, _41989_, _43634_);
  and _49005_ (_41990_, _41409_, _28271_);
  or _49006_ (_41991_, _41990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _49007_ (_41992_, _41991_, _41406_);
  nand _49008_ (_41993_, _41990_, _32431_);
  and _49009_ (_41994_, _41993_, _41992_);
  and _49010_ (_41995_, _41405_, _39307_);
  or _49011_ (_41996_, _41995_, _41994_);
  and _49012_ (_00168_, _41996_, _43634_);
  and _49013_ (_41997_, _41409_, _39768_);
  or _49014_ (_41998_, _41997_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _49015_ (_41999_, _41998_, _41406_);
  nand _49016_ (_42000_, _41997_, _32431_);
  and _49017_ (_42001_, _42000_, _41999_);
  nor _49018_ (_42002_, _41406_, _39298_);
  or _49019_ (_42003_, _42002_, _42001_);
  and _49020_ (_00170_, _42003_, _43634_);
  nand _49021_ (_42004_, _41409_, _40329_);
  and _49022_ (_42005_, _42004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _49023_ (_42006_, _42005_, _41405_);
  and _49024_ (_42007_, _34542_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _49025_ (_42008_, _42007_, _34531_);
  and _49026_ (_42009_, _42008_, _41409_);
  or _49027_ (_42010_, _42009_, _42006_);
  nand _49028_ (_42011_, _41405_, _39291_);
  and _49029_ (_42012_, _42011_, _43634_);
  and _49030_ (_00172_, _42012_, _42010_);
  and _49031_ (_42013_, _41409_, _35217_);
  or _49032_ (_42014_, _42013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _49033_ (_42015_, _42014_, _41406_);
  nand _49034_ (_42016_, _42013_, _32431_);
  and _49035_ (_42017_, _42016_, _42015_);
  nor _49036_ (_42018_, _41406_, _39284_);
  or _49037_ (_42019_, _42018_, _42017_);
  and _49038_ (_00174_, _42019_, _43634_);
  and _49039_ (_42020_, _41409_, _35978_);
  or _49040_ (_42021_, _42020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _49041_ (_42022_, _42021_, _41406_);
  nand _49042_ (_42023_, _42020_, _32431_);
  and _49043_ (_42024_, _42023_, _42022_);
  nor _49044_ (_42025_, _41406_, _39276_);
  or _49045_ (_42026_, _42025_, _42024_);
  and _49046_ (_00176_, _42026_, _43634_);
  and _49047_ (_42027_, _41409_, _36762_);
  or _49048_ (_42028_, _42027_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _49049_ (_42029_, _42028_, _41406_);
  nand _49050_ (_42030_, _42027_, _32431_);
  and _49051_ (_42031_, _42030_, _42029_);
  nor _49052_ (_42032_, _41406_, _39268_);
  or _49053_ (_42033_, _42032_, _42031_);
  and _49054_ (_00178_, _42033_, _43634_);
  and _49055_ (_42034_, _41409_, _37502_);
  or _49056_ (_42035_, _42034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _49057_ (_42036_, _42035_, _41406_);
  nand _49058_ (_42037_, _42034_, _32431_);
  and _49059_ (_42038_, _42037_, _42036_);
  nor _49060_ (_42039_, _41406_, _39261_);
  or _49061_ (_42040_, _42039_, _42038_);
  and _49062_ (_00180_, _42040_, _43634_);
  and _49063_ (_42041_, _41393_, _28271_);
  nand _49064_ (_42042_, _42041_, _32431_);
  or _49065_ (_42043_, _42041_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _49066_ (_42044_, _42043_, _41398_);
  and _49067_ (_42045_, _42044_, _42042_);
  and _49068_ (_42046_, _41397_, _39307_);
  or _49069_ (_42047_, _42046_, _42045_);
  and _49070_ (_00181_, _42047_, _43634_);
  and _49071_ (_42048_, _41393_, _39768_);
  nand _49072_ (_42049_, _42048_, _32431_);
  or _49073_ (_42050_, _42048_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _49074_ (_42051_, _42050_, _41398_);
  and _49075_ (_42052_, _42051_, _42049_);
  nor _49076_ (_42053_, _41398_, _39298_);
  or _49077_ (_42054_, _42053_, _42052_);
  and _49078_ (_00183_, _42054_, _43634_);
  and _49079_ (_42055_, _34542_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _49080_ (_42056_, _42055_, _34531_);
  and _49081_ (_42057_, _42056_, _41393_);
  nand _49082_ (_42058_, _41393_, _40329_);
  and _49083_ (_42059_, _42058_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _49084_ (_42060_, _42059_, _41397_);
  or _49085_ (_42061_, _42060_, _42057_);
  nand _49086_ (_42062_, _41397_, _39291_);
  and _49087_ (_42063_, _42062_, _43634_);
  and _49088_ (_00185_, _42063_, _42061_);
  and _49089_ (_42064_, _41393_, _35217_);
  nand _49090_ (_42065_, _42064_, _32431_);
  or _49091_ (_42066_, _42064_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _49092_ (_42067_, _42066_, _41398_);
  and _49093_ (_42068_, _42067_, _42065_);
  nor _49094_ (_42069_, _41398_, _39284_);
  or _49095_ (_42070_, _42069_, _42068_);
  and _49096_ (_00187_, _42070_, _43634_);
  and _49097_ (_42071_, _41393_, _35978_);
  nand _49098_ (_42072_, _42071_, _32431_);
  or _49099_ (_42073_, _42071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _49100_ (_42074_, _42073_, _41398_);
  and _49101_ (_42075_, _42074_, _42072_);
  nor _49102_ (_42076_, _41398_, _39276_);
  or _49103_ (_42077_, _42076_, _42075_);
  and _49104_ (_00189_, _42077_, _43634_);
  and _49105_ (_42078_, _41393_, _36762_);
  nand _49106_ (_42079_, _42078_, _32431_);
  or _49107_ (_42080_, _42078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _49108_ (_42081_, _42080_, _41398_);
  and _49109_ (_42082_, _42081_, _42079_);
  nor _49110_ (_42083_, _41398_, _39268_);
  or _49111_ (_42084_, _42083_, _42082_);
  and _49112_ (_00191_, _42084_, _43634_);
  and _49113_ (_42085_, _41393_, _37502_);
  nand _49114_ (_42086_, _42085_, _32431_);
  or _49115_ (_42087_, _42085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _49116_ (_42088_, _42087_, _42086_);
  or _49117_ (_42089_, _42088_, _41397_);
  nand _49118_ (_42090_, _41397_, _39261_);
  and _49119_ (_42091_, _42090_, _43634_);
  and _49120_ (_00192_, _42091_, _42089_);
  and _49121_ (_42092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _49122_ (_42093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _49123_ (_42094_, _41433_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _49124_ (_42095_, _42094_, _42093_);
  not _49125_ (_42096_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _49126_ (_42097_, _42096_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _49127_ (_42098_, _42097_, _42095_);
  nor _49128_ (_42099_, _42098_, _42092_);
  or _49129_ (_42100_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _49130_ (_42101_, _42100_, _43634_);
  nor _49131_ (_00552_, _42101_, _42099_);
  nor _49132_ (_42102_, _42099_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _49133_ (_42103_, _42102_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _49134_ (_42104_, _42102_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _49135_ (_42105_, _42104_, _43634_);
  and _49136_ (_00555_, _42105_, _42103_);
  not _49137_ (_42106_, rxd_i);
  and _49138_ (_42107_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _42106_);
  nor _49139_ (_42108_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _49140_ (_42109_, _42108_);
  and _49141_ (_42110_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _49142_ (_42111_, _42110_, _42109_);
  and _49143_ (_42112_, _42111_, _42107_);
  not _49144_ (_42113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _49145_ (_42114_, _42113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _49146_ (_42115_, _42114_, _42108_);
  or _49147_ (_42116_, _42115_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _49148_ (_42117_, _42116_, _42112_);
  and _49149_ (_42118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _43634_);
  and _49150_ (_00558_, _42118_, _42117_);
  and _49151_ (_42119_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _49152_ (_42120_, _42119_, _42109_);
  nor _49153_ (_42121_, _42108_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _49154_ (_42122_, _42121_, _42113_);
  nor _49155_ (_42123_, _42122_, _42120_);
  not _49156_ (_42124_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _49157_ (_42125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _42124_);
  not _49158_ (_42126_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _49159_ (_42127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _42126_);
  and _49160_ (_42128_, _42127_, _42125_);
  not _49161_ (_42129_, _42128_);
  or _49162_ (_42130_, _42129_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _49163_ (_42131_, _42128_, _42120_);
  and _49164_ (_42132_, _42120_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49165_ (_42133_, _42132_, _42131_);
  and _49166_ (_42134_, _42133_, _42130_);
  or _49167_ (_42135_, _42134_, _42123_);
  and _49168_ (_42136_, _42108_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _49169_ (_42137_, _42136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _49170_ (_42138_, _42137_);
  or _49171_ (_42139_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _49172_ (_42140_, _42139_, _42135_);
  nand _49173_ (_00561_, _42140_, _42118_);
  not _49174_ (_42141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _49175_ (_42142_, _42120_);
  nor _49176_ (_42143_, _42113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _49177_ (_42144_, _42143_);
  not _49178_ (_42145_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _49179_ (_42146_, _42108_, _42145_);
  and _49180_ (_42147_, _42146_, _42144_);
  and _49181_ (_42148_, _42147_, _42142_);
  nor _49182_ (_42149_, _42148_, _42141_);
  and _49183_ (_42150_, _42148_, rxd_i);
  or _49184_ (_42151_, _42150_, rst);
  or _49185_ (_00563_, _42151_, _42149_);
  nor _49186_ (_42152_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _49187_ (_42153_, _42152_, _42125_);
  and _49188_ (_42154_, _42153_, _42132_);
  nand _49189_ (_42155_, _42154_, _42106_);
  or _49190_ (_42156_, _42154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _49191_ (_42157_, _42156_, _43634_);
  and _49192_ (_00566_, _42157_, _42155_);
  and _49193_ (_42158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _49194_ (_42159_, _42158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _49195_ (_42160_, _42159_, _42124_);
  and _49196_ (_42161_, _42160_, _42132_);
  and _49197_ (_42162_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _49198_ (_42163_, _42162_, _42132_);
  nor _49199_ (_42164_, _42159_, _42142_);
  or _49200_ (_42165_, _42164_, _42163_);
  and _49201_ (_42166_, _42165_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _49202_ (_42167_, _42166_, _42161_);
  and _49203_ (_00569_, _42167_, _43634_);
  and _49204_ (_42168_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _43634_);
  nand _49205_ (_42169_, _42168_, _42145_);
  nand _49206_ (_42170_, _42118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _49207_ (_00571_, _42170_, _42169_);
  and _49208_ (_42171_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _42145_);
  not _49209_ (_42172_, _42111_);
  not _49210_ (_42173_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _49211_ (_42174_, _42115_, _42173_);
  and _49212_ (_42175_, _42174_, _42172_);
  and _49213_ (_42176_, _42175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _49214_ (_42177_, _42176_, _42120_);
  or _49215_ (_42178_, _42128_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _49216_ (_42179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _49217_ (_42180_, _42179_, _42131_);
  and _49218_ (_42181_, _42180_, _42178_);
  and _49219_ (_42182_, _42181_, _42177_);
  or _49220_ (_42183_, _42182_, _42137_);
  nand _49221_ (_42184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _49222_ (_42185_, _42184_, _42120_);
  or _49223_ (_42186_, _42185_, _42129_);
  and _49224_ (_42187_, _42186_, _42138_);
  or _49225_ (_42188_, _42187_, rxd_i);
  and _49226_ (_42189_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _49227_ (_42190_, _42189_, _42183_);
  or _49228_ (_42191_, _42190_, _42171_);
  and _49229_ (_00574_, _42191_, _43634_);
  and _49230_ (_42192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _49231_ (_42193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _49232_ (_42194_, _42094_, _42193_);
  or _49233_ (_42195_, _42194_, _42097_);
  nor _49234_ (_42196_, _42195_, _42192_);
  or _49235_ (_42197_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _49236_ (_42198_, _42197_, _43634_);
  nor _49237_ (_00577_, _42198_, _42196_);
  nor _49238_ (_42199_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _49239_ (_42200_, _42199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _49240_ (_42201_, _42199_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _49241_ (_42202_, _42201_, _43634_);
  and _49242_ (_00579_, _42202_, _42200_);
  not _49243_ (_42203_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _49244_ (_42204_, _41351_, _31886_);
  and _49245_ (_42205_, _42204_, _40067_);
  and _49246_ (_42206_, _42205_, _43634_);
  nand _49247_ (_42207_, _42206_, _42203_);
  and _49248_ (_42208_, _42136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _49249_ (_42209_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _49250_ (_42210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _49251_ (_42211_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _49252_ (_42212_, _42211_, _42210_);
  and _49253_ (_42213_, _42212_, _42209_);
  not _49254_ (_42214_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _49255_ (_42215_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _49256_ (_42216_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _49257_ (_42217_, _42216_, _42215_);
  and _49258_ (_42218_, _42217_, _42214_);
  and _49259_ (_42219_, _42218_, _42213_);
  or _49260_ (_42220_, _42219_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _49261_ (_42221_, _42219_, _42203_);
  nand _49262_ (_42222_, _42221_, _42220_);
  nand _49263_ (_42223_, _42222_, _42208_);
  nor _49264_ (_42224_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _49265_ (_42225_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _49266_ (_42226_, _42225_, _42224_);
  and _49267_ (_42227_, _42109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _49268_ (_42228_, _42227_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _49269_ (_42229_, _42228_, _42226_);
  not _49270_ (_42230_, _42229_);
  or _49271_ (_42231_, _42230_, _42220_);
  and _49272_ (_42232_, _42226_, _42227_);
  not _49273_ (_42233_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or _49274_ (_42234_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _42233_);
  or _49275_ (_42235_, _42234_, _42232_);
  or _49276_ (_42236_, _42235_, _42208_);
  and _49277_ (_42237_, _42236_, _42231_);
  nand _49278_ (_42238_, _42237_, _42223_);
  nor _49279_ (_42239_, _42205_, rst);
  nand _49280_ (_42240_, _42239_, _42238_);
  and _49281_ (_00582_, _42240_, _42207_);
  not _49282_ (_42241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and _49283_ (_42242_, _42219_, _42241_);
  nand _49284_ (_42243_, _42232_, _42242_);
  and _49285_ (_42244_, _42219_, _42208_);
  or _49286_ (_42245_, _42233_, rst);
  nor _49287_ (_42246_, _42245_, _42244_);
  and _49288_ (_42247_, _42246_, _42243_);
  or _49289_ (_00585_, _42247_, _42206_);
  or _49290_ (_42248_, _42230_, _42242_);
  or _49291_ (_42249_, _42232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _49292_ (_42250_, _42136_, _42233_);
  and _49293_ (_42251_, _42250_, _42249_);
  and _49294_ (_42252_, _42251_, _42248_);
  or _49295_ (_42253_, _42252_, _42244_);
  and _49296_ (_00587_, _42253_, _42239_);
  and _49297_ (_42254_, _42228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _49298_ (_42255_, _42254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _49299_ (_42256_, _42255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _49300_ (_42257_, _42256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _49301_ (_42258_, _42256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _49302_ (_42259_, _42258_, _42257_);
  and _49303_ (_00590_, _42259_, _42239_);
  nor _49304_ (_42260_, _42229_, _42208_);
  and _49305_ (_42261_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _49306_ (_42262_, _42261_, _42239_);
  and _49307_ (_42263_, _42206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _49308_ (_00593_, _42263_, _42262_);
  and _49309_ (_42264_, _41396_, _39242_);
  or _49310_ (_42265_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _49311_ (_42266_, _42265_, _43634_);
  nand _49312_ (_42267_, _42264_, _39327_);
  and _49313_ (_00595_, _42267_, _42266_);
  and _49314_ (_42268_, _41392_, _40045_);
  and _49315_ (_42269_, _42268_, _32463_);
  nand _49316_ (_42270_, _42269_, _32431_);
  and _49317_ (_42271_, _41404_, _40067_);
  not _49318_ (_42272_, _42271_);
  or _49319_ (_42273_, _42269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _49320_ (_42274_, _42273_, _42272_);
  and _49321_ (_42275_, _42274_, _42270_);
  nor _49322_ (_42276_, _42272_, _39327_);
  or _49323_ (_42277_, _42276_, _42275_);
  and _49324_ (_00598_, _42277_, _43634_);
  nor _49325_ (_42278_, _42137_, _42131_);
  not _49326_ (_42279_, _42278_);
  nor _49327_ (_42280_, _42175_, _42120_);
  nor _49328_ (_42281_, _42280_, _42279_);
  nor _49329_ (_42282_, _42281_, _42145_);
  or _49330_ (_42283_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _49331_ (_42284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _42145_);
  or _49332_ (_42285_, _42284_, _42278_);
  and _49333_ (_42286_, _42285_, _43634_);
  and _49334_ (_01218_, _42286_, _42283_);
  or _49335_ (_42287_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _49336_ (_42288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _42145_);
  or _49337_ (_42289_, _42288_, _42278_);
  and _49338_ (_42290_, _42289_, _43634_);
  and _49339_ (_01220_, _42290_, _42287_);
  or _49340_ (_42291_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _49341_ (_42292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _42145_);
  or _49342_ (_42293_, _42292_, _42278_);
  and _49343_ (_42294_, _42293_, _43634_);
  and _49344_ (_01222_, _42294_, _42291_);
  or _49345_ (_42295_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _49346_ (_42296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _42145_);
  or _49347_ (_42297_, _42296_, _42278_);
  and _49348_ (_42298_, _42297_, _43634_);
  and _49349_ (_01224_, _42298_, _42295_);
  or _49350_ (_42299_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _49351_ (_42300_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _42145_);
  or _49352_ (_42301_, _42300_, _42278_);
  and _49353_ (_42302_, _42301_, _43634_);
  and _49354_ (_01226_, _42302_, _42299_);
  or _49355_ (_42303_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _49356_ (_42304_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _42145_);
  or _49357_ (_42305_, _42304_, _42278_);
  and _49358_ (_42306_, _42305_, _43634_);
  and _49359_ (_01228_, _42306_, _42303_);
  or _49360_ (_42307_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _49361_ (_42308_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _42145_);
  or _49362_ (_42309_, _42308_, _42278_);
  and _49363_ (_42310_, _42309_, _43634_);
  and _49364_ (_01230_, _42310_, _42307_);
  or _49365_ (_42311_, _42282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _49366_ (_42312_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _42145_);
  or _49367_ (_42313_, _42312_, _42278_);
  and _49368_ (_42314_, _42313_, _43634_);
  and _49369_ (_01232_, _42314_, _42311_);
  nor _49370_ (_42315_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _49371_ (_42316_, _42315_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _49372_ (_42317_, _42129_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _49373_ (_42318_, _42128_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _49374_ (_42319_, _42318_, _42120_);
  and _49375_ (_42320_, _42319_, _42317_);
  or _49376_ (_42321_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _49377_ (_42322_, _42321_, _42174_);
  and _49378_ (_42323_, _42322_, _42142_);
  or _49379_ (_42324_, _42323_, _42320_);
  or _49380_ (_42325_, _42324_, _42137_);
  or _49381_ (_42326_, _42138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _49382_ (_42327_, _42326_, _42118_);
  and _49383_ (_42328_, _42327_, _42325_);
  or _49384_ (_01234_, _42328_, _42316_);
  and _49385_ (_42329_, _42128_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _49386_ (_42330_, _42329_, _42175_);
  or _49387_ (_42331_, _42330_, _42281_);
  and _49388_ (_42332_, _42331_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _49389_ (_42333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _42145_);
  nand _49390_ (_42334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _49391_ (_42335_, _42334_, _42278_);
  or _49392_ (_42336_, _42335_, _42333_);
  or _49393_ (_42337_, _42336_, _42332_);
  and _49394_ (_01236_, _42337_, _43634_);
  not _49395_ (_42338_, _42282_);
  and _49396_ (_42339_, _42338_, _42168_);
  or _49397_ (_42340_, _42330_, _42279_);
  and _49398_ (_42341_, _42118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _49399_ (_42342_, _42341_, _42340_);
  or _49400_ (_01238_, _42342_, _42339_);
  or _49401_ (_42343_, _42161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _49402_ (_42344_, _42161_, _42106_);
  and _49403_ (_42345_, _42344_, _43634_);
  and _49404_ (_01240_, _42345_, _42343_);
  or _49405_ (_42346_, _42163_, _42126_);
  or _49406_ (_42347_, _42132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _49407_ (_42348_, _42347_, _43634_);
  and _49408_ (_01242_, _42348_, _42346_);
  and _49409_ (_42349_, _42163_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _49410_ (_42350_, _42152_, _42158_);
  and _49411_ (_42351_, _42350_, _42132_);
  or _49412_ (_42353_, _42351_, _42349_);
  and _49413_ (_01244_, _42353_, _43634_);
  and _49414_ (_42356_, _42165_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _49415_ (_42358_, _42158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _49416_ (_42360_, _42358_, _42164_);
  or _49417_ (_42362_, _42360_, _42356_);
  and _49418_ (_01245_, _42362_, _43634_);
  and _49419_ (_42365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _42145_);
  and _49420_ (_42367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49421_ (_42369_, _42367_, _42365_);
  and _49422_ (_01247_, _42369_, _43634_);
  and _49423_ (_42372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _42145_);
  and _49424_ (_42374_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49425_ (_42376_, _42374_, _42372_);
  and _49426_ (_01249_, _42376_, _43634_);
  and _49427_ (_42379_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _42145_);
  and _49428_ (_42381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49429_ (_42383_, _42381_, _42379_);
  and _49430_ (_01251_, _42383_, _43634_);
  and _49431_ (_42386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _42145_);
  and _49432_ (_42388_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49433_ (_42390_, _42388_, _42386_);
  and _49434_ (_01253_, _42390_, _43634_);
  and _49435_ (_42393_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _42145_);
  and _49436_ (_42395_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49437_ (_42397_, _42395_, _42393_);
  and _49438_ (_01255_, _42397_, _43634_);
  and _49439_ (_42400_, _42118_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _49440_ (_01257_, _42400_, _42316_);
  and _49441_ (_42403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _49442_ (_42405_, _42403_, _42333_);
  and _49443_ (_01259_, _42405_, _43634_);
  nor _49444_ (_42408_, _42228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _49445_ (_42410_, _42408_, _42254_);
  and _49446_ (_01261_, _42410_, _42239_);
  nor _49447_ (_42412_, _42254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _49448_ (_42413_, _42412_, _42255_);
  and _49449_ (_01263_, _42413_, _42239_);
  nor _49450_ (_42414_, _42255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _49451_ (_42415_, _42414_, _42256_);
  and _49452_ (_01265_, _42415_, _42239_);
  and _49453_ (_42416_, _42229_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _49454_ (_42417_, _42208_, _42241_);
  nor _49455_ (_42418_, _42417_, _42229_);
  or _49456_ (_42419_, _42418_, _42416_);
  and _49457_ (_42420_, _42219_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _49458_ (_42421_, _42420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _49459_ (_42422_, _42421_, _42208_);
  nor _49460_ (_42423_, _42422_, _42419_);
  nor _49461_ (_42424_, _42423_, _42205_);
  nor _49462_ (_42425_, _42109_, _39306_);
  and _49463_ (_42426_, _42425_, _42205_);
  or _49464_ (_42427_, _42426_, _42424_);
  and _49465_ (_01267_, _42427_, _43634_);
  not _49466_ (_42428_, _42260_);
  and _49467_ (_42429_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _49468_ (_42430_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _49469_ (_42431_, _42430_, _42429_);
  and _49470_ (_42432_, _42431_, _42239_);
  nand _49471_ (_42433_, _42108_, _39298_);
  nand _49472_ (_42434_, _42109_, _39306_);
  and _49473_ (_42435_, _42434_, _42206_);
  and _49474_ (_42436_, _42435_, _42433_);
  or _49475_ (_01269_, _42436_, _42432_);
  nor _49476_ (_42437_, _42260_, _42214_);
  and _49477_ (_42438_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _49478_ (_42439_, _42438_, _42437_);
  and _49479_ (_42440_, _42439_, _42239_);
  nand _49480_ (_42441_, _42108_, _39291_);
  nand _49481_ (_42442_, _42109_, _39298_);
  and _49482_ (_42443_, _42442_, _42206_);
  and _49483_ (_42444_, _42443_, _42441_);
  or _49484_ (_01271_, _42444_, _42440_);
  nor _49485_ (_42445_, _42260_, _42210_);
  and _49486_ (_42446_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _49487_ (_42447_, _42446_, _42445_);
  and _49488_ (_42448_, _42447_, _42239_);
  nand _49489_ (_42449_, _42109_, _39291_);
  nand _49490_ (_42450_, _42108_, _39284_);
  and _49491_ (_42451_, _42450_, _42206_);
  and _49492_ (_42452_, _42451_, _42449_);
  or _49493_ (_01273_, _42452_, _42448_);
  and _49494_ (_42453_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _49495_ (_42454_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _49496_ (_42455_, _42454_, _42453_);
  and _49497_ (_42456_, _42455_, _42239_);
  nand _49498_ (_42457_, _42108_, _39276_);
  nand _49499_ (_42458_, _42109_, _39284_);
  and _49500_ (_42459_, _42458_, _42206_);
  and _49501_ (_42460_, _42459_, _42457_);
  or _49502_ (_01275_, _42460_, _42456_);
  and _49503_ (_42461_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _49504_ (_42462_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _49505_ (_42463_, _42462_, _42461_);
  and _49506_ (_42464_, _42463_, _42239_);
  nand _49507_ (_42465_, _42109_, _39276_);
  nand _49508_ (_42466_, _42108_, _39268_);
  and _49509_ (_42467_, _42466_, _42206_);
  and _49510_ (_42468_, _42467_, _42465_);
  or _49511_ (_01276_, _42468_, _42464_);
  and _49512_ (_42469_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _49513_ (_42470_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _49514_ (_42471_, _42470_, _42469_);
  and _49515_ (_42472_, _42471_, _42239_);
  nand _49516_ (_42473_, _42108_, _39261_);
  nand _49517_ (_42474_, _42109_, _39268_);
  and _49518_ (_42475_, _42474_, _42206_);
  and _49519_ (_42476_, _42475_, _42473_);
  or _49520_ (_01278_, _42476_, _42472_);
  and _49521_ (_42477_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _49522_ (_42478_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _49523_ (_42479_, _42478_, _42477_);
  and _49524_ (_42480_, _42479_, _42239_);
  nand _49525_ (_42481_, _42108_, _39327_);
  nand _49526_ (_42482_, _42109_, _39261_);
  and _49527_ (_42483_, _42482_, _42206_);
  and _49528_ (_42484_, _42483_, _42481_);
  or _49529_ (_01280_, _42484_, _42480_);
  and _49530_ (_42485_, _42205_, _42109_);
  nand _49531_ (_42486_, _42485_, _39327_);
  or _49532_ (_42487_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _49533_ (_42488_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _49534_ (_42489_, _42488_, _42487_);
  or _49535_ (_42490_, _42489_, _42205_);
  and _49536_ (_42491_, _42490_, _43634_);
  and _49537_ (_01282_, _42491_, _42486_);
  and _49538_ (_42492_, _42428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _49539_ (_42493_, _42260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _49540_ (_42494_, _42493_, _42492_);
  and _49541_ (_42495_, _42494_, _42239_);
  or _49542_ (_42496_, _42096_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _49543_ (_42497_, _42496_, _42109_);
  and _49544_ (_42498_, _42497_, _42206_);
  or _49545_ (_01284_, _42498_, _42495_);
  nand _49546_ (_42499_, _42264_, _39306_);
  or _49547_ (_42500_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _49548_ (_42501_, _42500_, _43634_);
  and _49549_ (_01286_, _42501_, _42499_);
  or _49550_ (_42502_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _49551_ (_42503_, _42502_, _43634_);
  nand _49552_ (_42504_, _42264_, _39298_);
  and _49553_ (_01288_, _42504_, _42503_);
  or _49554_ (_42505_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _49555_ (_42506_, _42505_, _43634_);
  nand _49556_ (_42507_, _42264_, _39291_);
  and _49557_ (_01290_, _42507_, _42506_);
  or _49558_ (_42508_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _49559_ (_42509_, _42508_, _43634_);
  nand _49560_ (_42510_, _42264_, _39284_);
  and _49561_ (_01292_, _42510_, _42509_);
  or _49562_ (_42511_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _49563_ (_42512_, _42511_, _43634_);
  nand _49564_ (_42513_, _42264_, _39276_);
  and _49565_ (_01294_, _42513_, _42512_);
  or _49566_ (_42514_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _49567_ (_42515_, _42514_, _43634_);
  nand _49568_ (_42516_, _42264_, _39268_);
  and _49569_ (_01296_, _42516_, _42515_);
  or _49570_ (_42517_, _42264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _49571_ (_42518_, _42517_, _43634_);
  nand _49572_ (_42519_, _42264_, _39261_);
  and _49573_ (_01298_, _42519_, _42518_);
  not _49574_ (_42520_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _49575_ (_42521_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _42520_);
  or _49576_ (_42522_, _42521_, _42108_);
  nor _49577_ (_42523_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _49578_ (_42524_, _42523_, _42522_);
  or _49579_ (_42525_, _42524_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _49580_ (_42526_, _42525_, _42268_);
  nand _49581_ (_42527_, _39957_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _49582_ (_42528_, _42527_, _42268_);
  or _49583_ (_42529_, _42528_, _39958_);
  and _49584_ (_42530_, _42529_, _42526_);
  or _49585_ (_42531_, _42530_, _42271_);
  nand _49586_ (_42532_, _42271_, _39306_);
  and _49587_ (_42533_, _42532_, _43634_);
  and _49588_ (_01299_, _42533_, _42531_);
  or _49589_ (_42534_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _49590_ (_42535_, _42534_, _42268_);
  nand _49591_ (_42536_, _39974_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _49592_ (_42537_, _42536_, _42268_);
  or _49593_ (_42538_, _42537_, _39975_);
  and _49594_ (_42539_, _42538_, _42535_);
  or _49595_ (_42540_, _42539_, _42271_);
  nand _49596_ (_42541_, _42271_, _39298_);
  and _49597_ (_42542_, _42541_, _43634_);
  and _49598_ (_01300_, _42542_, _42540_);
  not _49599_ (_42543_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _49600_ (_42544_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _49601_ (_42545_, _42121_, _42544_);
  nor _49602_ (_42546_, _42545_, _42543_);
  and _49603_ (_42547_, _42545_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _49604_ (_42548_, _42547_, _42546_);
  or _49605_ (_42549_, _42548_, _42268_);
  or _49606_ (_42550_, _34509_, _42543_);
  nand _49607_ (_42551_, _42550_, _42268_);
  or _49608_ (_42552_, _42551_, _34531_);
  and _49609_ (_42553_, _42552_, _42549_);
  or _49610_ (_42554_, _42553_, _42271_);
  nand _49611_ (_42555_, _42271_, _39291_);
  and _49612_ (_42556_, _42555_, _43634_);
  and _49613_ (_01301_, _42556_, _42554_);
  and _49614_ (_42557_, _42268_, _35217_);
  nand _49615_ (_42558_, _42557_, _32431_);
  or _49616_ (_42559_, _42557_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _49617_ (_42560_, _42559_, _42272_);
  and _49618_ (_42561_, _42560_, _42558_);
  nor _49619_ (_42562_, _42272_, _39284_);
  or _49620_ (_42563_, _42562_, _42561_);
  and _49621_ (_01303_, _42563_, _43634_);
  and _49622_ (_42564_, _42268_, _35978_);
  nand _49623_ (_42565_, _42564_, _32431_);
  or _49624_ (_42566_, _42564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _49625_ (_42567_, _42566_, _42272_);
  and _49626_ (_42568_, _42567_, _42565_);
  nor _49627_ (_42569_, _42272_, _39276_);
  or _49628_ (_42570_, _42569_, _42568_);
  and _49629_ (_01305_, _42570_, _43634_);
  and _49630_ (_42571_, _42268_, _36762_);
  nand _49631_ (_42572_, _42571_, _32431_);
  or _49632_ (_42573_, _42571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _49633_ (_42574_, _42573_, _42272_);
  and _49634_ (_42575_, _42574_, _42572_);
  nor _49635_ (_42576_, _42272_, _39268_);
  or _49636_ (_42577_, _42576_, _42575_);
  and _49637_ (_01307_, _42577_, _43634_);
  and _49638_ (_42578_, _42268_, _37502_);
  nand _49639_ (_42579_, _42578_, _32431_);
  or _49640_ (_42580_, _42578_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _49641_ (_42581_, _42580_, _42272_);
  and _49642_ (_42582_, _42581_, _42579_);
  nor _49643_ (_42583_, _42272_, _39261_);
  or _49644_ (_42584_, _42583_, _42582_);
  and _49645_ (_01309_, _42584_, _43634_);
  and _49646_ (_01615_, t2_i, _43634_);
  nor _49647_ (_42585_, t2_i, rst);
  and _49648_ (_01618_, _42585_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _49649_ (_42586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _43634_);
  nor _49650_ (_01621_, _42586_, t2ex_i);
  and _49651_ (_01624_, t2ex_i, _43634_);
  and _49652_ (_42587_, _39240_, _39760_);
  and _49653_ (_42588_, _42587_, _40845_);
  nand _49654_ (_42589_, _42588_, _39327_);
  and _49655_ (_42590_, _42587_, _40697_);
  not _49656_ (_42591_, _42590_);
  and _49657_ (_42592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _49658_ (_42593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _49659_ (_42594_, _42593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49660_ (_42595_, _42594_, _42592_);
  not _49661_ (_42596_, _42595_);
  and _49662_ (_42597_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _49663_ (_42598_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _49664_ (_42599_, _42598_, _42597_);
  or _49665_ (_42600_, _42588_, _42599_);
  and _49666_ (_42601_, _42600_, _42591_);
  and _49667_ (_42602_, _42601_, _42589_);
  and _49668_ (_42603_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _49669_ (_42604_, _42603_, _42602_);
  and _49670_ (_01627_, _42604_, _43634_);
  nand _49671_ (_42605_, _42590_, _39327_);
  nor _49672_ (_42606_, _42588_, _42596_);
  or _49673_ (_42607_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _49674_ (_42608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _49675_ (_42609_, _42606_, _42608_);
  and _49676_ (_42610_, _42609_, _42607_);
  or _49677_ (_42611_, _42610_, _42590_);
  and _49678_ (_42612_, _42611_, _43634_);
  and _49679_ (_01630_, _42612_, _42605_);
  and _49680_ (_42613_, _42587_, _36762_);
  and _49681_ (_42614_, _42613_, _40696_);
  and _49682_ (_42615_, _42587_, _40805_);
  nor _49683_ (_42616_, _42615_, _42614_);
  not _49684_ (_42617_, _42593_);
  or _49685_ (_42618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _49686_ (_42619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _49687_ (_42620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _42619_);
  and _49688_ (_42621_, _42620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _49689_ (_42622_, _42621_, _42618_);
  and _49690_ (_42623_, _42622_, _42617_);
  and _49691_ (_42624_, _42623_, _42616_);
  or _49692_ (_42625_, _42624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _49693_ (_42626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49694_ (_42627_, _42626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49695_ (_42628_, _42627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49696_ (_42629_, _42628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49697_ (_42630_, _42629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49698_ (_42631_, _42630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _49699_ (_42632_, _42631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _49700_ (_42633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _49701_ (_42634_, _42633_, _42632_);
  and _49702_ (_42635_, _42634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _49703_ (_42636_, _42635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _49704_ (_42637_, _42636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _49705_ (_42638_, _42637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _49706_ (_42639_, _42638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _49707_ (_42640_, _42639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _49708_ (_42641_, _42640_);
  nand _49709_ (_42642_, _42641_, _42624_);
  and _49710_ (_42643_, _42642_, _43634_);
  and _49711_ (_01633_, _42643_, _42625_);
  nand _49712_ (_42644_, _42615_, _39327_);
  not _49713_ (_42645_, _42614_);
  not _49714_ (_42646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49715_ (_42647_, _42592_, _42646_);
  and _49716_ (_42648_, _42647_, _42593_);
  and _49717_ (_42649_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _49718_ (_42650_, _42648_);
  not _49719_ (_42651_, _42594_);
  and _49720_ (_42652_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _49721_ (_42653_, _42640_, _42622_);
  and _49722_ (_42654_, _42653_, _42652_);
  and _49723_ (_42655_, _42631_, _42622_);
  nor _49724_ (_42656_, _42655_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _49725_ (_42657_, _42632_, _42622_);
  nor _49726_ (_42658_, _42657_, _42656_);
  or _49727_ (_42659_, _42658_, _42654_);
  and _49728_ (_42660_, _42659_, _42650_);
  or _49729_ (_42661_, _42660_, _42649_);
  or _49730_ (_42662_, _42661_, _42615_);
  and _49731_ (_42663_, _42662_, _42645_);
  and _49732_ (_42664_, _42663_, _42644_);
  and _49733_ (_42665_, _42614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _49734_ (_42666_, _42665_, _42664_);
  and _49735_ (_01636_, _42666_, _43634_);
  nand _49736_ (_42667_, _42614_, _39327_);
  nor _49737_ (_42668_, _42648_, _42608_);
  and _49738_ (_42669_, _42650_, _42622_);
  and _49739_ (_42670_, _42669_, _42639_);
  or _49740_ (_42671_, _42670_, _42668_);
  nand _49741_ (_42672_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _49742_ (_42673_, _42672_, _42653_);
  and _49743_ (_42674_, _42673_, _42671_);
  nand _49744_ (_42675_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _49745_ (_42676_, _42675_, _42616_);
  or _49746_ (_42677_, _42676_, _42674_);
  nand _49747_ (_42678_, _42615_, _42608_);
  and _49748_ (_42679_, _42678_, _43634_);
  and _49749_ (_42680_, _42679_, _42677_);
  and _49750_ (_01639_, _42680_, _42667_);
  and _49751_ (_42681_, _42593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _49752_ (_42682_, _42681_, _42670_);
  nand _49753_ (_42683_, _42682_, _42616_);
  or _49754_ (_42684_, _42616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49755_ (_42685_, _42684_, _43634_);
  and _49756_ (_01642_, _42685_, _42683_);
  or _49757_ (_42686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49758_ (_42687_, _41408_, _39742_);
  or _49759_ (_42688_, _42687_, _42686_);
  nand _49760_ (_42689_, _39745_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _49761_ (_42690_, _42689_, _42687_);
  or _49762_ (_42691_, _42690_, _39746_);
  and _49763_ (_42692_, _42691_, _42688_);
  and _49764_ (_42693_, _42587_, _41404_);
  or _49765_ (_42694_, _42693_, _42692_);
  nand _49766_ (_42695_, _42693_, _39327_);
  and _49767_ (_42696_, _42695_, _43634_);
  and _49768_ (_01645_, _42696_, _42694_);
  or _49769_ (_42697_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _49770_ (_42698_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49771_ (_42699_, _42698_, _42697_);
  or _49772_ (_42700_, _42699_, _42588_);
  nand _49773_ (_42701_, _42588_, _39306_);
  and _49774_ (_42702_, _42701_, _42700_);
  or _49775_ (_42703_, _42702_, _42590_);
  or _49776_ (_42704_, _42591_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _49777_ (_42705_, _42704_, _43634_);
  and _49778_ (_02131_, _42705_, _42703_);
  nand _49779_ (_42706_, _42588_, _39298_);
  and _49780_ (_42707_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49781_ (_42708_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _49782_ (_42709_, _42708_, _42707_);
  or _49783_ (_42710_, _42709_, _42588_);
  and _49784_ (_42711_, _42710_, _42591_);
  and _49785_ (_42712_, _42711_, _42706_);
  and _49786_ (_42713_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _49787_ (_42714_, _42713_, _42712_);
  and _49788_ (_02133_, _42714_, _43634_);
  nand _49789_ (_42715_, _42588_, _39291_);
  and _49790_ (_42716_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49791_ (_42717_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49792_ (_42718_, _42717_, _42716_);
  or _49793_ (_42719_, _42718_, _42588_);
  and _49794_ (_42720_, _42719_, _42591_);
  and _49795_ (_42721_, _42720_, _42715_);
  and _49796_ (_42722_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _49797_ (_42723_, _42722_, _42721_);
  and _49798_ (_02135_, _42723_, _43634_);
  nand _49799_ (_42724_, _42588_, _39284_);
  and _49800_ (_42725_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49801_ (_42726_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49802_ (_42727_, _42726_, _42725_);
  or _49803_ (_42728_, _42727_, _42588_);
  and _49804_ (_42729_, _42728_, _42591_);
  and _49805_ (_42730_, _42729_, _42724_);
  and _49806_ (_42731_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _49807_ (_42732_, _42731_, _42730_);
  and _49808_ (_02136_, _42732_, _43634_);
  nand _49809_ (_42733_, _42588_, _39276_);
  and _49810_ (_42734_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49811_ (_42735_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49812_ (_42736_, _42735_, _42734_);
  or _49813_ (_42737_, _42736_, _42588_);
  and _49814_ (_42738_, _42737_, _42591_);
  and _49815_ (_42739_, _42738_, _42733_);
  and _49816_ (_42740_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _49817_ (_42741_, _42740_, _42739_);
  and _49818_ (_02138_, _42741_, _43634_);
  nand _49819_ (_42742_, _42588_, _39268_);
  and _49820_ (_42743_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49821_ (_42744_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49822_ (_42745_, _42744_, _42743_);
  or _49823_ (_42746_, _42745_, _42588_);
  and _49824_ (_42747_, _42746_, _42591_);
  and _49825_ (_42748_, _42747_, _42742_);
  and _49826_ (_42749_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _49827_ (_42750_, _42749_, _42748_);
  and _49828_ (_02140_, _42750_, _43634_);
  nand _49829_ (_42751_, _42588_, _39261_);
  and _49830_ (_42752_, _42596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49831_ (_42753_, _42595_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _49832_ (_42754_, _42753_, _42752_);
  or _49833_ (_42755_, _42754_, _42588_);
  and _49834_ (_42756_, _42755_, _42591_);
  and _49835_ (_42757_, _42756_, _42751_);
  and _49836_ (_42758_, _42590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _49837_ (_42759_, _42758_, _42757_);
  and _49838_ (_02142_, _42759_, _43634_);
  or _49839_ (_42760_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _49840_ (_42761_, _42606_);
  or _49841_ (_42762_, _42761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _49842_ (_42763_, _42762_, _42760_);
  or _49843_ (_42764_, _42763_, _42590_);
  nand _49844_ (_42765_, _42590_, _39306_);
  and _49845_ (_42766_, _42765_, _43634_);
  and _49846_ (_02143_, _42766_, _42764_);
  or _49847_ (_42767_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not _49848_ (_42768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _49849_ (_42769_, _42606_, _42768_);
  and _49850_ (_42770_, _42769_, _42767_);
  or _49851_ (_42771_, _42770_, _42590_);
  nand _49852_ (_42772_, _42590_, _39298_);
  and _49853_ (_42773_, _42772_, _43634_);
  and _49854_ (_02145_, _42773_, _42771_);
  nand _49855_ (_42774_, _42590_, _39291_);
  and _49856_ (_42775_, _42761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49857_ (_42776_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49858_ (_42777_, _42776_, _42775_);
  or _49859_ (_42778_, _42777_, _42590_);
  and _49860_ (_42779_, _42778_, _43634_);
  and _49861_ (_02147_, _42779_, _42774_);
  nand _49862_ (_42780_, _42590_, _39284_);
  and _49863_ (_42781_, _42761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49864_ (_42782_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49865_ (_42783_, _42782_, _42781_);
  or _49866_ (_42784_, _42783_, _42590_);
  and _49867_ (_42785_, _42784_, _43634_);
  and _49868_ (_02149_, _42785_, _42780_);
  nand _49869_ (_42786_, _42590_, _39276_);
  or _49870_ (_42787_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  not _49871_ (_42788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand _49872_ (_42789_, _42606_, _42788_);
  and _49873_ (_42790_, _42789_, _42787_);
  or _49874_ (_42791_, _42790_, _42590_);
  and _49875_ (_42792_, _42791_, _43634_);
  and _49876_ (_02150_, _42792_, _42786_);
  nand _49877_ (_42793_, _42590_, _39268_);
  or _49878_ (_42794_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  not _49879_ (_42795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _49880_ (_42796_, _42606_, _42795_);
  and _49881_ (_42797_, _42796_, _42794_);
  or _49882_ (_42798_, _42797_, _42590_);
  and _49883_ (_42799_, _42798_, _43634_);
  and _49884_ (_02152_, _42799_, _42793_);
  nand _49885_ (_42800_, _42590_, _39261_);
  or _49886_ (_42801_, _42606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  not _49887_ (_42802_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _49888_ (_42803_, _42606_, _42802_);
  and _49889_ (_42804_, _42803_, _42801_);
  or _49890_ (_42805_, _42804_, _42590_);
  and _49891_ (_42806_, _42805_, _43634_);
  and _49892_ (_02154_, _42806_, _42800_);
  and _49893_ (_42807_, _42622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49894_ (_42808_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _49895_ (_42809_, _42808_, _42640_);
  nand _49896_ (_42810_, _42809_, _42807_);
  or _49897_ (_42811_, _42622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49898_ (_42812_, _42811_, _42650_);
  and _49899_ (_42813_, _42812_, _42810_);
  and _49900_ (_42814_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _49901_ (_42815_, _42814_, _42615_);
  or _49902_ (_42816_, _42815_, _42813_);
  and _49903_ (_42817_, _42615_, _39306_);
  nor _49904_ (_42818_, _42817_, _42614_);
  and _49905_ (_42819_, _42818_, _42816_);
  and _49906_ (_42820_, _42614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _49907_ (_42821_, _42820_, _42819_);
  and _49908_ (_02156_, _42821_, _43634_);
  and _49909_ (_42822_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49910_ (_42823_, _42822_, _42669_);
  and _49911_ (_42824_, _42823_, _42640_);
  and _49912_ (_42825_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not _49913_ (_42826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _49914_ (_42827_, _42807_, _42826_);
  and _49915_ (_42828_, _42807_, _42826_);
  or _49916_ (_42829_, _42828_, _42827_);
  and _49917_ (_42830_, _42829_, _42650_);
  nor _49918_ (_42831_, _42830_, _42825_);
  nand _49919_ (_42832_, _42831_, _42616_);
  or _49920_ (_42833_, _42832_, _42824_);
  nand _49921_ (_42834_, _42615_, _39298_);
  nand _49922_ (_42835_, _42614_, _42826_);
  and _49923_ (_42836_, _42835_, _43634_);
  and _49924_ (_42837_, _42836_, _42834_);
  and _49925_ (_02157_, _42837_, _42833_);
  and _49926_ (_42838_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49927_ (_42839_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49928_ (_42840_, _42839_, _42653_);
  nand _49929_ (_42841_, _42626_, _42622_);
  nor _49930_ (_42842_, _42841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49931_ (_42843_, _42841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49932_ (_42844_, _42843_, _42842_);
  or _49933_ (_42845_, _42844_, _42840_);
  and _49934_ (_42846_, _42845_, _42650_);
  or _49935_ (_42847_, _42846_, _42838_);
  or _49936_ (_42848_, _42847_, _42615_);
  nand _49937_ (_42849_, _42615_, _39291_);
  and _49938_ (_42850_, _42849_, _42645_);
  and _49939_ (_42851_, _42850_, _42848_);
  and _49940_ (_42852_, _42614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49941_ (_42853_, _42852_, _42851_);
  and _49942_ (_02159_, _42853_, _43634_);
  and _49943_ (_42854_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49944_ (_42855_, _42854_, _42653_);
  nand _49945_ (_42856_, _42627_, _42622_);
  nor _49946_ (_42857_, _42856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49947_ (_42858_, _42856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49948_ (_42859_, _42858_, _42857_);
  or _49949_ (_42860_, _42859_, _42855_);
  and _49950_ (_42861_, _42860_, _42650_);
  nand _49951_ (_42862_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand _49952_ (_42863_, _42862_, _42616_);
  or _49953_ (_42864_, _42863_, _42861_);
  nand _49954_ (_42865_, _42615_, _39284_);
  or _49955_ (_42866_, _42645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49956_ (_42867_, _42866_, _43634_);
  and _49957_ (_42868_, _42867_, _42865_);
  and _49958_ (_02161_, _42868_, _42864_);
  nand _49959_ (_42869_, _42615_, _39276_);
  or _49960_ (_42870_, _42645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49961_ (_42871_, _42870_, _43634_);
  and _49962_ (_42872_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49963_ (_42873_, _42872_, _42653_);
  nand _49964_ (_42874_, _42628_, _42622_);
  nor _49965_ (_42875_, _42874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49966_ (_42876_, _42874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49967_ (_42877_, _42876_, _42875_);
  or _49968_ (_42878_, _42877_, _42873_);
  and _49969_ (_42879_, _42878_, _42650_);
  nand _49970_ (_42880_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _49971_ (_42881_, _42880_, _42616_);
  or _49972_ (_42882_, _42881_, _42879_);
  and _49973_ (_42883_, _42882_, _42871_);
  and _49974_ (_02163_, _42883_, _42869_);
  and _49975_ (_42884_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49976_ (_42885_, _42884_, _42653_);
  nand _49977_ (_42886_, _42629_, _42622_);
  nor _49978_ (_42887_, _42886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49979_ (_42888_, _42886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49980_ (_42889_, _42888_, _42887_);
  or _49981_ (_42890_, _42889_, _42885_);
  and _49982_ (_42891_, _42890_, _42650_);
  nand _49983_ (_42892_, _42648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand _49984_ (_42893_, _42892_, _42616_);
  or _49985_ (_42894_, _42893_, _42891_);
  nand _49986_ (_42895_, _42615_, _39268_);
  or _49987_ (_42896_, _42645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49988_ (_42897_, _42896_, _43634_);
  and _49989_ (_42898_, _42897_, _42895_);
  and _49990_ (_02164_, _42898_, _42894_);
  not _49991_ (_42899_, _39261_);
  and _49992_ (_42900_, _42615_, _42899_);
  and _49993_ (_42901_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49994_ (_42902_, _42901_, _42653_);
  and _49995_ (_42903_, _42630_, _42622_);
  nor _49996_ (_42904_, _42903_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _49997_ (_42905_, _42904_, _42655_);
  or _49998_ (_42906_, _42905_, _42648_);
  or _49999_ (_42907_, _42906_, _42902_);
  or _50000_ (_42908_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _50001_ (_42909_, _42908_, _42616_);
  and _50002_ (_42910_, _42909_, _42907_);
  and _50003_ (_42911_, _42614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _50004_ (_42912_, _42911_, _42910_);
  or _50005_ (_42913_, _42912_, _42900_);
  and _50006_ (_02166_, _42913_, _43634_);
  and _50007_ (_42914_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _50008_ (_42915_, _42914_, _42653_);
  or _50009_ (_42916_, _42657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _50010_ (_42917_, _42657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _50011_ (_42918_, _42917_, _42916_);
  or _50012_ (_42919_, _42918_, _42648_);
  or _50013_ (_42920_, _42919_, _42915_);
  or _50014_ (_42921_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _50015_ (_42922_, _42921_, _42616_);
  and _50016_ (_42923_, _42922_, _42920_);
  and _50017_ (_42924_, _42615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _50018_ (_42925_, _42614_, _39307_);
  or _50019_ (_42926_, _42925_, _42924_);
  or _50020_ (_42927_, _42926_, _42923_);
  and _50021_ (_02168_, _42927_, _43634_);
  and _50022_ (_42928_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _50023_ (_42929_, _42928_, _42653_);
  nand _50024_ (_42930_, _42917_, _42768_);
  nand _50025_ (_42931_, _42634_, _42622_);
  and _50026_ (_42932_, _42931_, _42930_);
  or _50027_ (_42933_, _42932_, _42648_);
  or _50028_ (_42934_, _42933_, _42929_);
  not _50029_ (_42935_, _42616_);
  nor _50030_ (_42936_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _50031_ (_42937_, _42936_, _42935_);
  and _50032_ (_42938_, _42937_, _42934_);
  and _50033_ (_42939_, _42615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _50034_ (_42940_, _42645_, _39298_);
  or _50035_ (_42941_, _42940_, _42939_);
  or _50036_ (_42942_, _42941_, _42938_);
  and _50037_ (_02170_, _42942_, _43634_);
  and _50038_ (_42943_, _40705_, _33748_);
  and _50039_ (_42944_, _42587_, _42943_);
  and _50040_ (_42945_, _42944_, _31886_);
  not _50041_ (_42946_, _42945_);
  and _50042_ (_42947_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _50043_ (_42948_, _42947_, _42653_);
  and _50044_ (_42949_, _42931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _50045_ (_42950_, _42931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _50046_ (_42951_, _42950_, _42648_);
  or _50047_ (_42952_, _42951_, _42949_);
  or _50048_ (_42953_, _42952_, _42948_);
  nor _50049_ (_42954_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _50050_ (_42955_, _42954_, _42615_);
  and _50051_ (_42956_, _42955_, _42953_);
  and _50052_ (_42957_, _40705_, _28260_);
  and _50053_ (_42958_, _42587_, _42957_);
  and _50054_ (_42959_, _42958_, _31886_);
  and _50055_ (_42960_, _42959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _50056_ (_42961_, _42960_, _42956_);
  and _50057_ (_42962_, _42961_, _42946_);
  nor _50058_ (_42963_, _42946_, _39291_);
  or _50059_ (_42964_, _42963_, _42962_);
  and _50060_ (_02171_, _42964_, _43634_);
  and _50061_ (_42965_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _50062_ (_42966_, _42965_, _42653_);
  nand _50063_ (_42967_, _42635_, _42622_);
  nor _50064_ (_42968_, _42967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _50065_ (_42969_, _42967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _50066_ (_42970_, _42969_, _42648_);
  or _50067_ (_42971_, _42970_, _42968_);
  or _50068_ (_42972_, _42971_, _42966_);
  or _50069_ (_42973_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _50070_ (_42974_, _42973_, _42616_);
  and _50071_ (_42975_, _42974_, _42972_);
  and _50072_ (_42976_, _42615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _50073_ (_42977_, _42976_, _42975_);
  nor _50074_ (_42978_, _42645_, _39284_);
  or _50075_ (_42979_, _42978_, _42977_);
  and _50076_ (_02173_, _42979_, _43634_);
  and _50077_ (_42980_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _50078_ (_42981_, _42980_, _42653_);
  and _50079_ (_42982_, _42636_, _42622_);
  and _50080_ (_42983_, _42982_, _42788_);
  nor _50081_ (_42984_, _42982_, _42788_);
  or _50082_ (_42985_, _42984_, _42648_);
  or _50083_ (_42986_, _42985_, _42983_);
  or _50084_ (_42987_, _42986_, _42981_);
  or _50085_ (_42988_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _50086_ (_42989_, _42988_, _42616_);
  and _50087_ (_42990_, _42989_, _42987_);
  and _50088_ (_42991_, _42615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _50089_ (_42992_, _42991_, _42990_);
  nor _50090_ (_42993_, _42645_, _39276_);
  or _50091_ (_42994_, _42993_, _42992_);
  and _50092_ (_02175_, _42994_, _43634_);
  and _50093_ (_42995_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _50094_ (_42996_, _42995_, _42653_);
  and _50095_ (_42997_, _42637_, _42622_);
  nor _50096_ (_42998_, _42997_, _42795_);
  and _50097_ (_42999_, _42997_, _42795_);
  or _50098_ (_43000_, _42999_, _42648_);
  or _50099_ (_43001_, _43000_, _42998_);
  or _50100_ (_43002_, _43001_, _42996_);
  nor _50101_ (_43003_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _50102_ (_43004_, _43003_, _42615_);
  and _50103_ (_43005_, _43004_, _43002_);
  and _50104_ (_43006_, _42959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _50105_ (_43007_, _43006_, _43005_);
  and _50106_ (_43008_, _43007_, _42946_);
  nor _50107_ (_43009_, _42946_, _39268_);
  or _50108_ (_43010_, _43009_, _43008_);
  and _50109_ (_02177_, _43010_, _43634_);
  and _50110_ (_43011_, _42615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _50111_ (_43012_, _42651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _50112_ (_43013_, _43012_, _42653_);
  and _50113_ (_43014_, _42638_, _42622_);
  nor _50114_ (_43015_, _43014_, _42802_);
  and _50115_ (_43016_, _43014_, _42802_);
  or _50116_ (_43017_, _43016_, _42648_);
  or _50117_ (_43018_, _43017_, _43015_);
  or _50118_ (_43019_, _43018_, _43013_);
  or _50119_ (_43020_, _42650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _50120_ (_43021_, _43020_, _42616_);
  and _50121_ (_43022_, _43021_, _43019_);
  or _50122_ (_43023_, _43022_, _43011_);
  nor _50123_ (_43024_, _42645_, _39261_);
  or _50124_ (_43025_, _43024_, _43023_);
  and _50125_ (_02178_, _43025_, _43634_);
  not _50126_ (_43026_, _42693_);
  and _50127_ (_43027_, _42687_, _28271_);
  or _50128_ (_43028_, _43027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _50129_ (_43029_, _43028_, _43026_);
  nand _50130_ (_43030_, _43027_, _32431_);
  and _50131_ (_43031_, _43030_, _43029_);
  and _50132_ (_43032_, _42693_, _39307_);
  or _50133_ (_43033_, _43032_, _43031_);
  and _50134_ (_02180_, _43033_, _43634_);
  and _50135_ (_43034_, _42687_, _39768_);
  or _50136_ (_43035_, _43034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _50137_ (_43036_, _43035_, _43026_);
  nand _50138_ (_43037_, _43034_, _32431_);
  and _50139_ (_43038_, _43037_, _43036_);
  nor _50140_ (_43039_, _43026_, _39298_);
  or _50141_ (_43040_, _43039_, _43038_);
  and _50142_ (_02182_, _43040_, _43634_);
  nand _50143_ (_43041_, _42687_, _40329_);
  and _50144_ (_43042_, _43041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _50145_ (_43043_, _43042_, _42693_);
  and _50146_ (_43044_, _34542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _50147_ (_43045_, _43044_, _34531_);
  and _50148_ (_43046_, _43045_, _42687_);
  or _50149_ (_43047_, _43046_, _43043_);
  nand _50150_ (_43048_, _42693_, _39291_);
  and _50151_ (_43049_, _43048_, _43634_);
  and _50152_ (_02184_, _43049_, _43047_);
  and _50153_ (_43050_, _42687_, _35217_);
  or _50154_ (_43051_, _43050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _50155_ (_43052_, _43051_, _43026_);
  nand _50156_ (_43053_, _43050_, _32431_);
  and _50157_ (_43054_, _43053_, _43052_);
  nor _50158_ (_43055_, _43026_, _39284_);
  or _50159_ (_43056_, _43055_, _43054_);
  and _50160_ (_02185_, _43056_, _43634_);
  and _50161_ (_43057_, _42687_, _35978_);
  or _50162_ (_43058_, _43057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _50163_ (_43059_, _43058_, _43026_);
  nand _50164_ (_43060_, _43057_, _32431_);
  and _50165_ (_43061_, _43060_, _43059_);
  nor _50166_ (_43062_, _43026_, _39276_);
  or _50167_ (_43063_, _43062_, _43061_);
  and _50168_ (_02186_, _43063_, _43634_);
  and _50169_ (_43064_, _42687_, _36762_);
  or _50170_ (_43065_, _43064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _50171_ (_43066_, _43065_, _43026_);
  nand _50172_ (_43067_, _43064_, _32431_);
  and _50173_ (_43068_, _43067_, _43066_);
  nor _50174_ (_43069_, _43026_, _39268_);
  or _50175_ (_43070_, _43069_, _43068_);
  and _50176_ (_02187_, _43070_, _43634_);
  not _50177_ (_43071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _50178_ (_43072_, _42592_, _43071_);
  or _50179_ (_43073_, _43072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _50180_ (_43074_, _43073_, _42687_);
  nand _50181_ (_43075_, _39910_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _50182_ (_43076_, _43075_, _42687_);
  or _50183_ (_43077_, _43076_, _39911_);
  and _50184_ (_43078_, _43077_, _43074_);
  or _50185_ (_43079_, _43078_, _42693_);
  nand _50186_ (_43080_, _42693_, _39261_);
  and _50187_ (_43081_, _43080_, _43634_);
  and _50188_ (_02188_, _43081_, _43079_);
  nor _50189_ (_43082_, _39148_, _39135_);
  nor _50190_ (_43083_, _39128_, _39120_);
  and _50191_ (_43084_, _43083_, _39172_);
  and _50192_ (_43085_, _43084_, _43082_);
  not _50193_ (_43086_, _39140_);
  and _50194_ (_43087_, _43086_, _39127_);
  and _50195_ (_43088_, _43087_, _39182_);
  and _50196_ (_43089_, _43088_, _43085_);
  nor _50197_ (_43090_, _43089_, _37633_);
  or _50198_ (_43091_, _39175_, _39133_);
  and _50199_ (_43092_, _39092_, _43091_);
  or _50200_ (_43093_, _43092_, _43090_);
  not _50201_ (_43094_, _39237_);
  and _50202_ (_43095_, _43094_, _39205_);
  and _50203_ (_43096_, _43095_, _39105_);
  and _50204_ (_43097_, _38124_, _28250_);
  nor _50205_ (_43098_, _38124_, _28250_);
  not _50206_ (_43099_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _50207_ (_43100_, _31853_, _43099_);
  and _50208_ (_43101_, _43100_, _34542_);
  nand _50209_ (_43102_, _43101_, _28765_);
  or _50210_ (_43103_, _43102_, _43098_);
  nor _50211_ (_43104_, _43103_, _43097_);
  and _50212_ (_43105_, _39759_, _39760_);
  and _50213_ (_43106_, _43105_, _39761_);
  not _50214_ (_43107_, _43106_);
  and _50215_ (_43108_, _43107_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _50216_ (_43109_, _43108_, _39851_);
  and _50217_ (_43110_, _43109_, _28929_);
  nor _50218_ (_43111_, _43109_, _28929_);
  nor _50219_ (_43112_, _43111_, _43110_);
  and _50220_ (_43113_, _43112_, _43104_);
  and _50221_ (_43114_, _43109_, _38124_);
  and _50222_ (_43115_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _50223_ (_43116_, _43109_, _38124_);
  and _50224_ (_43117_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _50225_ (_43118_, _43117_, _43115_);
  nor _50226_ (_43119_, _43109_, _39118_);
  and _50227_ (_43120_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _50228_ (_43121_, _43109_, _39118_);
  and _50229_ (_43122_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _50230_ (_43123_, _43122_, _43120_);
  and _50231_ (_43124_, _43123_, _43118_);
  nor _50232_ (_43125_, _43124_, _43113_);
  not _50233_ (_43126_, _39291_);
  and _50234_ (_43127_, _43113_, _43126_);
  nor _50235_ (_43128_, _43127_, _43125_);
  not _50236_ (_43129_, _43128_);
  and _50237_ (_43130_, _43129_, _43096_);
  not _50238_ (_43131_, _43130_);
  not _50239_ (_43132_, _39349_);
  and _50240_ (_43133_, _43132_, _39239_);
  not _50241_ (_43134_, _43133_);
  and _50242_ (_43135_, _39105_, _39237_);
  and _50243_ (_43136_, _43135_, _39205_);
  and _50244_ (_43137_, _43136_, _38832_);
  nor _50245_ (_43138_, _43094_, _39205_);
  and _50246_ (_43139_, _43138_, _39105_);
  not _50247_ (_43140_, _37676_);
  and _50248_ (_43141_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  nor _50249_ (_43142_, _37742_, _43140_);
  not _50250_ (_43143_, _43142_);
  and _50251_ (_43144_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _50252_ (_43145_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _50253_ (_43146_, _43145_, _43144_);
  and _50254_ (_43147_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _50255_ (_43148_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _50256_ (_43149_, _43148_, _43147_);
  and _50257_ (_43150_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _50258_ (_43151_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _50259_ (_43152_, _43151_, _43150_);
  and _50260_ (_43153_, _43152_, _43149_);
  and _50261_ (_43154_, _43153_, _43146_);
  nor _50262_ (_43155_, _43154_, _43143_);
  nor _50263_ (_43156_, _43155_, _43141_);
  not _50264_ (_43157_, _43156_);
  and _50265_ (_43158_, _43157_, _43139_);
  nor _50266_ (_43159_, _43158_, _43137_);
  and _50267_ (_43160_, _43159_, _43134_);
  and _50268_ (_43161_, _43160_, _43131_);
  nor _50269_ (_43162_, _43161_, _43093_);
  not _50270_ (_43163_, _39105_);
  and _50271_ (_43164_, _43163_, _39237_);
  and _50272_ (_43165_, _43164_, _39205_);
  not _50273_ (_43166_, _39367_);
  and _50274_ (_43167_, _43166_, _39239_);
  nor _50275_ (_43168_, _43167_, _43165_);
  and _50276_ (_43169_, _39238_, _43163_);
  not _50277_ (_43170_, _43169_);
  and _50278_ (_43171_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _50279_ (_43172_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _50280_ (_43173_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _50281_ (_43174_, _43173_, _43172_);
  and _50282_ (_43175_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _50283_ (_43176_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _50284_ (_43177_, _43176_, _43175_);
  and _50285_ (_43178_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _50286_ (_43179_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _50287_ (_43180_, _43179_, _43178_);
  and _50288_ (_43181_, _43180_, _43177_);
  and _50289_ (_43182_, _43181_, _43174_);
  nor _50290_ (_43183_, _43182_, _43143_);
  nor _50291_ (_43184_, _43183_, _43171_);
  not _50292_ (_43185_, _43184_);
  and _50293_ (_43186_, _43185_, _43139_);
  and _50294_ (_43187_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not _50295_ (_43188_, _43187_);
  and _50296_ (_43189_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _50297_ (_43190_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _50298_ (_43191_, _43190_, _43189_);
  and _50299_ (_43192_, _43191_, _43188_);
  and _50300_ (_43193_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _50301_ (_43194_, _43193_, _43113_);
  and _50302_ (_43195_, _43194_, _43192_);
  and _50303_ (_43196_, _43113_, _39268_);
  or _50304_ (_43197_, _43196_, _43195_);
  not _50305_ (_43198_, _43197_);
  and _50306_ (_43199_, _43198_, _43096_);
  nor _50307_ (_43200_, _43199_, _43186_);
  and _50308_ (_43201_, _43200_, _43170_);
  and _50309_ (_43202_, _43201_, _43168_);
  not _50310_ (_43203_, _43202_);
  nor _50311_ (_43204_, _39180_, _39176_);
  not _50312_ (_43205_, _39091_);
  nor _50313_ (_43206_, _43205_, _43204_);
  nor _50314_ (_43207_, _43206_, _43090_);
  not _50315_ (_43208_, _43207_);
  and _50316_ (_43209_, _39329_, _39239_);
  not _50317_ (_43210_, _43209_);
  and _50318_ (_43211_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _50319_ (_43212_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _50320_ (_43213_, _43212_, _43211_);
  and _50321_ (_43214_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _50322_ (_43215_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _50323_ (_43216_, _43215_, _43214_);
  and _50324_ (_43217_, _43216_, _43213_);
  nor _50325_ (_43218_, _43217_, _43113_);
  not _50326_ (_43219_, _39327_);
  and _50327_ (_43220_, _43113_, _43219_);
  nor _50328_ (_43221_, _43220_, _43218_);
  not _50329_ (_43222_, _43221_);
  and _50330_ (_43223_, _43222_, _43095_);
  not _50331_ (_43224_, _43223_);
  and _50332_ (_43225_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _50333_ (_43226_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _50334_ (_43227_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _50335_ (_43228_, _43227_, _43226_);
  and _50336_ (_43229_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _50337_ (_43230_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _50338_ (_43231_, _43230_, _43229_);
  and _50339_ (_43232_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _50340_ (_43233_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _50341_ (_43234_, _43233_, _43232_);
  and _50342_ (_43235_, _43234_, _43231_);
  and _50343_ (_43236_, _43235_, _43228_);
  nor _50344_ (_43237_, _43236_, _43143_);
  nor _50345_ (_43238_, _43237_, _43225_);
  not _50346_ (_43239_, _43238_);
  and _50347_ (_43240_, _43239_, _43138_);
  nor _50348_ (_43241_, _43240_, _43163_);
  and _50349_ (_43242_, _43241_, _43224_);
  and _50350_ (_43243_, _43242_, _43210_);
  and _50351_ (_43244_, _43243_, _43208_);
  and _50352_ (_43245_, _43244_, _43203_);
  nor _50353_ (_43246_, _43245_, _43162_);
  not _50354_ (_43247_, _43246_);
  and _50355_ (_43248_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _50356_ (_43249_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _50357_ (_43250_, _43249_, _43248_);
  and _50358_ (_43251_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _50359_ (_43252_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _50360_ (_43253_, _43252_, _43251_);
  and _50361_ (_43254_, _43253_, _43250_);
  nor _50362_ (_43255_, _43254_, _43113_);
  not _50363_ (_43256_, _39298_);
  and _50364_ (_43257_, _43113_, _43256_);
  nor _50365_ (_43258_, _43257_, _43255_);
  not _50366_ (_43259_, _43258_);
  and _50367_ (_43260_, _43259_, _43096_);
  not _50368_ (_43261_, _43260_);
  and _50369_ (_43262_, _43095_, _43163_);
  and _50370_ (_43263_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _50371_ (_43264_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _50372_ (_43265_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _50373_ (_43266_, _43265_, _43264_);
  and _50374_ (_43267_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _50375_ (_43268_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _50376_ (_43269_, _43268_, _43267_);
  and _50377_ (_43270_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _50378_ (_43271_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _50379_ (_43272_, _43271_, _43270_);
  and _50380_ (_43273_, _43272_, _43269_);
  and _50381_ (_43274_, _43273_, _43266_);
  nor _50382_ (_43275_, _43274_, _43143_);
  nor _50383_ (_43276_, _43275_, _43263_);
  not _50384_ (_43277_, _43276_);
  and _50385_ (_43278_, _43277_, _43139_);
  nor _50386_ (_43279_, _43278_, _43262_);
  not _50387_ (_43280_, _39343_);
  and _50388_ (_43281_, _43280_, _39239_);
  and _50389_ (_43282_, _43136_, _38337_);
  nor _50390_ (_43283_, _43282_, _43281_);
  and _50391_ (_43284_, _43283_, _43279_);
  and _50392_ (_43285_, _43284_, _43261_);
  nor _50393_ (_43286_, _43285_, _43093_);
  and _50394_ (_43287_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _50395_ (_43288_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _50396_ (_43289_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _50397_ (_43290_, _43289_, _43288_);
  and _50398_ (_43291_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _50399_ (_43292_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _50400_ (_43293_, _43292_, _43291_);
  and _50401_ (_43294_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _50402_ (_43295_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _50403_ (_43296_, _43295_, _43294_);
  and _50404_ (_43297_, _43296_, _43293_);
  and _50405_ (_43298_, _43297_, _43290_);
  nor _50406_ (_43299_, _43298_, _43143_);
  nor _50407_ (_43300_, _43299_, _43287_);
  not _50408_ (_43301_, _43300_);
  and _50409_ (_43302_, _43301_, _43139_);
  and _50410_ (_43303_, _43107_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _50411_ (_43304_, _43303_, _39861_);
  not _50412_ (_43305_, _43304_);
  and _50413_ (_43306_, _43305_, _43136_);
  nor _50414_ (_43307_, _43306_, _43302_);
  not _50415_ (_43308_, _39276_);
  and _50416_ (_43309_, _43113_, _43308_);
  and _50417_ (_43310_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _50418_ (_43311_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _50419_ (_43312_, _43311_, _43310_);
  and _50420_ (_43313_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _50421_ (_43314_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _50422_ (_43315_, _43314_, _43313_);
  and _50423_ (_43316_, _43315_, _43312_);
  nor _50424_ (_43317_, _43316_, _43113_);
  nor _50425_ (_43318_, _43317_, _43309_);
  not _50426_ (_43319_, _43318_);
  and _50427_ (_43320_, _43319_, _43096_);
  not _50428_ (_43321_, _43320_);
  not _50429_ (_43322_, _39361_);
  and _50430_ (_43323_, _43322_, _39239_);
  nor _50431_ (_43324_, _43323_, _43164_);
  and _50432_ (_43325_, _43324_, _43321_);
  and _50433_ (_43326_, _43325_, _43307_);
  not _50434_ (_43327_, _43326_);
  and _50435_ (_43328_, _43327_, _43244_);
  nor _50436_ (_43329_, _43328_, _43286_);
  and _50437_ (_43330_, _43113_, _39307_);
  and _50438_ (_43331_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _50439_ (_43332_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor _50440_ (_43333_, _43332_, _43331_);
  and _50441_ (_43334_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _50442_ (_43335_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _50443_ (_43336_, _43335_, _43334_);
  and _50444_ (_43337_, _43336_, _43333_);
  nor _50445_ (_43338_, _43337_, _43113_);
  nor _50446_ (_43339_, _43338_, _43330_);
  not _50447_ (_43340_, _43339_);
  and _50448_ (_43341_, _43340_, _43096_);
  not _50449_ (_43342_, _43341_);
  and _50450_ (_43343_, _43136_, _38124_);
  not _50451_ (_43344_, _43343_);
  not _50452_ (_43345_, _39337_);
  and _50453_ (_43346_, _43345_, _39239_);
  and _50454_ (_43347_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _50455_ (_43348_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _50456_ (_43349_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _50457_ (_43350_, _43349_, _43348_);
  and _50458_ (_43351_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _50459_ (_43352_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _50460_ (_43353_, _43352_, _43351_);
  and _50461_ (_43354_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _50462_ (_43355_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _50463_ (_43356_, _43355_, _43354_);
  and _50464_ (_43357_, _43356_, _43353_);
  and _50465_ (_43358_, _43357_, _43350_);
  nor _50466_ (_43359_, _43358_, _43143_);
  nor _50467_ (_43360_, _43359_, _43347_);
  not _50468_ (_43361_, _43360_);
  and _50469_ (_43362_, _43361_, _43139_);
  nor _50470_ (_43363_, _43362_, _43346_);
  and _50471_ (_43364_, _43363_, _43344_);
  and _50472_ (_43365_, _43364_, _43342_);
  nor _50473_ (_43366_, _43365_, _43093_);
  not _50474_ (_43367_, _39284_);
  and _50475_ (_43368_, _43113_, _43367_);
  and _50476_ (_43369_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _50477_ (_43370_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _50478_ (_43371_, _43370_, _43369_);
  and _50479_ (_43372_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _50480_ (_43373_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _50481_ (_43374_, _43373_, _43372_);
  and _50482_ (_43375_, _43374_, _43371_);
  nor _50483_ (_43376_, _43375_, _43113_);
  nor _50484_ (_43377_, _43376_, _43368_);
  not _50485_ (_43378_, _43377_);
  and _50486_ (_43379_, _43378_, _43096_);
  not _50487_ (_43380_, _43379_);
  not _50488_ (_43381_, _39355_);
  and _50489_ (_43382_, _43381_, _39239_);
  not _50490_ (_43383_, _43382_);
  not _50491_ (_43384_, _43109_);
  and _50492_ (_43385_, _43136_, _43384_);
  and _50493_ (_43386_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _50494_ (_43387_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _50495_ (_43388_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _50496_ (_43389_, _43388_, _43387_);
  and _50497_ (_43390_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _50498_ (_43391_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _50499_ (_43392_, _43391_, _43390_);
  and _50500_ (_43393_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _50501_ (_43394_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _50502_ (_43395_, _43394_, _43393_);
  and _50503_ (_43396_, _43395_, _43392_);
  and _50504_ (_43397_, _43396_, _43389_);
  nor _50505_ (_43398_, _43397_, _43143_);
  nor _50506_ (_43399_, _43398_, _43386_);
  not _50507_ (_43400_, _43399_);
  and _50508_ (_43401_, _43400_, _43139_);
  nor _50509_ (_43402_, _43401_, _43385_);
  and _50510_ (_43403_, _43402_, _43383_);
  and _50511_ (_43404_, _43403_, _43380_);
  not _50512_ (_43405_, _43404_);
  and _50513_ (_43406_, _43405_, _43244_);
  nor _50514_ (_43407_, _43406_, _43366_);
  or _50515_ (_43408_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _50516_ (_43409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _50517_ (_43410_, _43407_, _43409_);
  and _50518_ (_43411_, _43410_, _43408_);
  or _50519_ (_43412_, _43411_, _43329_);
  not _50520_ (_43413_, _43244_);
  and _50521_ (_43414_, _43404_, _43413_);
  not _50522_ (_43415_, _39373_);
  and _50523_ (_43416_, _43415_, _39239_);
  not _50524_ (_43417_, _43416_);
  and _50525_ (_43418_, _43113_, _42899_);
  and _50526_ (_43419_, _43119_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _50527_ (_43420_, _43114_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _50528_ (_43421_, _43420_, _43419_);
  and _50529_ (_43422_, _43121_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _50530_ (_43423_, _43116_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _50531_ (_43424_, _43423_, _43422_);
  and _50532_ (_43425_, _43424_, _43421_);
  nor _50533_ (_43426_, _43425_, _43113_);
  nor _50534_ (_43427_, _43426_, _43418_);
  not _50535_ (_43428_, _43427_);
  and _50536_ (_43429_, _43428_, _43096_);
  not _50537_ (_43430_, _43429_);
  nor _50538_ (_43431_, _43095_, _39105_);
  and _50539_ (_43432_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _50540_ (_43433_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _50541_ (_43434_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _50542_ (_43435_, _43434_, _43433_);
  and _50543_ (_43436_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _50544_ (_43437_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _50545_ (_43438_, _43437_, _43436_);
  and _50546_ (_43439_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _50547_ (_43440_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _50548_ (_43441_, _43440_, _43439_);
  and _50549_ (_43442_, _43441_, _43438_);
  and _50550_ (_43443_, _43442_, _43435_);
  nor _50551_ (_43444_, _43443_, _43143_);
  nor _50552_ (_43445_, _43444_, _43432_);
  not _50553_ (_43446_, _43445_);
  and _50554_ (_43447_, _43446_, _43138_);
  nor _50555_ (_43448_, _43447_, _43431_);
  and _50556_ (_43449_, _43448_, _43430_);
  and _50557_ (_43450_, _43449_, _43417_);
  and _50558_ (_43451_, _43450_, _43244_);
  nor _50559_ (_43452_, _43451_, _43414_);
  not _50560_ (_43453_, _43329_);
  not _50561_ (_43454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _50562_ (_43455_, _43407_, _43454_);
  or _50563_ (_43456_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _50564_ (_43457_, _43456_, _43455_);
  or _50565_ (_43458_, _43457_, _43453_);
  and _50566_ (_43459_, _43458_, _43452_);
  and _50567_ (_43460_, _43459_, _43412_);
  and _50568_ (_43461_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not _50569_ (_43462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor _50570_ (_43463_, _43407_, _43462_);
  or _50571_ (_43464_, _43463_, _43453_);
  or _50572_ (_43465_, _43464_, _43461_);
  not _50573_ (_43466_, _43452_);
  not _50574_ (_43467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _50575_ (_43468_, _43407_, _43467_);
  and _50576_ (_43469_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _50577_ (_43470_, _43469_, _43329_);
  or _50578_ (_43471_, _43470_, _43468_);
  and _50579_ (_43472_, _43471_, _43466_);
  and _50580_ (_43473_, _43472_, _43465_);
  or _50581_ (_43474_, _43473_, _43460_);
  and _50582_ (_43475_, _43474_, _43247_);
  nor _50583_ (_43476_, _28765_, _27745_);
  nor _50584_ (_43477_, _43476_, _31864_);
  not _50585_ (_43478_, _29061_);
  and _50586_ (_43479_, _28765_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50587_ (_43480_, _43479_, _43478_);
  nor _50588_ (_43481_, _28139_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _50589_ (_43482_, _43481_, _43480_);
  nand _50590_ (_43483_, _43482_, _43329_);
  or _50591_ (_43484_, _43482_, _43329_);
  and _50592_ (_43485_, _43484_, _43483_);
  not _50593_ (_43486_, _43485_);
  and _50594_ (_43487_, _43479_, _28929_);
  nor _50595_ (_43488_, _28250_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _50596_ (_43489_, _43488_, _43487_);
  not _50597_ (_43490_, _43489_);
  and _50598_ (_43491_, _43490_, _43407_);
  nor _50599_ (_43492_, _43490_, _43407_);
  nor _50600_ (_43493_, _43492_, _43491_);
  and _50601_ (_43494_, _43493_, _43486_);
  nor _50602_ (_43495_, _43479_, _28929_);
  and _50603_ (_43496_, _43479_, _28490_);
  nor _50604_ (_43497_, _43496_, _43495_);
  not _50605_ (_43498_, _43497_);
  and _50606_ (_43499_, _43498_, _43452_);
  nor _50607_ (_43500_, _43498_, _43452_);
  nor _50608_ (_43501_, _43500_, _43499_);
  and _50609_ (_43502_, _43479_, _39741_);
  nor _50610_ (_43503_, _28008_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _50611_ (_43504_, _43503_, _43502_);
  not _50612_ (_43505_, _43504_);
  nor _50613_ (_43506_, _43505_, _43246_);
  and _50614_ (_43507_, _43505_, _43246_);
  nor _50615_ (_43508_, _43507_, _43506_);
  and _50616_ (_43509_, _43508_, _43501_);
  and _50617_ (_43510_, _43509_, _43494_);
  and _50618_ (_43511_, _43510_, _43477_);
  or _50619_ (_43512_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not _50620_ (_43513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _50621_ (_43514_, _43407_, _43513_);
  and _50622_ (_43515_, _43514_, _43512_);
  or _50623_ (_43516_, _43515_, _43329_);
  not _50624_ (_43517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _50625_ (_43518_, _43407_, _43517_);
  or _50626_ (_43519_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _50627_ (_43520_, _43519_, _43518_);
  or _50628_ (_43521_, _43520_, _43453_);
  and _50629_ (_43522_, _43521_, _43452_);
  and _50630_ (_43523_, _43522_, _43516_);
  and _50631_ (_43524_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not _50632_ (_43525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _50633_ (_43526_, _43407_, _43525_);
  or _50634_ (_43527_, _43526_, _43453_);
  or _50635_ (_43528_, _43527_, _43524_);
  not _50636_ (_43529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _50637_ (_43530_, _43407_, _43529_);
  and _50638_ (_43531_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _50639_ (_43532_, _43531_, _43329_);
  or _50640_ (_43533_, _43532_, _43530_);
  and _50641_ (_43534_, _43533_, _43466_);
  and _50642_ (_43535_, _43534_, _43528_);
  or _50643_ (_43536_, _43535_, _43523_);
  and _50644_ (_43537_, _43536_, _43246_);
  or _50645_ (_43538_, _43537_, _43511_);
  or _50646_ (_43539_, _43538_, _43475_);
  nor _50647_ (_43540_, _43326_, _43244_);
  nor _50648_ (_43541_, _43479_, _29061_);
  not _50649_ (_43542_, _43541_);
  and _50650_ (_43543_, _43542_, _43540_);
  nor _50651_ (_43544_, _43542_, _43540_);
  nor _50652_ (_43545_, _43544_, _43543_);
  and _50653_ (_43546_, _43413_, _43202_);
  nor _50654_ (_43547_, _43479_, _39741_);
  not _50655_ (_43548_, _43547_);
  nor _50656_ (_43549_, _43548_, _43546_);
  and _50657_ (_43550_, _43548_, _43546_);
  nor _50658_ (_43551_, _43550_, _43549_);
  and _50659_ (_43552_, _43551_, _43545_);
  nor _50660_ (_43553_, _43243_, _28776_);
  and _50661_ (_43554_, _43243_, _28776_);
  nor _50662_ (_43555_, _43554_, _43553_);
  nor _50663_ (_43556_, _43450_, _43244_);
  nor _50664_ (_43557_, _43479_, _28490_);
  not _50665_ (_43558_, _43557_);
  and _50666_ (_43559_, _43558_, _43556_);
  nor _50667_ (_43560_, _43558_, _43556_);
  nor _50668_ (_43561_, _43560_, _43559_);
  and _50669_ (_43562_, _43561_, _43555_);
  and _50670_ (_43563_, _43562_, _43552_);
  and _50671_ (_43564_, _43563_, _43511_);
  not _50672_ (_43565_, _43564_);
  or _50673_ (_43566_, _43565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not _50674_ (_43567_, _43511_);
  nor _50675_ (_43568_, _43563_, _43567_);
  nor _50676_ (_43569_, _43568_, rst);
  and _50677_ (_43570_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _50678_ (_43571_, _43570_, _29817_);
  nor _50679_ (_43573_, _43571_, _32431_);
  nor _50680_ (_43574_, _39327_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50681_ (_43576_, _29817_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50682_ (_43578_, _21293_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50683_ (_43579_, _43578_, _43576_);
  or _50684_ (_43581_, _43579_, _43574_);
  or _50685_ (_43583_, _43581_, _43573_);
  and _50686_ (_40752_, _43583_, _43634_);
  or _50687_ (_43586_, _40752_, _43569_);
  and _50688_ (_43587_, _43586_, _43566_);
  and _50689_ (_02564_, _43587_, _43539_);
  not _50690_ (_43588_, _43477_);
  nor _50691_ (_43589_, _43489_, _43588_);
  nor _50692_ (_43590_, _43588_, _43482_);
  and _50693_ (_43591_, _43590_, _43589_);
  and _50694_ (_43592_, _43497_, _43477_);
  nor _50695_ (_43593_, _43588_, _43504_);
  and _50696_ (_43594_, _43593_, _43592_);
  and _50697_ (_43595_, _43594_, _43591_);
  and _50698_ (_43596_, _43583_, _43477_);
  and _50699_ (_43597_, _43596_, _43595_);
  not _50700_ (_43598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _50701_ (_43599_, _43595_, _43598_);
  or _50702_ (_02576_, _43599_, _43597_);
  nor _50703_ (_43600_, _43593_, _43592_);
  nor _50704_ (_43601_, _43590_, _43589_);
  and _50705_ (_43602_, _43601_, _43477_);
  and _50706_ (_43603_, _43602_, _43600_);
  and _50707_ (_43604_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _29806_);
  and _50708_ (_43605_, _43604_, _29850_);
  nand _50709_ (_43606_, _43605_, _32431_);
  not _50710_ (_43607_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50711_ (_43608_, _39306_, _43607_);
  or _50712_ (_43609_, _20140_, _43607_);
  and _50713_ (_43610_, _43609_, _43608_);
  or _50714_ (_43611_, _43610_, _43605_);
  and _50715_ (_43612_, _43611_, _43606_);
  and _50716_ (_43613_, _43612_, _43603_);
  not _50717_ (_43614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _50718_ (_43615_, _43603_, _43614_);
  or _50719_ (_02812_, _43615_, _43613_);
  nand _50720_ (_43616_, _43604_, _29894_);
  nor _50721_ (_43617_, _43616_, _32431_);
  nor _50722_ (_43618_, _39298_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50723_ (_43619_, _43604_, _29916_);
  and _50724_ (_43621_, _43604_, _29817_);
  or _50725_ (_43623_, _43621_, _43570_);
  or _50726_ (_43625_, _43623_, _43619_);
  and _50727_ (_43627_, _43625_, _21119_);
  or _50728_ (_43629_, _43627_, _43618_);
  or _50729_ (_43631_, _43629_, _43617_);
  and _50730_ (_43633_, _43631_, _43603_);
  not _50731_ (_43635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _50732_ (_43636_, _43603_, _43635_);
  or _50733_ (_02816_, _43636_, _43633_);
  not _50734_ (_43639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _50735_ (_43640_, _43603_, _43639_);
  nand _50736_ (_43641_, _43604_, _29927_);
  nor _50737_ (_43642_, _43641_, _32431_);
  nor _50738_ (_43643_, _39291_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50739_ (_43644_, _43604_, _29883_);
  or _50740_ (_43645_, _43644_, _43623_);
  and _50741_ (_43646_, _43645_, _19791_);
  or _50742_ (_43647_, _43646_, _43643_);
  or _50743_ (_43648_, _43647_, _43642_);
  and _50744_ (_43649_, _43648_, _43603_);
  or _50745_ (_02821_, _43649_, _43640_);
  and _50746_ (_43650_, _43621_, _33040_);
  nor _50747_ (_43651_, _39284_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _50748_ (_43652_, _43619_, _43570_);
  or _50749_ (_43653_, _43652_, _43644_);
  and _50750_ (_43654_, _43653_, _20803_);
  or _50751_ (_43655_, _43654_, _43651_);
  or _50752_ (_43656_, _43655_, _43650_);
  and _50753_ (_43657_, _43656_, _43603_);
  not _50754_ (_43658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _50755_ (_43659_, _43603_, _43658_);
  or _50756_ (_02826_, _43659_, _43657_);
  nand _50757_ (_43660_, _43570_, _29850_);
  nor _50758_ (_43661_, _43660_, _32431_);
  nor _50759_ (_43662_, _39276_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50760_ (_43663_, _29850_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50761_ (_43664_, _19977_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50762_ (_43665_, _43664_, _43663_);
  or _50763_ (_43666_, _43665_, _43662_);
  or _50764_ (_43667_, _43666_, _43661_);
  and _50765_ (_43668_, _43667_, _43603_);
  not _50766_ (_43669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _50767_ (_43670_, _43603_, _43669_);
  or _50768_ (_02831_, _43670_, _43668_);
  nand _50769_ (_43671_, _43570_, _29894_);
  nor _50770_ (_43672_, _43671_, _32431_);
  nor _50771_ (_43673_, _39268_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50772_ (_43674_, _29894_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50773_ (_43675_, _20955_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50774_ (_43676_, _43675_, _43674_);
  or _50775_ (_43677_, _43676_, _43673_);
  or _50776_ (_43678_, _43677_, _43672_);
  and _50777_ (_43679_, _43678_, _43603_);
  not _50778_ (_43680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _50779_ (_43681_, _43603_, _43680_);
  or _50780_ (_02835_, _43681_, _43679_);
  nand _50781_ (_43682_, _43570_, _29927_);
  nor _50782_ (_43683_, _43682_, _32431_);
  nor _50783_ (_43684_, _39261_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50784_ (_43685_, _29927_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50785_ (_43686_, _20314_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50786_ (_43687_, _43686_, _43685_);
  or _50787_ (_43688_, _43687_, _43684_);
  or _50788_ (_43689_, _43688_, _43683_);
  and _50789_ (_43690_, _43689_, _43603_);
  not _50790_ (_43691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _50791_ (_43692_, _43603_, _43691_);
  or _50792_ (_02840_, _43692_, _43690_);
  not _50793_ (_43693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _50794_ (_43694_, _43603_, _43693_);
  and _50795_ (_43695_, _43603_, _43583_);
  or _50796_ (_02843_, _43695_, _43694_);
  and _50797_ (_43696_, _43612_, _43477_);
  and _50798_ (_43697_, _43589_, _43482_);
  and _50799_ (_43698_, _43697_, _43600_);
  and _50800_ (_43699_, _43698_, _43696_);
  not _50801_ (_43700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _50802_ (_43701_, _43698_, _43700_);
  or _50803_ (_02850_, _43701_, _43699_);
  and _50804_ (_43702_, _43631_, _43477_);
  and _50805_ (_43703_, _43698_, _43702_);
  not _50806_ (_43704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _50807_ (_43705_, _43698_, _43704_);
  or _50808_ (_02853_, _43705_, _43703_);
  and _50809_ (_43706_, _43648_, _43477_);
  and _50810_ (_43707_, _43698_, _43706_);
  not _50811_ (_43708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _50812_ (_43709_, _43698_, _43708_);
  or _50813_ (_02856_, _43709_, _43707_);
  and _50814_ (_43710_, _43656_, _43477_);
  and _50815_ (_43711_, _43698_, _43710_);
  not _50816_ (_43712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _50817_ (_43713_, _43698_, _43712_);
  or _50818_ (_02861_, _43713_, _43711_);
  and _50819_ (_43714_, _43667_, _43477_);
  and _50820_ (_43715_, _43698_, _43714_);
  not _50821_ (_43716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _50822_ (_43717_, _43698_, _43716_);
  or _50823_ (_02864_, _43717_, _43715_);
  and _50824_ (_43718_, _43678_, _43477_);
  and _50825_ (_43719_, _43698_, _43718_);
  not _50826_ (_43720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _50827_ (_43721_, _43698_, _43720_);
  or _50828_ (_02867_, _43721_, _43719_);
  and _50829_ (_43722_, _43689_, _43477_);
  and _50830_ (_43723_, _43698_, _43722_);
  not _50831_ (_43724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _50832_ (_43725_, _43698_, _43724_);
  or _50833_ (_02870_, _43725_, _43723_);
  and _50834_ (_43726_, _43698_, _43596_);
  nor _50835_ (_43727_, _43698_, _43525_);
  or _50836_ (_02873_, _43727_, _43726_);
  and _50837_ (_43728_, _43590_, _43489_);
  and _50838_ (_43729_, _43728_, _43600_);
  and _50839_ (_43730_, _43729_, _43696_);
  not _50840_ (_43731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _50841_ (_43732_, _43729_, _43731_);
  or _50842_ (_02879_, _43732_, _43730_);
  and _50843_ (_43733_, _43729_, _43702_);
  not _50844_ (_43734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _50845_ (_43735_, _43729_, _43734_);
  or _50846_ (_02883_, _43735_, _43733_);
  and _50847_ (_43736_, _43729_, _43706_);
  not _50848_ (_43737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _50849_ (_43738_, _43729_, _43737_);
  or _50850_ (_02887_, _43738_, _43736_);
  and _50851_ (_43739_, _43729_, _43710_);
  not _50852_ (_43740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _50853_ (_43741_, _43729_, _43740_);
  or _50854_ (_02890_, _43741_, _43739_);
  and _50855_ (_43742_, _43729_, _43714_);
  not _50856_ (_43743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _50857_ (_43744_, _43729_, _43743_);
  or _50858_ (_02895_, _43744_, _43742_);
  and _50859_ (_43745_, _43729_, _43718_);
  not _50860_ (_43746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _50861_ (_43747_, _43729_, _43746_);
  or _50862_ (_02898_, _43747_, _43745_);
  and _50863_ (_43748_, _43729_, _43722_);
  not _50864_ (_43749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _50865_ (_43750_, _43729_, _43749_);
  or _50866_ (_02902_, _43750_, _43748_);
  and _50867_ (_43751_, _43729_, _43596_);
  not _50868_ (_43752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _50869_ (_43753_, _43729_, _43752_);
  or _50870_ (_02905_, _43753_, _43751_);
  and _50871_ (_43754_, _43600_, _43591_);
  and _50872_ (_43755_, _43754_, _43696_);
  not _50873_ (_43756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _50874_ (_43757_, _43754_, _43756_);
  or _50875_ (_02911_, _43757_, _43755_);
  and _50876_ (_43758_, _43754_, _43702_);
  not _50877_ (_43759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _50878_ (_43760_, _43754_, _43759_);
  or _50879_ (_02914_, _43760_, _43758_);
  and _50880_ (_43761_, _43754_, _43706_);
  not _50881_ (_43762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _50882_ (_43763_, _43754_, _43762_);
  or _50883_ (_02918_, _43763_, _43761_);
  and _50884_ (_43764_, _43754_, _43710_);
  not _50885_ (_43765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _50886_ (_43766_, _43754_, _43765_);
  or _50887_ (_02922_, _43766_, _43764_);
  and _50888_ (_43767_, _43754_, _43714_);
  not _50889_ (_43768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _50890_ (_43769_, _43754_, _43768_);
  or _50891_ (_02925_, _43769_, _43767_);
  and _50892_ (_43770_, _43754_, _43718_);
  not _50893_ (_43771_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _50894_ (_43772_, _43754_, _43771_);
  or _50895_ (_02929_, _43772_, _43770_);
  and _50896_ (_43773_, _43754_, _43722_);
  not _50897_ (_43774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _50898_ (_43775_, _43754_, _43774_);
  or _50899_ (_02933_, _43775_, _43773_);
  and _50900_ (_43776_, _43754_, _43596_);
  nor _50901_ (_43777_, _43754_, _43529_);
  or _50902_ (_02936_, _43777_, _43776_);
  and _50903_ (_43778_, _43593_, _43498_);
  and _50904_ (_43779_, _43778_, _43601_);
  and _50905_ (_43780_, _43779_, _43696_);
  not _50906_ (_43781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _50907_ (_43782_, _43779_, _43781_);
  or _50908_ (_02944_, _43782_, _43780_);
  and _50909_ (_43783_, _43779_, _43702_);
  not _50910_ (_43784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _50911_ (_43785_, _43779_, _43784_);
  or _50912_ (_02948_, _43785_, _43783_);
  and _50913_ (_43786_, _43779_, _43706_);
  not _50914_ (_43787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _50915_ (_43788_, _43779_, _43787_);
  or _50916_ (_02951_, _43788_, _43786_);
  and _50917_ (_43789_, _43779_, _43710_);
  not _50918_ (_43790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _50919_ (_43791_, _43779_, _43790_);
  or _50920_ (_02956_, _43791_, _43789_);
  and _50921_ (_43792_, _43779_, _43714_);
  not _50922_ (_43793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _50923_ (_43794_, _43779_, _43793_);
  or _50924_ (_02959_, _43794_, _43792_);
  and _50925_ (_43795_, _43779_, _43718_);
  not _50926_ (_43796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _50927_ (_43797_, _43779_, _43796_);
  or _50928_ (_02963_, _43797_, _43795_);
  and _50929_ (_43798_, _43779_, _43722_);
  not _50930_ (_43799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _50931_ (_43800_, _43779_, _43799_);
  or _50932_ (_02966_, _43800_, _43798_);
  and _50933_ (_43801_, _43779_, _43596_);
  not _50934_ (_43802_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _50935_ (_43803_, _43779_, _43802_);
  or _50936_ (_02970_, _43803_, _43801_);
  and _50937_ (_43804_, _43778_, _43697_);
  and _50938_ (_43805_, _43804_, _43696_);
  not _50939_ (_43806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _50940_ (_43807_, _43804_, _43806_);
  or _50941_ (_02974_, _43807_, _43805_);
  and _50942_ (_43808_, _43804_, _43702_);
  not _50943_ (_43809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _50944_ (_43810_, _43804_, _43809_);
  or _50945_ (_02977_, _43810_, _43808_);
  and _50946_ (_43811_, _43804_, _43706_);
  not _50947_ (_43812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _50948_ (_43813_, _43804_, _43812_);
  or _50949_ (_02982_, _43813_, _43811_);
  and _50950_ (_43814_, _43804_, _43710_);
  not _50951_ (_43815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _50952_ (_43816_, _43804_, _43815_);
  or _50953_ (_02985_, _43816_, _43814_);
  and _50954_ (_43817_, _43804_, _43714_);
  not _50955_ (_43818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _50956_ (_43819_, _43804_, _43818_);
  or _50957_ (_02988_, _43819_, _43817_);
  and _50958_ (_43820_, _43804_, _43718_);
  not _50959_ (_43821_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _50960_ (_43822_, _43804_, _43821_);
  or _50961_ (_02993_, _43822_, _43820_);
  and _50962_ (_43823_, _43804_, _43722_);
  not _50963_ (_43824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _50964_ (_43825_, _43804_, _43824_);
  or _50965_ (_02996_, _43825_, _43823_);
  and _50966_ (_43826_, _43804_, _43596_);
  nor _50967_ (_43827_, _43804_, _43462_);
  or _50968_ (_02999_, _43827_, _43826_);
  and _50969_ (_43828_, _43778_, _43728_);
  and _50970_ (_43829_, _43828_, _43696_);
  not _50971_ (_43830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _50972_ (_43831_, _43828_, _43830_);
  or _50973_ (_03003_, _43831_, _43829_);
  and _50974_ (_43832_, _43828_, _43702_);
  not _50975_ (_43833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _50976_ (_43834_, _43828_, _43833_);
  or _50977_ (_03007_, _43834_, _43832_);
  and _50978_ (_43835_, _43828_, _43706_);
  not _50979_ (_43836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _50980_ (_43837_, _43828_, _43836_);
  or _50981_ (_03010_, _43837_, _43835_);
  and _50982_ (_43838_, _43828_, _43710_);
  not _50983_ (_43839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor _50984_ (_43840_, _43828_, _43839_);
  or _50985_ (_03014_, _43840_, _43838_);
  and _50986_ (_43841_, _43828_, _43714_);
  not _50987_ (_43842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _50988_ (_43843_, _43828_, _43842_);
  or _50989_ (_03018_, _43843_, _43841_);
  and _50990_ (_43844_, _43828_, _43718_);
  not _50991_ (_43845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _50992_ (_43846_, _43828_, _43845_);
  or _50993_ (_03021_, _43846_, _43844_);
  and _50994_ (_43847_, _43828_, _43722_);
  not _50995_ (_43848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _50996_ (_43849_, _43828_, _43848_);
  or _50997_ (_03024_, _43849_, _43847_);
  and _50998_ (_43850_, _43828_, _43596_);
  not _50999_ (_43851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _51000_ (_43852_, _43828_, _43851_);
  or _51001_ (_03027_, _43852_, _43850_);
  and _51002_ (_43853_, _43778_, _43591_);
  and _51003_ (_43854_, _43853_, _43696_);
  not _51004_ (_43855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _51005_ (_43856_, _43853_, _43855_);
  or _51006_ (_03032_, _43856_, _43854_);
  and _51007_ (_43857_, _43853_, _43702_);
  not _51008_ (_43858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _51009_ (_43859_, _43853_, _43858_);
  or _51010_ (_03035_, _43859_, _43857_);
  and _51011_ (_43860_, _43853_, _43706_);
  not _51012_ (_43861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _51013_ (_43862_, _43853_, _43861_);
  or _51014_ (_03038_, _43862_, _43860_);
  and _51015_ (_43863_, _43853_, _43710_);
  not _51016_ (_43864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _51017_ (_43865_, _43853_, _43864_);
  or _51018_ (_03042_, _43865_, _43863_);
  and _51019_ (_43866_, _43853_, _43714_);
  not _51020_ (_43867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _51021_ (_43868_, _43853_, _43867_);
  or _51022_ (_03045_, _43868_, _43866_);
  and _51023_ (_43869_, _43853_, _43718_);
  not _51024_ (_43870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _51025_ (_43871_, _43853_, _43870_);
  or _51026_ (_03048_, _43871_, _43869_);
  and _51027_ (_43872_, _43853_, _43722_);
  not _51028_ (_43873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _51029_ (_43874_, _43853_, _43873_);
  or _51030_ (_03051_, _43874_, _43872_);
  and _51031_ (_43875_, _43853_, _43596_);
  nor _51032_ (_43876_, _43853_, _43467_);
  or _51033_ (_03054_, _43876_, _43875_);
  and _51034_ (_43877_, _43592_, _43504_);
  and _51035_ (_43878_, _43877_, _43601_);
  and _51036_ (_43879_, _43878_, _43696_);
  not _51037_ (_43880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _51038_ (_43881_, _43878_, _43880_);
  or _51039_ (_03060_, _43881_, _43879_);
  and _51040_ (_43882_, _43878_, _43702_);
  not _51041_ (_43883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _51042_ (_43884_, _43878_, _43883_);
  or _51043_ (_03063_, _43884_, _43882_);
  and _51044_ (_43885_, _43878_, _43706_);
  not _51045_ (_43886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _51046_ (_43887_, _43878_, _43886_);
  or _51047_ (_03067_, _43887_, _43885_);
  and _51048_ (_43888_, _43878_, _43710_);
  not _51049_ (_43889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _51050_ (_43890_, _43878_, _43889_);
  or _51051_ (_03069_, _43890_, _43888_);
  and _51052_ (_43891_, _43878_, _43714_);
  not _51053_ (_43892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _51054_ (_43893_, _43878_, _43892_);
  or _51055_ (_03073_, _43893_, _43891_);
  and _51056_ (_43894_, _43878_, _43718_);
  not _51057_ (_43895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _51058_ (_43896_, _43878_, _43895_);
  or _51059_ (_03076_, _43896_, _43894_);
  and _51060_ (_43897_, _43878_, _43722_);
  not _51061_ (_43898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _51062_ (_43899_, _43878_, _43898_);
  or _51063_ (_03080_, _43899_, _43897_);
  and _51064_ (_43900_, _43878_, _43596_);
  nor _51065_ (_43901_, _43878_, _43517_);
  or _51066_ (_03083_, _43901_, _43900_);
  and _51067_ (_43902_, _43877_, _43697_);
  and _51068_ (_43903_, _43902_, _43696_);
  not _51069_ (_43904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _51070_ (_43905_, _43902_, _43904_);
  or _51071_ (_03087_, _43905_, _43903_);
  and _51072_ (_43906_, _43902_, _43702_);
  not _51073_ (_43907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _51074_ (_43908_, _43902_, _43907_);
  or _51075_ (_03091_, _43908_, _43906_);
  and _51076_ (_43909_, _43902_, _43706_);
  not _51077_ (_43910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _51078_ (_43911_, _43902_, _43910_);
  or _51079_ (_03095_, _43911_, _43909_);
  and _51080_ (_43912_, _43902_, _43710_);
  not _51081_ (_43913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _51082_ (_43914_, _43902_, _43913_);
  or _51083_ (_03099_, _43914_, _43912_);
  and _51084_ (_43915_, _43902_, _43714_);
  not _51085_ (_43916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _51086_ (_43917_, _43902_, _43916_);
  or _51087_ (_03102_, _43917_, _43915_);
  and _51088_ (_43918_, _43902_, _43718_);
  not _51089_ (_43919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _51090_ (_43920_, _43902_, _43919_);
  or _51091_ (_03106_, _43920_, _43918_);
  and _51092_ (_43921_, _43902_, _43722_);
  not _51093_ (_43922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _51094_ (_43923_, _43902_, _43922_);
  or _51095_ (_03109_, _43923_, _43921_);
  and _51096_ (_43924_, _43902_, _43596_);
  not _51097_ (_43925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _51098_ (_43926_, _43902_, _43925_);
  or _51099_ (_03112_, _43926_, _43924_);
  and _51100_ (_43927_, _43877_, _43728_);
  and _51101_ (_43928_, _43927_, _43696_);
  not _51102_ (_43929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _51103_ (_43930_, _43927_, _43929_);
  or _51104_ (_03116_, _43930_, _43928_);
  and _51105_ (_43931_, _43927_, _43702_);
  not _51106_ (_43932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _51107_ (_43933_, _43927_, _43932_);
  or _51108_ (_03119_, _43933_, _43931_);
  and _51109_ (_43934_, _43927_, _43706_);
  not _51110_ (_43935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _51111_ (_43936_, _43927_, _43935_);
  or _51112_ (_03122_, _43936_, _43934_);
  and _51113_ (_43937_, _43927_, _43710_);
  not _51114_ (_43938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _51115_ (_43939_, _43927_, _43938_);
  or _51116_ (_03125_, _43939_, _43937_);
  and _51117_ (_43940_, _43927_, _43714_);
  not _51118_ (_43941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _51119_ (_43942_, _43927_, _43941_);
  or _51120_ (_03130_, _43942_, _43940_);
  and _51121_ (_43943_, _43927_, _43718_);
  not _51122_ (_43944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _51123_ (_43945_, _43927_, _43944_);
  or _51124_ (_03133_, _43945_, _43943_);
  and _51125_ (_43946_, _43927_, _43722_);
  not _51126_ (_43947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _51127_ (_43948_, _43927_, _43947_);
  or _51128_ (_03136_, _43948_, _43946_);
  and _51129_ (_43949_, _43927_, _43596_);
  nor _51130_ (_43950_, _43927_, _43513_);
  or _51131_ (_03139_, _43950_, _43949_);
  and _51132_ (_43951_, _43877_, _43591_);
  and _51133_ (_43952_, _43951_, _43696_);
  not _51134_ (_43953_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _51135_ (_43954_, _43951_, _43953_);
  or _51136_ (_03143_, _43954_, _43952_);
  and _51137_ (_43955_, _43951_, _43702_);
  not _51138_ (_43956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _51139_ (_43957_, _43951_, _43956_);
  or _51140_ (_03147_, _43957_, _43955_);
  and _51141_ (_43958_, _43951_, _43706_);
  not _51142_ (_43959_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _51143_ (_43960_, _43951_, _43959_);
  or _51144_ (_03150_, _43960_, _43958_);
  and _51145_ (_43961_, _43951_, _43710_);
  not _51146_ (_43962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _51147_ (_43963_, _43951_, _43962_);
  or _51148_ (_03154_, _43963_, _43961_);
  and _51149_ (_43964_, _43951_, _43714_);
  not _51150_ (_43965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _51151_ (_43966_, _43951_, _43965_);
  or _51152_ (_03157_, _43966_, _43964_);
  and _51153_ (_43967_, _43951_, _43718_);
  not _51154_ (_43968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _51155_ (_43969_, _43951_, _43968_);
  or _51156_ (_03161_, _43969_, _43967_);
  and _51157_ (_43970_, _43951_, _43722_);
  not _51158_ (_43971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _51159_ (_43972_, _43951_, _43971_);
  or _51160_ (_03164_, _43972_, _43970_);
  and _51161_ (_43973_, _43951_, _43596_);
  not _51162_ (_43974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _51163_ (_43975_, _43951_, _43974_);
  or _51164_ (_03167_, _43975_, _43973_);
  and _51165_ (_43976_, _43601_, _43594_);
  and _51166_ (_43977_, _43976_, _43696_);
  not _51167_ (_43978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _51168_ (_43979_, _43976_, _43978_);
  or _51169_ (_03172_, _43979_, _43977_);
  and _51170_ (_43980_, _43976_, _43702_);
  not _51171_ (_43981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _51172_ (_43982_, _43976_, _43981_);
  or _51173_ (_03176_, _43982_, _43980_);
  and _51174_ (_43983_, _43976_, _43706_);
  not _51175_ (_43984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _51176_ (_43985_, _43976_, _43984_);
  or _51177_ (_03180_, _43985_, _43983_);
  and _51178_ (_43986_, _43976_, _43710_);
  not _51179_ (_43987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _51180_ (_43988_, _43976_, _43987_);
  or _51181_ (_03183_, _43988_, _43986_);
  and _51182_ (_43989_, _43976_, _43714_);
  not _51183_ (_43990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _51184_ (_43991_, _43976_, _43990_);
  or _51185_ (_03187_, _43991_, _43989_);
  and _51186_ (_43992_, _43976_, _43718_);
  not _51187_ (_43993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _51188_ (_43994_, _43976_, _43993_);
  or _51189_ (_03190_, _43994_, _43992_);
  and _51190_ (_43995_, _43976_, _43722_);
  not _51191_ (_43996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _51192_ (_43997_, _43976_, _43996_);
  or _51193_ (_03194_, _43997_, _43995_);
  and _51194_ (_43998_, _43976_, _43596_);
  nor _51195_ (_43999_, _43976_, _43454_);
  or _51196_ (_03197_, _43999_, _43998_);
  and _51197_ (_44000_, _43697_, _43594_);
  and _51198_ (_44001_, _44000_, _43696_);
  not _51199_ (_44002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _51200_ (_44003_, _44000_, _44002_);
  or _51201_ (_03201_, _44003_, _44001_);
  and _51202_ (_44004_, _44000_, _43702_);
  not _51203_ (_44005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _51204_ (_44006_, _44000_, _44005_);
  or _51205_ (_03205_, _44006_, _44004_);
  and _51206_ (_44007_, _44000_, _43706_);
  not _51207_ (_44008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _51208_ (_44009_, _44000_, _44008_);
  or _51209_ (_03208_, _44009_, _44007_);
  and _51210_ (_44010_, _44000_, _43710_);
  not _51211_ (_44011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _51212_ (_44012_, _44000_, _44011_);
  or _51213_ (_03212_, _44012_, _44010_);
  and _51214_ (_44013_, _44000_, _43714_);
  not _51215_ (_44014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _51216_ (_44015_, _44000_, _44014_);
  or _51217_ (_03215_, _44015_, _44013_);
  and _51218_ (_44016_, _44000_, _43718_);
  not _51219_ (_44017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _51220_ (_44018_, _44000_, _44017_);
  or _51221_ (_03219_, _44018_, _44016_);
  and _51222_ (_44019_, _44000_, _43722_);
  not _51223_ (_44020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _51224_ (_44021_, _44000_, _44020_);
  or _51225_ (_03222_, _44021_, _44019_);
  and _51226_ (_44022_, _44000_, _43596_);
  not _51227_ (_44023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _51228_ (_44024_, _44000_, _44023_);
  or _51229_ (_03225_, _44024_, _44022_);
  and _51230_ (_44025_, _43728_, _43594_);
  and _51231_ (_44026_, _44025_, _43696_);
  not _51232_ (_44027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _51233_ (_44028_, _44025_, _44027_);
  or _51234_ (_03230_, _44028_, _44026_);
  and _51235_ (_44029_, _44025_, _43702_);
  not _51236_ (_44030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _51237_ (_44031_, _44025_, _44030_);
  or _51238_ (_03233_, _44031_, _44029_);
  and _51239_ (_44032_, _44025_, _43706_);
  not _51240_ (_44033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _51241_ (_44034_, _44025_, _44033_);
  or _51242_ (_03237_, _44034_, _44032_);
  and _51243_ (_44035_, _44025_, _43710_);
  not _51244_ (_44036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _51245_ (_44037_, _44025_, _44036_);
  or _51246_ (_03240_, _44037_, _44035_);
  and _51247_ (_44038_, _44025_, _43714_);
  not _51248_ (_44039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _51249_ (_44040_, _44025_, _44039_);
  or _51250_ (_03244_, _44040_, _44038_);
  and _51251_ (_44041_, _44025_, _43718_);
  not _51252_ (_44042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _51253_ (_44043_, _44025_, _44042_);
  or _51254_ (_03247_, _44043_, _44041_);
  and _51255_ (_44044_, _44025_, _43722_);
  not _51256_ (_44045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _51257_ (_44046_, _44025_, _44045_);
  or _51258_ (_03251_, _44046_, _44044_);
  and _51259_ (_44047_, _44025_, _43596_);
  nor _51260_ (_44048_, _44025_, _43409_);
  or _51261_ (_03254_, _44048_, _44047_);
  and _51262_ (_44049_, _43696_, _43595_);
  not _51263_ (_44050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _51264_ (_44051_, _43595_, _44050_);
  or _51265_ (_03258_, _44051_, _44049_);
  and _51266_ (_44052_, _43702_, _43595_);
  not _51267_ (_44053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _51268_ (_44054_, _43595_, _44053_);
  or _51269_ (_03262_, _44054_, _44052_);
  and _51270_ (_44055_, _43706_, _43595_);
  not _51271_ (_44056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _51272_ (_44057_, _43595_, _44056_);
  or _51273_ (_03265_, _44057_, _44055_);
  and _51274_ (_44058_, _43710_, _43595_);
  not _51275_ (_44059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _51276_ (_44060_, _43595_, _44059_);
  or _51277_ (_03269_, _44060_, _44058_);
  and _51278_ (_44061_, _43714_, _43595_);
  not _51279_ (_44062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _51280_ (_44063_, _43595_, _44062_);
  or _51281_ (_03273_, _44063_, _44061_);
  and _51282_ (_44064_, _43718_, _43595_);
  not _51283_ (_44065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _51284_ (_44066_, _43595_, _44065_);
  or _51285_ (_03276_, _44066_, _44064_);
  and _51286_ (_44067_, _43722_, _43595_);
  not _51287_ (_44068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _51288_ (_44069_, _43595_, _44068_);
  or _51289_ (_03279_, _44069_, _44067_);
  and _51290_ (_44070_, _43563_, _43510_);
  and _51291_ (_44071_, _44070_, _43477_);
  not _51292_ (_44072_, _44071_);
  nor _51293_ (_44073_, _43407_, _43756_);
  and _51294_ (_44074_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _51295_ (_44075_, _44074_, _43329_);
  or _51296_ (_44076_, _44075_, _44073_);
  and _51297_ (_44077_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _51298_ (_44078_, _43407_, _43700_);
  or _51299_ (_44079_, _44078_, _43453_);
  or _51300_ (_44080_, _44079_, _44077_);
  and _51301_ (_44081_, _44080_, _44076_);
  or _51302_ (_44082_, _44081_, _43247_);
  nor _51303_ (_44083_, _43407_, _43855_);
  and _51304_ (_44084_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _51305_ (_44085_, _44084_, _43329_);
  or _51306_ (_44086_, _44085_, _44083_);
  and _51307_ (_44087_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _51308_ (_44088_, _43407_, _43806_);
  or _51309_ (_44089_, _44088_, _43453_);
  or _51310_ (_44090_, _44089_, _44087_);
  and _51311_ (_44091_, _44090_, _44086_);
  or _51312_ (_44092_, _44091_, _43246_);
  and _51313_ (_44093_, _44092_, _43466_);
  and _51314_ (_44094_, _44093_, _44082_);
  nand _51315_ (_44095_, _43407_, _43880_);
  or _51316_ (_44096_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _51317_ (_44097_, _44096_, _44095_);
  or _51318_ (_44098_, _44097_, _43453_);
  or _51319_ (_44099_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand _51320_ (_44100_, _43407_, _43929_);
  and _51321_ (_44101_, _44100_, _44099_);
  or _51322_ (_44102_, _44101_, _43329_);
  and _51323_ (_44103_, _44102_, _44098_);
  or _51324_ (_44104_, _44103_, _43247_);
  nand _51325_ (_44105_, _43407_, _43978_);
  or _51326_ (_44106_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _51327_ (_44107_, _44106_, _44105_);
  or _51328_ (_44108_, _44107_, _43453_);
  or _51329_ (_44109_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand _51330_ (_44110_, _43407_, _44027_);
  and _51331_ (_44111_, _44110_, _44109_);
  or _51332_ (_44112_, _44111_, _43329_);
  and _51333_ (_44113_, _44112_, _44108_);
  or _51334_ (_44114_, _44113_, _43246_);
  and _51335_ (_44120_, _44114_, _43452_);
  and _51336_ (_44124_, _44120_, _44104_);
  or _51337_ (_44131_, _44124_, _44094_);
  and _51338_ (_44139_, _44131_, _44072_);
  and _51339_ (_44143_, _43564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or _51340_ (_44148_, _44143_, _43568_);
  or _51341_ (_44156_, _44148_, _44139_);
  and _51342_ (_40772_, _43612_, _43634_);
  or _51343_ (_44165_, _40772_, _43569_);
  and _51344_ (_05076_, _44165_, _44156_);
  nor _51345_ (_44179_, _43407_, _43759_);
  and _51346_ (_44183_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _51347_ (_44188_, _44183_, _43329_);
  or _51348_ (_44196_, _44188_, _44179_);
  and _51349_ (_44202_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _51350_ (_44205_, _43407_, _43704_);
  or _51351_ (_44209_, _44205_, _43453_);
  or _51352_ (_44220_, _44209_, _44202_);
  and _51353_ (_44224_, _44220_, _44196_);
  or _51354_ (_44231_, _44224_, _43247_);
  nor _51355_ (_44239_, _43407_, _43858_);
  and _51356_ (_44243_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _51357_ (_44248_, _44243_, _43329_);
  or _51358_ (_44256_, _44248_, _44239_);
  and _51359_ (_44262_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _51360_ (_44266_, _43407_, _43809_);
  or _51361_ (_44273_, _44266_, _43453_);
  or _51362_ (_44281_, _44273_, _44262_);
  and _51363_ (_44285_, _44281_, _44256_);
  or _51364_ (_44290_, _44285_, _43246_);
  and _51365_ (_44298_, _44290_, _43466_);
  and _51366_ (_44304_, _44298_, _44231_);
  nand _51367_ (_44308_, _43407_, _43883_);
  or _51368_ (_44315_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _51369_ (_44323_, _44315_, _44308_);
  or _51370_ (_44327_, _44323_, _43453_);
  or _51371_ (_44332_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand _51372_ (_44340_, _43407_, _43932_);
  and _51373_ (_44341_, _44340_, _44332_);
  or _51374_ (_44342_, _44341_, _43329_);
  and _51375_ (_44343_, _44342_, _44327_);
  or _51376_ (_44344_, _44343_, _43247_);
  nand _51377_ (_44345_, _43407_, _43981_);
  or _51378_ (_44346_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _51379_ (_44347_, _44346_, _44345_);
  or _51380_ (_44348_, _44347_, _43453_);
  or _51381_ (_44349_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand _51382_ (_44350_, _43407_, _44030_);
  and _51383_ (_44351_, _44350_, _44349_);
  or _51384_ (_44352_, _44351_, _43329_);
  and _51385_ (_44353_, _44352_, _44348_);
  or _51386_ (_44354_, _44353_, _43246_);
  and _51387_ (_44355_, _44354_, _43452_);
  and _51388_ (_44356_, _44355_, _44344_);
  or _51389_ (_44357_, _44356_, _44304_);
  and _51390_ (_44358_, _44357_, _44072_);
  and _51391_ (_44359_, _43564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _51392_ (_44360_, _44359_, _43568_);
  or _51393_ (_44361_, _44360_, _44358_);
  and _51394_ (_40773_, _43631_, _43634_);
  or _51395_ (_44362_, _40773_, _43569_);
  and _51396_ (_05078_, _44362_, _44361_);
  nor _51397_ (_44363_, _43407_, _43762_);
  and _51398_ (_44364_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _51399_ (_44365_, _44364_, _43329_);
  or _51400_ (_44366_, _44365_, _44363_);
  and _51401_ (_44367_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _51402_ (_44368_, _43407_, _43708_);
  or _51403_ (_44369_, _44368_, _43453_);
  or _51404_ (_44370_, _44369_, _44367_);
  and _51405_ (_44371_, _44370_, _44366_);
  or _51406_ (_44372_, _44371_, _43247_);
  nor _51407_ (_44373_, _43407_, _43861_);
  and _51408_ (_44374_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _51409_ (_44375_, _44374_, _43329_);
  or _51410_ (_44376_, _44375_, _44373_);
  and _51411_ (_44377_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _51412_ (_44378_, _43407_, _43812_);
  or _51413_ (_44379_, _44378_, _43453_);
  or _51414_ (_44380_, _44379_, _44377_);
  and _51415_ (_44381_, _44380_, _44376_);
  or _51416_ (_44382_, _44381_, _43246_);
  and _51417_ (_44383_, _44382_, _43466_);
  and _51418_ (_44384_, _44383_, _44372_);
  nand _51419_ (_44385_, _43407_, _43886_);
  or _51420_ (_44386_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _51421_ (_44387_, _44386_, _44385_);
  or _51422_ (_44388_, _44387_, _43453_);
  or _51423_ (_44389_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _51424_ (_44390_, _43407_, _43935_);
  and _51425_ (_44391_, _44390_, _44389_);
  or _51426_ (_44392_, _44391_, _43329_);
  and _51427_ (_44393_, _44392_, _44388_);
  or _51428_ (_44394_, _44393_, _43247_);
  nand _51429_ (_44395_, _43407_, _43984_);
  or _51430_ (_44396_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _51431_ (_44397_, _44396_, _44395_);
  or _51432_ (_44398_, _44397_, _43453_);
  or _51433_ (_44399_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _51434_ (_44400_, _43407_, _44033_);
  and _51435_ (_44401_, _44400_, _44399_);
  or _51436_ (_44402_, _44401_, _43329_);
  and _51437_ (_44403_, _44402_, _44398_);
  or _51438_ (_44404_, _44403_, _43246_);
  and _51439_ (_44405_, _44404_, _43452_);
  and _51440_ (_44406_, _44405_, _44394_);
  or _51441_ (_44407_, _44406_, _44384_);
  or _51442_ (_44408_, _44407_, _43564_);
  or _51443_ (_44409_, _43565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _51444_ (_44410_, _44409_, _43569_);
  and _51445_ (_44411_, _44410_, _44408_);
  and _51446_ (_40774_, _43648_, _43634_);
  and _51447_ (_44412_, _40774_, _43568_);
  or _51448_ (_05080_, _44412_, _44411_);
  nor _51449_ (_44413_, _43407_, _43765_);
  and _51450_ (_44414_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _51451_ (_44415_, _44414_, _43329_);
  or _51452_ (_44416_, _44415_, _44413_);
  and _51453_ (_44417_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _51454_ (_44418_, _43407_, _43712_);
  or _51455_ (_44419_, _44418_, _43453_);
  or _51456_ (_44420_, _44419_, _44417_);
  and _51457_ (_44421_, _44420_, _44416_);
  or _51458_ (_44422_, _44421_, _43247_);
  nor _51459_ (_44423_, _43407_, _43864_);
  and _51460_ (_44424_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _51461_ (_44425_, _44424_, _43329_);
  or _51462_ (_44426_, _44425_, _44423_);
  and _51463_ (_44427_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _51464_ (_44428_, _43407_, _43815_);
  or _51465_ (_44429_, _44428_, _43453_);
  or _51466_ (_44430_, _44429_, _44427_);
  and _51467_ (_44431_, _44430_, _44426_);
  or _51468_ (_44432_, _44431_, _43246_);
  and _51469_ (_44433_, _44432_, _43466_);
  and _51470_ (_44434_, _44433_, _44422_);
  nand _51471_ (_44435_, _43407_, _43889_);
  or _51472_ (_44436_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _51473_ (_44437_, _44436_, _44435_);
  or _51474_ (_44438_, _44437_, _43453_);
  or _51475_ (_44439_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _51476_ (_44440_, _43407_, _43938_);
  and _51477_ (_44441_, _44440_, _44439_);
  or _51478_ (_44442_, _44441_, _43329_);
  and _51479_ (_44443_, _44442_, _44438_);
  or _51480_ (_44444_, _44443_, _43247_);
  nand _51481_ (_44445_, _43407_, _43987_);
  or _51482_ (_44446_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _51483_ (_44447_, _44446_, _44445_);
  or _51484_ (_44448_, _44447_, _43453_);
  or _51485_ (_44449_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _51486_ (_44450_, _43407_, _44036_);
  and _51487_ (_44451_, _44450_, _44449_);
  or _51488_ (_44452_, _44451_, _43329_);
  and _51489_ (_44453_, _44452_, _44448_);
  or _51490_ (_44454_, _44453_, _43246_);
  and _51491_ (_44455_, _44454_, _43452_);
  and _51492_ (_44456_, _44455_, _44444_);
  or _51493_ (_44457_, _44456_, _44434_);
  and _51494_ (_44458_, _44457_, _44072_);
  and _51495_ (_44459_, _43564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _51496_ (_44460_, _44459_, _43568_);
  or _51497_ (_44461_, _44460_, _44458_);
  and _51498_ (_40775_, _43656_, _43634_);
  or _51499_ (_44462_, _40775_, _43569_);
  and _51500_ (_05082_, _44462_, _44461_);
  and _51501_ (_44463_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _51502_ (_44464_, _43407_, _43716_);
  or _51503_ (_44465_, _44464_, _43453_);
  or _51504_ (_44466_, _44465_, _44463_);
  nor _51505_ (_44467_, _43407_, _43768_);
  and _51506_ (_44468_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _51507_ (_44469_, _44468_, _43329_);
  or _51508_ (_44470_, _44469_, _44467_);
  and _51509_ (_44471_, _44470_, _44466_);
  or _51510_ (_44472_, _44471_, _43247_);
  nor _51511_ (_44473_, _43407_, _43867_);
  and _51512_ (_44474_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _51513_ (_44475_, _44474_, _43329_);
  or _51514_ (_44476_, _44475_, _44473_);
  and _51515_ (_44477_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _51516_ (_44478_, _43407_, _43818_);
  or _51517_ (_44479_, _44478_, _43453_);
  or _51518_ (_44480_, _44479_, _44477_);
  and _51519_ (_44481_, _44480_, _44476_);
  or _51520_ (_44482_, _44481_, _43246_);
  and _51521_ (_44483_, _44482_, _43466_);
  and _51522_ (_44484_, _44483_, _44472_);
  nor _51523_ (_44485_, _43407_, _43965_);
  and _51524_ (_44486_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _51525_ (_44487_, _44486_, _43329_);
  or _51526_ (_44488_, _44487_, _44485_);
  and _51527_ (_44489_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _51528_ (_44490_, _43407_, _43916_);
  or _51529_ (_44491_, _44490_, _43453_);
  or _51530_ (_44492_, _44491_, _44489_);
  and _51531_ (_44493_, _44492_, _44488_);
  or _51532_ (_44494_, _44493_, _43247_);
  nor _51533_ (_44495_, _43407_, _44062_);
  and _51534_ (_44496_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _51535_ (_44497_, _44496_, _43329_);
  or _51536_ (_44498_, _44497_, _44495_);
  and _51537_ (_44499_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _51538_ (_44500_, _43407_, _44014_);
  or _51539_ (_44501_, _44500_, _43453_);
  or _51540_ (_44502_, _44501_, _44499_);
  and _51541_ (_44503_, _44502_, _44498_);
  or _51542_ (_44504_, _44503_, _43246_);
  and _51543_ (_44505_, _44504_, _43452_);
  and _51544_ (_44506_, _44505_, _44494_);
  or _51545_ (_44507_, _44506_, _44484_);
  and _51546_ (_44508_, _44507_, _43567_);
  and _51547_ (_44509_, _43667_, _43568_);
  and _51548_ (_44510_, _43564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _51549_ (_44511_, _44510_, _44509_);
  or _51550_ (_44512_, _44511_, _44508_);
  and _51551_ (_05084_, _44512_, _43634_);
  nor _51552_ (_44513_, _43407_, _43771_);
  and _51553_ (_44514_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _51554_ (_44515_, _44514_, _43329_);
  or _51555_ (_44516_, _44515_, _44513_);
  and _51556_ (_44517_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _51557_ (_44518_, _43407_, _43720_);
  or _51558_ (_44519_, _44518_, _43453_);
  or _51559_ (_44520_, _44519_, _44517_);
  and _51560_ (_44521_, _44520_, _44516_);
  or _51561_ (_44522_, _44521_, _43247_);
  nor _51562_ (_44523_, _43407_, _43870_);
  and _51563_ (_44524_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _51564_ (_44525_, _44524_, _43329_);
  or _51565_ (_44526_, _44525_, _44523_);
  and _51566_ (_44527_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _51567_ (_44528_, _43407_, _43821_);
  or _51568_ (_44529_, _44528_, _43453_);
  or _51569_ (_44530_, _44529_, _44527_);
  and _51570_ (_44531_, _44530_, _44526_);
  or _51571_ (_44532_, _44531_, _43246_);
  and _51572_ (_44533_, _44532_, _43466_);
  and _51573_ (_44534_, _44533_, _44522_);
  nand _51574_ (_44535_, _43407_, _43895_);
  or _51575_ (_44536_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _51576_ (_44537_, _44536_, _44535_);
  or _51577_ (_44538_, _44537_, _43453_);
  or _51578_ (_44539_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _51579_ (_44540_, _43407_, _43944_);
  and _51580_ (_44541_, _44540_, _44539_);
  or _51581_ (_44542_, _44541_, _43329_);
  and _51582_ (_44543_, _44542_, _44538_);
  or _51583_ (_44544_, _44543_, _43247_);
  nand _51584_ (_44545_, _43407_, _43993_);
  or _51585_ (_44546_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _51586_ (_44547_, _44546_, _44545_);
  or _51587_ (_44548_, _44547_, _43453_);
  or _51588_ (_44549_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _51589_ (_44550_, _43407_, _44042_);
  and _51590_ (_44551_, _44550_, _44549_);
  or _51591_ (_44552_, _44551_, _43329_);
  and _51592_ (_44553_, _44552_, _44548_);
  or _51593_ (_44554_, _44553_, _43246_);
  and _51594_ (_44555_, _44554_, _43452_);
  and _51595_ (_44556_, _44555_, _44544_);
  or _51596_ (_44557_, _44556_, _44534_);
  or _51597_ (_44558_, _44557_, _43564_);
  or _51598_ (_44559_, _43565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _51599_ (_44560_, _44559_, _43569_);
  and _51600_ (_44561_, _44560_, _44558_);
  and _51601_ (_40777_, _43678_, _43634_);
  and _51602_ (_44562_, _40777_, _43568_);
  or _51603_ (_05086_, _44562_, _44561_);
  nor _51604_ (_44563_, _43407_, _43774_);
  and _51605_ (_44564_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _51606_ (_44565_, _44564_, _43329_);
  or _51607_ (_44566_, _44565_, _44563_);
  and _51608_ (_44567_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _51609_ (_44568_, _43407_, _43724_);
  or _51610_ (_44569_, _44568_, _43453_);
  or _51611_ (_44570_, _44569_, _44567_);
  and _51612_ (_44571_, _44570_, _44566_);
  or _51613_ (_44572_, _44571_, _43247_);
  nor _51614_ (_44573_, _43407_, _43873_);
  and _51615_ (_44574_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _51616_ (_44575_, _44574_, _43329_);
  or _51617_ (_44576_, _44575_, _44573_);
  and _51618_ (_44577_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _51619_ (_44578_, _43407_, _43824_);
  or _51620_ (_44579_, _44578_, _43453_);
  or _51621_ (_44580_, _44579_, _44577_);
  and _51622_ (_44581_, _44580_, _44576_);
  or _51623_ (_44582_, _44581_, _43246_);
  and _51624_ (_44583_, _44582_, _43466_);
  and _51625_ (_44584_, _44583_, _44572_);
  nand _51626_ (_44585_, _43407_, _43898_);
  or _51627_ (_44586_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _51628_ (_44587_, _44586_, _44585_);
  or _51629_ (_44588_, _44587_, _43453_);
  or _51630_ (_44589_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _51631_ (_44590_, _43407_, _43947_);
  and _51632_ (_00006_, _44590_, _44589_);
  or _51633_ (_00007_, _00006_, _43329_);
  and _51634_ (_00008_, _00007_, _44588_);
  or _51635_ (_00009_, _00008_, _43247_);
  nand _51636_ (_00010_, _43407_, _43996_);
  or _51637_ (_00011_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _51638_ (_00012_, _00011_, _00010_);
  or _51639_ (_00013_, _00012_, _43453_);
  or _51640_ (_00014_, _43407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _51641_ (_00015_, _43407_, _44045_);
  and _51642_ (_00016_, _00015_, _00014_);
  or _51643_ (_00017_, _00016_, _43329_);
  and _51644_ (_00018_, _00017_, _00013_);
  or _51645_ (_00019_, _00018_, _43246_);
  and _51646_ (_00020_, _00019_, _43452_);
  and _51647_ (_00021_, _00020_, _00009_);
  or _51648_ (_00022_, _00021_, _44584_);
  or _51649_ (_00023_, _00022_, _43564_);
  or _51650_ (_00024_, _43565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _51651_ (_00025_, _00024_, _43569_);
  and _51652_ (_00026_, _00025_, _00023_);
  and _51653_ (_40778_, _43689_, _43634_);
  and _51654_ (_00027_, _40778_, _43568_);
  or _51655_ (_05088_, _00027_, _00026_);
  or _51656_ (_00028_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _51657_ (_00029_, \oc8051_gm_cxrom_1.cell0.valid );
  or _51658_ (_00030_, _00029_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _51659_ (_00031_, _00030_, _00028_);
  nand _51660_ (_00032_, _00031_, _43634_);
  or _51661_ (_00033_, \oc8051_gm_cxrom_1.cell0.data [7], _43634_);
  and _51662_ (_05096_, _00033_, _00032_);
  or _51663_ (_00034_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _51664_ (_00035_, \oc8051_gm_cxrom_1.cell0.data [0], _00029_);
  nand _51665_ (_00036_, _00035_, _00034_);
  nand _51666_ (_00037_, _00036_, _43634_);
  or _51667_ (_00038_, \oc8051_gm_cxrom_1.cell0.data [0], _43634_);
  and _51668_ (_05103_, _00038_, _00037_);
  or _51669_ (_00039_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _51670_ (_00040_, \oc8051_gm_cxrom_1.cell0.data [1], _00029_);
  nand _51671_ (_00041_, _00040_, _00039_);
  nand _51672_ (_00042_, _00041_, _43634_);
  or _51673_ (_00043_, \oc8051_gm_cxrom_1.cell0.data [1], _43634_);
  and _51674_ (_05107_, _00043_, _00042_);
  or _51675_ (_00044_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _51676_ (_00045_, \oc8051_gm_cxrom_1.cell0.data [2], _00029_);
  nand _51677_ (_00046_, _00045_, _00044_);
  nand _51678_ (_00047_, _00046_, _43634_);
  or _51679_ (_00048_, \oc8051_gm_cxrom_1.cell0.data [2], _43634_);
  and _51680_ (_05111_, _00048_, _00047_);
  or _51681_ (_00049_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _51682_ (_00050_, \oc8051_gm_cxrom_1.cell0.data [3], _00029_);
  nand _51683_ (_00051_, _00050_, _00049_);
  nand _51684_ (_00052_, _00051_, _43634_);
  or _51685_ (_00053_, \oc8051_gm_cxrom_1.cell0.data [3], _43634_);
  and _51686_ (_05115_, _00053_, _00052_);
  or _51687_ (_00054_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _51688_ (_00055_, \oc8051_gm_cxrom_1.cell0.data [4], _00029_);
  nand _51689_ (_00056_, _00055_, _00054_);
  nand _51690_ (_00057_, _00056_, _43634_);
  or _51691_ (_00058_, \oc8051_gm_cxrom_1.cell0.data [4], _43634_);
  and _51692_ (_05118_, _00058_, _00057_);
  nor _51693_ (_00059_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  nor _51694_ (_00060_, \oc8051_gm_cxrom_1.cell0.data [5], _00029_);
  or _51695_ (_00061_, _00060_, _00059_);
  nand _51696_ (_00062_, _00061_, _43634_);
  or _51697_ (_00063_, \oc8051_gm_cxrom_1.cell0.data [5], _43634_);
  and _51698_ (_05122_, _00063_, _00062_);
  or _51699_ (_00064_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _51700_ (_00065_, \oc8051_gm_cxrom_1.cell0.data [6], _00029_);
  nand _51701_ (_00066_, _00065_, _00064_);
  nand _51702_ (_00067_, _00066_, _43634_);
  or _51703_ (_00068_, \oc8051_gm_cxrom_1.cell0.data [6], _43634_);
  and _51704_ (_05126_, _00068_, _00067_);
  or _51705_ (_00069_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _51706_ (_00070_, \oc8051_gm_cxrom_1.cell1.valid );
  or _51707_ (_00071_, _00070_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _51708_ (_00072_, _00071_, _00069_);
  nand _51709_ (_00073_, _00072_, _43634_);
  or _51710_ (_00074_, \oc8051_gm_cxrom_1.cell1.data [7], _43634_);
  and _51711_ (_05148_, _00074_, _00073_);
  or _51712_ (_00075_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _51713_ (_00076_, \oc8051_gm_cxrom_1.cell1.data [0], _00070_);
  nand _51714_ (_00077_, _00076_, _00075_);
  nand _51715_ (_00078_, _00077_, _43634_);
  or _51716_ (_00079_, \oc8051_gm_cxrom_1.cell1.data [0], _43634_);
  and _51717_ (_05154_, _00079_, _00078_);
  or _51718_ (_00080_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _51719_ (_00081_, \oc8051_gm_cxrom_1.cell1.data [1], _00070_);
  nand _51720_ (_00082_, _00081_, _00080_);
  nand _51721_ (_00083_, _00082_, _43634_);
  or _51722_ (_00084_, \oc8051_gm_cxrom_1.cell1.data [1], _43634_);
  and _51723_ (_05158_, _00084_, _00083_);
  or _51724_ (_00085_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _51725_ (_00086_, \oc8051_gm_cxrom_1.cell1.data [2], _00070_);
  nand _51726_ (_00087_, _00086_, _00085_);
  nand _51727_ (_00088_, _00087_, _43634_);
  or _51728_ (_00089_, \oc8051_gm_cxrom_1.cell1.data [2], _43634_);
  and _51729_ (_05162_, _00089_, _00088_);
  or _51730_ (_00090_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _51731_ (_00091_, \oc8051_gm_cxrom_1.cell1.data [3], _00070_);
  nand _51732_ (_00092_, _00091_, _00090_);
  nand _51733_ (_00093_, _00092_, _43634_);
  or _51734_ (_00094_, \oc8051_gm_cxrom_1.cell1.data [3], _43634_);
  and _51735_ (_05166_, _00094_, _00093_);
  or _51736_ (_00095_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _51737_ (_00096_, \oc8051_gm_cxrom_1.cell1.data [4], _00070_);
  nand _51738_ (_00097_, _00096_, _00095_);
  nand _51739_ (_00098_, _00097_, _43634_);
  or _51740_ (_00099_, \oc8051_gm_cxrom_1.cell1.data [4], _43634_);
  and _51741_ (_05170_, _00099_, _00098_);
  nor _51742_ (_00100_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  nor _51743_ (_00101_, \oc8051_gm_cxrom_1.cell1.data [5], _00070_);
  or _51744_ (_00102_, _00101_, _00100_);
  nand _51745_ (_00103_, _00102_, _43634_);
  or _51746_ (_00104_, \oc8051_gm_cxrom_1.cell1.data [5], _43634_);
  and _51747_ (_05174_, _00104_, _00103_);
  or _51748_ (_00105_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _51749_ (_00106_, \oc8051_gm_cxrom_1.cell1.data [6], _00070_);
  nand _51750_ (_00107_, _00106_, _00105_);
  nand _51751_ (_00108_, _00107_, _43634_);
  or _51752_ (_00109_, \oc8051_gm_cxrom_1.cell1.data [6], _43634_);
  and _51753_ (_05178_, _00109_, _00108_);
  or _51754_ (_00110_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _51755_ (_00111_, \oc8051_gm_cxrom_1.cell2.valid );
  or _51756_ (_00112_, _00111_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _51757_ (_00113_, _00112_, _00110_);
  nand _51758_ (_00114_, _00113_, _43634_);
  or _51759_ (_00115_, \oc8051_gm_cxrom_1.cell2.data [7], _43634_);
  and _51760_ (_05199_, _00115_, _00114_);
  or _51761_ (_00116_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _51762_ (_00117_, \oc8051_gm_cxrom_1.cell2.data [0], _00111_);
  nand _51763_ (_00118_, _00117_, _00116_);
  nand _51764_ (_00119_, _00118_, _43634_);
  or _51765_ (_00120_, \oc8051_gm_cxrom_1.cell2.data [0], _43634_);
  and _51766_ (_05206_, _00120_, _00119_);
  or _51767_ (_00121_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _51768_ (_00122_, \oc8051_gm_cxrom_1.cell2.data [1], _00111_);
  nand _51769_ (_00123_, _00122_, _00121_);
  nand _51770_ (_00124_, _00123_, _43634_);
  or _51771_ (_00125_, \oc8051_gm_cxrom_1.cell2.data [1], _43634_);
  and _51772_ (_05210_, _00125_, _00124_);
  or _51773_ (_00126_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _51774_ (_00127_, \oc8051_gm_cxrom_1.cell2.data [2], _00111_);
  nand _51775_ (_00128_, _00127_, _00126_);
  nand _51776_ (_00129_, _00128_, _43634_);
  or _51777_ (_00130_, \oc8051_gm_cxrom_1.cell2.data [2], _43634_);
  and _51778_ (_05214_, _00130_, _00129_);
  or _51779_ (_00131_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _51780_ (_00132_, \oc8051_gm_cxrom_1.cell2.data [3], _00111_);
  nand _51781_ (_00133_, _00132_, _00131_);
  nand _51782_ (_00134_, _00133_, _43634_);
  or _51783_ (_00135_, \oc8051_gm_cxrom_1.cell2.data [3], _43634_);
  and _51784_ (_05218_, _00135_, _00134_);
  or _51785_ (_00136_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _51786_ (_00138_, \oc8051_gm_cxrom_1.cell2.data [4], _00111_);
  nand _51787_ (_00140_, _00138_, _00136_);
  nand _51788_ (_00142_, _00140_, _43634_);
  or _51789_ (_00144_, \oc8051_gm_cxrom_1.cell2.data [4], _43634_);
  and _51790_ (_05222_, _00144_, _00142_);
  nor _51791_ (_00147_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  nor _51792_ (_00149_, \oc8051_gm_cxrom_1.cell2.data [5], _00111_);
  or _51793_ (_00151_, _00149_, _00147_);
  nand _51794_ (_00153_, _00151_, _43634_);
  or _51795_ (_00155_, \oc8051_gm_cxrom_1.cell2.data [5], _43634_);
  and _51796_ (_05225_, _00155_, _00153_);
  or _51797_ (_00158_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _51798_ (_00160_, \oc8051_gm_cxrom_1.cell2.data [6], _00111_);
  nand _51799_ (_00162_, _00160_, _00158_);
  nand _51800_ (_00164_, _00162_, _43634_);
  or _51801_ (_00166_, \oc8051_gm_cxrom_1.cell2.data [6], _43634_);
  and _51802_ (_05229_, _00166_, _00164_);
  or _51803_ (_00169_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _51804_ (_00171_, \oc8051_gm_cxrom_1.cell3.valid );
  or _51805_ (_00173_, _00171_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _51806_ (_00175_, _00173_, _00169_);
  nand _51807_ (_00177_, _00175_, _43634_);
  or _51808_ (_00179_, \oc8051_gm_cxrom_1.cell3.data [7], _43634_);
  and _51809_ (_05251_, _00179_, _00177_);
  or _51810_ (_00182_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _51811_ (_00184_, \oc8051_gm_cxrom_1.cell3.data [0], _00171_);
  nand _51812_ (_00186_, _00184_, _00182_);
  nand _51813_ (_00188_, _00186_, _43634_);
  or _51814_ (_00190_, \oc8051_gm_cxrom_1.cell3.data [0], _43634_);
  and _51815_ (_05258_, _00190_, _00188_);
  or _51816_ (_00193_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _51817_ (_00194_, \oc8051_gm_cxrom_1.cell3.data [1], _00171_);
  nand _51818_ (_00195_, _00194_, _00193_);
  nand _51819_ (_00196_, _00195_, _43634_);
  or _51820_ (_00197_, \oc8051_gm_cxrom_1.cell3.data [1], _43634_);
  and _51821_ (_05261_, _00197_, _00196_);
  or _51822_ (_00198_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _51823_ (_00199_, \oc8051_gm_cxrom_1.cell3.data [2], _00171_);
  nand _51824_ (_00200_, _00199_, _00198_);
  nand _51825_ (_00201_, _00200_, _43634_);
  or _51826_ (_00202_, \oc8051_gm_cxrom_1.cell3.data [2], _43634_);
  and _51827_ (_05265_, _00202_, _00201_);
  or _51828_ (_00203_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _51829_ (_00204_, \oc8051_gm_cxrom_1.cell3.data [3], _00171_);
  nand _51830_ (_00205_, _00204_, _00203_);
  nand _51831_ (_00206_, _00205_, _43634_);
  or _51832_ (_00207_, \oc8051_gm_cxrom_1.cell3.data [3], _43634_);
  and _51833_ (_05269_, _00207_, _00206_);
  or _51834_ (_00208_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _51835_ (_00209_, \oc8051_gm_cxrom_1.cell3.data [4], _00171_);
  nand _51836_ (_00210_, _00209_, _00208_);
  nand _51837_ (_00211_, _00210_, _43634_);
  or _51838_ (_00212_, \oc8051_gm_cxrom_1.cell3.data [4], _43634_);
  and _51839_ (_05273_, _00212_, _00211_);
  nor _51840_ (_00213_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  nor _51841_ (_00214_, \oc8051_gm_cxrom_1.cell3.data [5], _00171_);
  or _51842_ (_00215_, _00214_, _00213_);
  nand _51843_ (_00216_, _00215_, _43634_);
  or _51844_ (_00217_, \oc8051_gm_cxrom_1.cell3.data [5], _43634_);
  and _51845_ (_05277_, _00217_, _00216_);
  or _51846_ (_00218_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _51847_ (_00219_, \oc8051_gm_cxrom_1.cell3.data [6], _00171_);
  nand _51848_ (_00220_, _00219_, _00218_);
  nand _51849_ (_00221_, _00220_, _43634_);
  or _51850_ (_00222_, \oc8051_gm_cxrom_1.cell3.data [6], _43634_);
  and _51851_ (_05281_, _00222_, _00221_);
  or _51852_ (_00223_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _51853_ (_00224_, \oc8051_gm_cxrom_1.cell4.valid );
  or _51854_ (_00225_, _00224_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _51855_ (_00226_, _00225_, _00223_);
  nand _51856_ (_00227_, _00226_, _43634_);
  or _51857_ (_00228_, \oc8051_gm_cxrom_1.cell4.data [7], _43634_);
  and _51858_ (_05302_, _00228_, _00227_);
  or _51859_ (_00229_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _51860_ (_00230_, \oc8051_gm_cxrom_1.cell4.data [0], _00224_);
  nand _51861_ (_00231_, _00230_, _00229_);
  nand _51862_ (_00232_, _00231_, _43634_);
  or _51863_ (_00233_, \oc8051_gm_cxrom_1.cell4.data [0], _43634_);
  and _51864_ (_05309_, _00233_, _00232_);
  or _51865_ (_00234_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _51866_ (_00235_, \oc8051_gm_cxrom_1.cell4.data [1], _00224_);
  nand _51867_ (_00236_, _00235_, _00234_);
  nand _51868_ (_00237_, _00236_, _43634_);
  or _51869_ (_00238_, \oc8051_gm_cxrom_1.cell4.data [1], _43634_);
  and _51870_ (_05313_, _00238_, _00237_);
  or _51871_ (_00239_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _51872_ (_00240_, \oc8051_gm_cxrom_1.cell4.data [2], _00224_);
  nand _51873_ (_00241_, _00240_, _00239_);
  nand _51874_ (_00242_, _00241_, _43634_);
  or _51875_ (_00243_, \oc8051_gm_cxrom_1.cell4.data [2], _43634_);
  and _51876_ (_05317_, _00243_, _00242_);
  or _51877_ (_00244_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _51878_ (_00245_, \oc8051_gm_cxrom_1.cell4.data [3], _00224_);
  nand _51879_ (_00246_, _00245_, _00244_);
  nand _51880_ (_00247_, _00246_, _43634_);
  or _51881_ (_00248_, \oc8051_gm_cxrom_1.cell4.data [3], _43634_);
  and _51882_ (_05321_, _00248_, _00247_);
  or _51883_ (_00249_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _51884_ (_00250_, \oc8051_gm_cxrom_1.cell4.data [4], _00224_);
  nand _51885_ (_00251_, _00250_, _00249_);
  nand _51886_ (_00252_, _00251_, _43634_);
  or _51887_ (_00253_, \oc8051_gm_cxrom_1.cell4.data [4], _43634_);
  and _51888_ (_05325_, _00253_, _00252_);
  nor _51889_ (_00254_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  nor _51890_ (_00255_, \oc8051_gm_cxrom_1.cell4.data [5], _00224_);
  or _51891_ (_00256_, _00255_, _00254_);
  nand _51892_ (_00257_, _00256_, _43634_);
  or _51893_ (_00258_, \oc8051_gm_cxrom_1.cell4.data [5], _43634_);
  and _51894_ (_05329_, _00258_, _00257_);
  or _51895_ (_00259_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _51896_ (_00260_, \oc8051_gm_cxrom_1.cell4.data [6], _00224_);
  nand _51897_ (_00261_, _00260_, _00259_);
  nand _51898_ (_00262_, _00261_, _43634_);
  or _51899_ (_00263_, \oc8051_gm_cxrom_1.cell4.data [6], _43634_);
  and _51900_ (_05333_, _00263_, _00262_);
  or _51901_ (_00264_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _51902_ (_00265_, \oc8051_gm_cxrom_1.cell5.valid );
  or _51903_ (_00266_, _00265_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _51904_ (_00267_, _00266_, _00264_);
  nand _51905_ (_00268_, _00267_, _43634_);
  or _51906_ (_00269_, \oc8051_gm_cxrom_1.cell5.data [7], _43634_);
  and _51907_ (_05354_, _00269_, _00268_);
  or _51908_ (_00270_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _51909_ (_00271_, \oc8051_gm_cxrom_1.cell5.data [0], _00265_);
  nand _51910_ (_00272_, _00271_, _00270_);
  nand _51911_ (_00273_, _00272_, _43634_);
  or _51912_ (_00274_, \oc8051_gm_cxrom_1.cell5.data [0], _43634_);
  and _51913_ (_05361_, _00274_, _00273_);
  or _51914_ (_00275_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _51915_ (_00276_, \oc8051_gm_cxrom_1.cell5.data [1], _00265_);
  nand _51916_ (_00277_, _00276_, _00275_);
  nand _51917_ (_00278_, _00277_, _43634_);
  or _51918_ (_00279_, \oc8051_gm_cxrom_1.cell5.data [1], _43634_);
  and _51919_ (_05365_, _00279_, _00278_);
  or _51920_ (_00280_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _51921_ (_00281_, \oc8051_gm_cxrom_1.cell5.data [2], _00265_);
  nand _51922_ (_00282_, _00281_, _00280_);
  nand _51923_ (_00283_, _00282_, _43634_);
  or _51924_ (_00284_, \oc8051_gm_cxrom_1.cell5.data [2], _43634_);
  and _51925_ (_05369_, _00284_, _00283_);
  or _51926_ (_00285_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _51927_ (_00286_, \oc8051_gm_cxrom_1.cell5.data [3], _00265_);
  nand _51928_ (_00287_, _00286_, _00285_);
  nand _51929_ (_00288_, _00287_, _43634_);
  or _51930_ (_00289_, \oc8051_gm_cxrom_1.cell5.data [3], _43634_);
  and _51931_ (_05372_, _00289_, _00288_);
  or _51932_ (_00290_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _51933_ (_00291_, \oc8051_gm_cxrom_1.cell5.data [4], _00265_);
  nand _51934_ (_00292_, _00291_, _00290_);
  nand _51935_ (_00293_, _00292_, _43634_);
  or _51936_ (_00294_, \oc8051_gm_cxrom_1.cell5.data [4], _43634_);
  and _51937_ (_05376_, _00294_, _00293_);
  nor _51938_ (_00295_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  nor _51939_ (_00296_, \oc8051_gm_cxrom_1.cell5.data [5], _00265_);
  or _51940_ (_00297_, _00296_, _00295_);
  nand _51941_ (_00298_, _00297_, _43634_);
  or _51942_ (_00299_, \oc8051_gm_cxrom_1.cell5.data [5], _43634_);
  and _51943_ (_05380_, _00299_, _00298_);
  or _51944_ (_00300_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _51945_ (_00301_, \oc8051_gm_cxrom_1.cell5.data [6], _00265_);
  nand _51946_ (_00302_, _00301_, _00300_);
  nand _51947_ (_00303_, _00302_, _43634_);
  or _51948_ (_00304_, \oc8051_gm_cxrom_1.cell5.data [6], _43634_);
  and _51949_ (_05384_, _00304_, _00303_);
  or _51950_ (_00305_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _51951_ (_00306_, \oc8051_gm_cxrom_1.cell6.valid );
  or _51952_ (_00307_, _00306_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _51953_ (_00308_, _00307_, _00305_);
  nand _51954_ (_00309_, _00308_, _43634_);
  or _51955_ (_00310_, \oc8051_gm_cxrom_1.cell6.data [7], _43634_);
  and _51956_ (_05405_, _00310_, _00309_);
  or _51957_ (_00311_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _51958_ (_00312_, \oc8051_gm_cxrom_1.cell6.data [0], _00306_);
  nand _51959_ (_00313_, _00312_, _00311_);
  nand _51960_ (_00314_, _00313_, _43634_);
  or _51961_ (_00315_, \oc8051_gm_cxrom_1.cell6.data [0], _43634_);
  and _51962_ (_05412_, _00315_, _00314_);
  or _51963_ (_00316_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _51964_ (_00317_, \oc8051_gm_cxrom_1.cell6.data [1], _00306_);
  nand _51965_ (_00318_, _00317_, _00316_);
  nand _51966_ (_00319_, _00318_, _43634_);
  or _51967_ (_00320_, \oc8051_gm_cxrom_1.cell6.data [1], _43634_);
  and _51968_ (_05416_, _00320_, _00319_);
  or _51969_ (_00321_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _51970_ (_00322_, \oc8051_gm_cxrom_1.cell6.data [2], _00306_);
  nand _51971_ (_00323_, _00322_, _00321_);
  nand _51972_ (_00324_, _00323_, _43634_);
  or _51973_ (_00325_, \oc8051_gm_cxrom_1.cell6.data [2], _43634_);
  and _51974_ (_05420_, _00325_, _00324_);
  or _51975_ (_00326_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _51976_ (_00327_, \oc8051_gm_cxrom_1.cell6.data [3], _00306_);
  nand _51977_ (_00328_, _00327_, _00326_);
  nand _51978_ (_00329_, _00328_, _43634_);
  or _51979_ (_00330_, \oc8051_gm_cxrom_1.cell6.data [3], _43634_);
  and _51980_ (_05424_, _00330_, _00329_);
  or _51981_ (_00331_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _51982_ (_00332_, \oc8051_gm_cxrom_1.cell6.data [4], _00306_);
  nand _51983_ (_00333_, _00332_, _00331_);
  nand _51984_ (_00334_, _00333_, _43634_);
  or _51985_ (_00335_, \oc8051_gm_cxrom_1.cell6.data [4], _43634_);
  and _51986_ (_05428_, _00335_, _00334_);
  nor _51987_ (_00336_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  nor _51988_ (_00337_, \oc8051_gm_cxrom_1.cell6.data [5], _00306_);
  or _51989_ (_00338_, _00337_, _00336_);
  nand _51990_ (_00339_, _00338_, _43634_);
  or _51991_ (_00340_, \oc8051_gm_cxrom_1.cell6.data [5], _43634_);
  and _51992_ (_05432_, _00340_, _00339_);
  or _51993_ (_00341_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _51994_ (_00342_, \oc8051_gm_cxrom_1.cell6.data [6], _00306_);
  nand _51995_ (_00343_, _00342_, _00341_);
  nand _51996_ (_00344_, _00343_, _43634_);
  or _51997_ (_00345_, \oc8051_gm_cxrom_1.cell6.data [6], _43634_);
  and _51998_ (_05436_, _00345_, _00344_);
  or _51999_ (_00346_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _52000_ (_00347_, \oc8051_gm_cxrom_1.cell7.valid );
  or _52001_ (_00348_, _00347_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _52002_ (_00349_, _00348_, _00346_);
  nand _52003_ (_00350_, _00349_, _43634_);
  or _52004_ (_00351_, \oc8051_gm_cxrom_1.cell7.data [7], _43634_);
  and _52005_ (_05457_, _00351_, _00350_);
  or _52006_ (_00352_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _52007_ (_00353_, \oc8051_gm_cxrom_1.cell7.data [0], _00347_);
  nand _52008_ (_00354_, _00353_, _00352_);
  nand _52009_ (_00355_, _00354_, _43634_);
  or _52010_ (_00356_, \oc8051_gm_cxrom_1.cell7.data [0], _43634_);
  and _52011_ (_05464_, _00356_, _00355_);
  or _52012_ (_00357_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _52013_ (_00358_, \oc8051_gm_cxrom_1.cell7.data [1], _00347_);
  nand _52014_ (_00359_, _00358_, _00357_);
  nand _52015_ (_00360_, _00359_, _43634_);
  or _52016_ (_00361_, \oc8051_gm_cxrom_1.cell7.data [1], _43634_);
  and _52017_ (_05468_, _00361_, _00360_);
  or _52018_ (_00362_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _52019_ (_00363_, \oc8051_gm_cxrom_1.cell7.data [2], _00347_);
  nand _52020_ (_00364_, _00363_, _00362_);
  nand _52021_ (_00365_, _00364_, _43634_);
  or _52022_ (_00366_, \oc8051_gm_cxrom_1.cell7.data [2], _43634_);
  and _52023_ (_05472_, _00366_, _00365_);
  or _52024_ (_00367_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _52025_ (_00368_, \oc8051_gm_cxrom_1.cell7.data [3], _00347_);
  nand _52026_ (_00369_, _00368_, _00367_);
  nand _52027_ (_00370_, _00369_, _43634_);
  or _52028_ (_00371_, \oc8051_gm_cxrom_1.cell7.data [3], _43634_);
  and _52029_ (_05476_, _00371_, _00370_);
  or _52030_ (_00372_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _52031_ (_00373_, \oc8051_gm_cxrom_1.cell7.data [4], _00347_);
  nand _52032_ (_00374_, _00373_, _00372_);
  nand _52033_ (_00375_, _00374_, _43634_);
  or _52034_ (_00376_, \oc8051_gm_cxrom_1.cell7.data [4], _43634_);
  and _52035_ (_05479_, _00376_, _00375_);
  nor _52036_ (_00377_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  nor _52037_ (_00378_, \oc8051_gm_cxrom_1.cell7.data [5], _00347_);
  or _52038_ (_00379_, _00378_, _00377_);
  nand _52039_ (_00380_, _00379_, _43634_);
  or _52040_ (_00381_, \oc8051_gm_cxrom_1.cell7.data [5], _43634_);
  and _52041_ (_05483_, _00381_, _00380_);
  or _52042_ (_00382_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _52043_ (_00383_, \oc8051_gm_cxrom_1.cell7.data [6], _00347_);
  nand _52044_ (_00384_, _00383_, _00382_);
  nand _52045_ (_00385_, _00384_, _43634_);
  or _52046_ (_00386_, \oc8051_gm_cxrom_1.cell7.data [6], _43634_);
  and _52047_ (_05487_, _00386_, _00385_);
  or _52048_ (_00387_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _52049_ (_00388_, \oc8051_gm_cxrom_1.cell8.valid );
  or _52050_ (_00389_, _00388_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _52051_ (_00390_, _00389_, _00387_);
  nand _52052_ (_00391_, _00390_, _43634_);
  or _52053_ (_00392_, \oc8051_gm_cxrom_1.cell8.data [7], _43634_);
  and _52054_ (_05509_, _00392_, _00391_);
  or _52055_ (_00393_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _52056_ (_00394_, \oc8051_gm_cxrom_1.cell8.data [0], _00388_);
  nand _52057_ (_00395_, _00394_, _00393_);
  nand _52058_ (_00396_, _00395_, _43634_);
  or _52059_ (_00397_, \oc8051_gm_cxrom_1.cell8.data [0], _43634_);
  and _52060_ (_05515_, _00397_, _00396_);
  or _52061_ (_00398_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _52062_ (_00399_, \oc8051_gm_cxrom_1.cell8.data [1], _00388_);
  nand _52063_ (_00400_, _00399_, _00398_);
  nand _52064_ (_00401_, _00400_, _43634_);
  or _52065_ (_00402_, \oc8051_gm_cxrom_1.cell8.data [1], _43634_);
  and _52066_ (_05519_, _00402_, _00401_);
  or _52067_ (_00403_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _52068_ (_00404_, \oc8051_gm_cxrom_1.cell8.data [2], _00388_);
  nand _52069_ (_00405_, _00404_, _00403_);
  nand _52070_ (_00406_, _00405_, _43634_);
  or _52071_ (_00407_, \oc8051_gm_cxrom_1.cell8.data [2], _43634_);
  and _52072_ (_05523_, _00407_, _00406_);
  or _52073_ (_00408_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _52074_ (_00409_, \oc8051_gm_cxrom_1.cell8.data [3], _00388_);
  nand _52075_ (_00410_, _00409_, _00408_);
  nand _52076_ (_00411_, _00410_, _43634_);
  or _52077_ (_00412_, \oc8051_gm_cxrom_1.cell8.data [3], _43634_);
  and _52078_ (_05527_, _00412_, _00411_);
  or _52079_ (_00413_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _52080_ (_00414_, \oc8051_gm_cxrom_1.cell8.data [4], _00388_);
  nand _52081_ (_00415_, _00414_, _00413_);
  nand _52082_ (_00416_, _00415_, _43634_);
  or _52083_ (_00417_, \oc8051_gm_cxrom_1.cell8.data [4], _43634_);
  and _52084_ (_05531_, _00417_, _00416_);
  nor _52085_ (_00418_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  nor _52086_ (_00419_, \oc8051_gm_cxrom_1.cell8.data [5], _00388_);
  or _52087_ (_00420_, _00419_, _00418_);
  nand _52088_ (_00421_, _00420_, _43634_);
  or _52089_ (_00422_, \oc8051_gm_cxrom_1.cell8.data [5], _43634_);
  and _52090_ (_05535_, _00422_, _00421_);
  or _52091_ (_00423_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _52092_ (_00424_, \oc8051_gm_cxrom_1.cell8.data [6], _00388_);
  nand _52093_ (_00425_, _00424_, _00423_);
  nand _52094_ (_00426_, _00425_, _43634_);
  or _52095_ (_00427_, \oc8051_gm_cxrom_1.cell8.data [6], _43634_);
  and _52096_ (_05539_, _00427_, _00426_);
  or _52097_ (_00428_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _52098_ (_00429_, \oc8051_gm_cxrom_1.cell9.valid );
  or _52099_ (_00430_, _00429_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _52100_ (_00431_, _00430_, _00428_);
  nand _52101_ (_00432_, _00431_, _43634_);
  or _52102_ (_00433_, \oc8051_gm_cxrom_1.cell9.data [7], _43634_);
  and _52103_ (_05560_, _00433_, _00432_);
  or _52104_ (_00434_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _52105_ (_00435_, \oc8051_gm_cxrom_1.cell9.data [0], _00429_);
  nand _52106_ (_00436_, _00435_, _00434_);
  nand _52107_ (_00437_, _00436_, _43634_);
  or _52108_ (_00438_, \oc8051_gm_cxrom_1.cell9.data [0], _43634_);
  and _52109_ (_05567_, _00438_, _00437_);
  or _52110_ (_00439_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _52111_ (_00440_, \oc8051_gm_cxrom_1.cell9.data [1], _00429_);
  nand _52112_ (_00441_, _00440_, _00439_);
  nand _52113_ (_00442_, _00441_, _43634_);
  or _52114_ (_00443_, \oc8051_gm_cxrom_1.cell9.data [1], _43634_);
  and _52115_ (_05571_, _00443_, _00442_);
  or _52116_ (_00444_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _52117_ (_00445_, \oc8051_gm_cxrom_1.cell9.data [2], _00429_);
  nand _52118_ (_00446_, _00445_, _00444_);
  nand _52119_ (_00447_, _00446_, _43634_);
  or _52120_ (_00448_, \oc8051_gm_cxrom_1.cell9.data [2], _43634_);
  and _52121_ (_05575_, _00448_, _00447_);
  or _52122_ (_00449_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _52123_ (_00450_, \oc8051_gm_cxrom_1.cell9.data [3], _00429_);
  nand _52124_ (_00451_, _00450_, _00449_);
  nand _52125_ (_00452_, _00451_, _43634_);
  or _52126_ (_00453_, \oc8051_gm_cxrom_1.cell9.data [3], _43634_);
  and _52127_ (_05579_, _00453_, _00452_);
  or _52128_ (_00454_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _52129_ (_00455_, \oc8051_gm_cxrom_1.cell9.data [4], _00429_);
  nand _52130_ (_00456_, _00455_, _00454_);
  nand _52131_ (_00457_, _00456_, _43634_);
  or _52132_ (_00458_, \oc8051_gm_cxrom_1.cell9.data [4], _43634_);
  and _52133_ (_05583_, _00458_, _00457_);
  nor _52134_ (_00459_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  nor _52135_ (_00460_, \oc8051_gm_cxrom_1.cell9.data [5], _00429_);
  or _52136_ (_00461_, _00460_, _00459_);
  nand _52137_ (_00462_, _00461_, _43634_);
  or _52138_ (_00463_, \oc8051_gm_cxrom_1.cell9.data [5], _43634_);
  and _52139_ (_05587_, _00463_, _00462_);
  or _52140_ (_00464_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _52141_ (_00465_, \oc8051_gm_cxrom_1.cell9.data [6], _00429_);
  nand _52142_ (_00466_, _00465_, _00464_);
  nand _52143_ (_00467_, _00466_, _43634_);
  or _52144_ (_00468_, \oc8051_gm_cxrom_1.cell9.data [6], _43634_);
  and _52145_ (_05590_, _00468_, _00467_);
  or _52146_ (_00469_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _52147_ (_00470_, \oc8051_gm_cxrom_1.cell10.valid );
  or _52148_ (_00471_, _00470_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _52149_ (_00472_, _00471_, _00469_);
  nand _52150_ (_00473_, _00472_, _43634_);
  or _52151_ (_00474_, \oc8051_gm_cxrom_1.cell10.data [7], _43634_);
  and _52152_ (_05612_, _00474_, _00473_);
  or _52153_ (_00475_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _52154_ (_00476_, \oc8051_gm_cxrom_1.cell10.data [0], _00470_);
  nand _52155_ (_00477_, _00476_, _00475_);
  nand _52156_ (_00478_, _00477_, _43634_);
  or _52157_ (_00479_, \oc8051_gm_cxrom_1.cell10.data [0], _43634_);
  and _52158_ (_05619_, _00479_, _00478_);
  or _52159_ (_00480_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _52160_ (_00481_, \oc8051_gm_cxrom_1.cell10.data [1], _00470_);
  nand _52161_ (_00482_, _00481_, _00480_);
  nand _52162_ (_00483_, _00482_, _43634_);
  or _52163_ (_00484_, \oc8051_gm_cxrom_1.cell10.data [1], _43634_);
  and _52164_ (_05623_, _00484_, _00483_);
  or _52165_ (_00485_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _52166_ (_00486_, \oc8051_gm_cxrom_1.cell10.data [2], _00470_);
  nand _52167_ (_00487_, _00486_, _00485_);
  nand _52168_ (_00488_, _00487_, _43634_);
  or _52169_ (_00489_, \oc8051_gm_cxrom_1.cell10.data [2], _43634_);
  and _52170_ (_05626_, _00489_, _00488_);
  or _52171_ (_00490_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _52172_ (_00491_, \oc8051_gm_cxrom_1.cell10.data [3], _00470_);
  nand _52173_ (_00492_, _00491_, _00490_);
  nand _52174_ (_00493_, _00492_, _43634_);
  or _52175_ (_00494_, \oc8051_gm_cxrom_1.cell10.data [3], _43634_);
  and _52176_ (_05630_, _00494_, _00493_);
  or _52177_ (_00495_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _52178_ (_00496_, \oc8051_gm_cxrom_1.cell10.data [4], _00470_);
  nand _52179_ (_00497_, _00496_, _00495_);
  nand _52180_ (_00498_, _00497_, _43634_);
  or _52181_ (_00499_, \oc8051_gm_cxrom_1.cell10.data [4], _43634_);
  and _52182_ (_05634_, _00499_, _00498_);
  nor _52183_ (_00500_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  nor _52184_ (_00501_, \oc8051_gm_cxrom_1.cell10.data [5], _00470_);
  or _52185_ (_00502_, _00501_, _00500_);
  nand _52186_ (_00503_, _00502_, _43634_);
  or _52187_ (_00504_, \oc8051_gm_cxrom_1.cell10.data [5], _43634_);
  and _52188_ (_05638_, _00504_, _00503_);
  or _52189_ (_00505_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _52190_ (_00506_, \oc8051_gm_cxrom_1.cell10.data [6], _00470_);
  nand _52191_ (_00507_, _00506_, _00505_);
  nand _52192_ (_00508_, _00507_, _43634_);
  or _52193_ (_00509_, \oc8051_gm_cxrom_1.cell10.data [6], _43634_);
  and _52194_ (_05642_, _00509_, _00508_);
  or _52195_ (_00510_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _52196_ (_00511_, \oc8051_gm_cxrom_1.cell11.valid );
  or _52197_ (_00512_, _00511_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _52198_ (_00513_, _00512_, _00510_);
  nand _52199_ (_00514_, _00513_, _43634_);
  or _52200_ (_00515_, \oc8051_gm_cxrom_1.cell11.data [7], _43634_);
  and _52201_ (_05663_, _00515_, _00514_);
  or _52202_ (_00516_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _52203_ (_00517_, \oc8051_gm_cxrom_1.cell11.data [0], _00511_);
  nand _52204_ (_00518_, _00517_, _00516_);
  nand _52205_ (_00519_, _00518_, _43634_);
  or _52206_ (_00520_, \oc8051_gm_cxrom_1.cell11.data [0], _43634_);
  and _52207_ (_05670_, _00520_, _00519_);
  or _52208_ (_00521_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _52209_ (_00522_, \oc8051_gm_cxrom_1.cell11.data [1], _00511_);
  nand _52210_ (_00523_, _00522_, _00521_);
  nand _52211_ (_00524_, _00523_, _43634_);
  or _52212_ (_00525_, \oc8051_gm_cxrom_1.cell11.data [1], _43634_);
  and _52213_ (_05674_, _00525_, _00524_);
  or _52214_ (_00526_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _52215_ (_00527_, \oc8051_gm_cxrom_1.cell11.data [2], _00511_);
  nand _52216_ (_00528_, _00527_, _00526_);
  nand _52217_ (_00529_, _00528_, _43634_);
  or _52218_ (_00530_, \oc8051_gm_cxrom_1.cell11.data [2], _43634_);
  and _52219_ (_05678_, _00530_, _00529_);
  or _52220_ (_00531_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _52221_ (_00532_, \oc8051_gm_cxrom_1.cell11.data [3], _00511_);
  nand _52222_ (_00533_, _00532_, _00531_);
  nand _52223_ (_00534_, _00533_, _43634_);
  or _52224_ (_00535_, \oc8051_gm_cxrom_1.cell11.data [3], _43634_);
  and _52225_ (_05682_, _00535_, _00534_);
  or _52226_ (_00536_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _52227_ (_00537_, \oc8051_gm_cxrom_1.cell11.data [4], _00511_);
  nand _52228_ (_00538_, _00537_, _00536_);
  nand _52229_ (_00539_, _00538_, _43634_);
  or _52230_ (_00540_, \oc8051_gm_cxrom_1.cell11.data [4], _43634_);
  and _52231_ (_05686_, _00540_, _00539_);
  nor _52232_ (_00541_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  nor _52233_ (_00542_, \oc8051_gm_cxrom_1.cell11.data [5], _00511_);
  or _52234_ (_00543_, _00542_, _00541_);
  nand _52235_ (_00544_, _00543_, _43634_);
  or _52236_ (_00545_, \oc8051_gm_cxrom_1.cell11.data [5], _43634_);
  and _52237_ (_05690_, _00545_, _00544_);
  or _52238_ (_00546_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _52239_ (_00547_, \oc8051_gm_cxrom_1.cell11.data [6], _00511_);
  nand _52240_ (_00548_, _00547_, _00546_);
  nand _52241_ (_00549_, _00548_, _43634_);
  or _52242_ (_00551_, \oc8051_gm_cxrom_1.cell11.data [6], _43634_);
  and _52243_ (_05694_, _00551_, _00549_);
  or _52244_ (_00553_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _52245_ (_00554_, \oc8051_gm_cxrom_1.cell12.valid );
  or _52246_ (_00556_, _00554_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _52247_ (_00557_, _00556_, _00553_);
  nand _52248_ (_00559_, _00557_, _43634_);
  or _52249_ (_00560_, \oc8051_gm_cxrom_1.cell12.data [7], _43634_);
  and _52250_ (_05716_, _00560_, _00559_);
  or _52251_ (_00562_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _52252_ (_00564_, \oc8051_gm_cxrom_1.cell12.data [0], _00554_);
  nand _52253_ (_00565_, _00564_, _00562_);
  nand _52254_ (_00567_, _00565_, _43634_);
  or _52255_ (_00568_, \oc8051_gm_cxrom_1.cell12.data [0], _43634_);
  and _52256_ (_05723_, _00568_, _00567_);
  or _52257_ (_00570_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _52258_ (_00572_, \oc8051_gm_cxrom_1.cell12.data [1], _00554_);
  nand _52259_ (_00573_, _00572_, _00570_);
  nand _52260_ (_00575_, _00573_, _43634_);
  or _52261_ (_00576_, \oc8051_gm_cxrom_1.cell12.data [1], _43634_);
  and _52262_ (_05727_, _00576_, _00575_);
  or _52263_ (_00578_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _52264_ (_00580_, \oc8051_gm_cxrom_1.cell12.data [2], _00554_);
  nand _52265_ (_00581_, _00580_, _00578_);
  nand _52266_ (_00583_, _00581_, _43634_);
  or _52267_ (_00584_, \oc8051_gm_cxrom_1.cell12.data [2], _43634_);
  and _52268_ (_05731_, _00584_, _00583_);
  or _52269_ (_00586_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _52270_ (_00588_, \oc8051_gm_cxrom_1.cell12.data [3], _00554_);
  nand _52271_ (_00589_, _00588_, _00586_);
  nand _52272_ (_00591_, _00589_, _43634_);
  or _52273_ (_00592_, \oc8051_gm_cxrom_1.cell12.data [3], _43634_);
  and _52274_ (_05735_, _00592_, _00591_);
  or _52275_ (_00594_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _52276_ (_00596_, \oc8051_gm_cxrom_1.cell12.data [4], _00554_);
  nand _52277_ (_00597_, _00596_, _00594_);
  nand _52278_ (_00599_, _00597_, _43634_);
  or _52279_ (_00600_, \oc8051_gm_cxrom_1.cell12.data [4], _43634_);
  and _52280_ (_05739_, _00600_, _00599_);
  nor _52281_ (_00601_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  nor _52282_ (_00602_, \oc8051_gm_cxrom_1.cell12.data [5], _00554_);
  or _52283_ (_00603_, _00602_, _00601_);
  nand _52284_ (_00604_, _00603_, _43634_);
  or _52285_ (_00605_, \oc8051_gm_cxrom_1.cell12.data [5], _43634_);
  and _52286_ (_05743_, _00605_, _00604_);
  or _52287_ (_00606_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _52288_ (_00607_, \oc8051_gm_cxrom_1.cell12.data [6], _00554_);
  nand _52289_ (_00608_, _00607_, _00606_);
  nand _52290_ (_00609_, _00608_, _43634_);
  or _52291_ (_00610_, \oc8051_gm_cxrom_1.cell12.data [6], _43634_);
  and _52292_ (_05747_, _00610_, _00609_);
  or _52293_ (_00611_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _52294_ (_00612_, \oc8051_gm_cxrom_1.cell13.valid );
  or _52295_ (_00613_, _00612_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _52296_ (_00614_, _00613_, _00611_);
  nand _52297_ (_00615_, _00614_, _43634_);
  or _52298_ (_00616_, \oc8051_gm_cxrom_1.cell13.data [7], _43634_);
  and _52299_ (_05769_, _00616_, _00615_);
  or _52300_ (_00617_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _52301_ (_00618_, \oc8051_gm_cxrom_1.cell13.data [0], _00612_);
  nand _52302_ (_00619_, _00618_, _00617_);
  nand _52303_ (_00620_, _00619_, _43634_);
  or _52304_ (_00621_, \oc8051_gm_cxrom_1.cell13.data [0], _43634_);
  and _52305_ (_05776_, _00621_, _00620_);
  or _52306_ (_00622_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _52307_ (_00623_, \oc8051_gm_cxrom_1.cell13.data [1], _00612_);
  nand _52308_ (_00624_, _00623_, _00622_);
  nand _52309_ (_00625_, _00624_, _43634_);
  or _52310_ (_00626_, \oc8051_gm_cxrom_1.cell13.data [1], _43634_);
  and _52311_ (_05780_, _00626_, _00625_);
  or _52312_ (_00627_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _52313_ (_00628_, \oc8051_gm_cxrom_1.cell13.data [2], _00612_);
  nand _52314_ (_00629_, _00628_, _00627_);
  nand _52315_ (_00630_, _00629_, _43634_);
  or _52316_ (_00631_, \oc8051_gm_cxrom_1.cell13.data [2], _43634_);
  and _52317_ (_05784_, _00631_, _00630_);
  or _52318_ (_00632_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _52319_ (_00633_, \oc8051_gm_cxrom_1.cell13.data [3], _00612_);
  nand _52320_ (_00634_, _00633_, _00632_);
  nand _52321_ (_00635_, _00634_, _43634_);
  or _52322_ (_00636_, \oc8051_gm_cxrom_1.cell13.data [3], _43634_);
  and _52323_ (_05788_, _00636_, _00635_);
  or _52324_ (_00637_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _52325_ (_00638_, \oc8051_gm_cxrom_1.cell13.data [4], _00612_);
  nand _52326_ (_00639_, _00638_, _00637_);
  nand _52327_ (_00640_, _00639_, _43634_);
  or _52328_ (_00641_, \oc8051_gm_cxrom_1.cell13.data [4], _43634_);
  and _52329_ (_05792_, _00641_, _00640_);
  nor _52330_ (_00642_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  nor _52331_ (_00643_, \oc8051_gm_cxrom_1.cell13.data [5], _00612_);
  or _52332_ (_00644_, _00643_, _00642_);
  nand _52333_ (_00645_, _00644_, _43634_);
  or _52334_ (_00646_, \oc8051_gm_cxrom_1.cell13.data [5], _43634_);
  and _52335_ (_05796_, _00646_, _00645_);
  or _52336_ (_00647_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _52337_ (_00648_, \oc8051_gm_cxrom_1.cell13.data [6], _00612_);
  nand _52338_ (_00649_, _00648_, _00647_);
  nand _52339_ (_00650_, _00649_, _43634_);
  or _52340_ (_00651_, \oc8051_gm_cxrom_1.cell13.data [6], _43634_);
  and _52341_ (_05800_, _00651_, _00650_);
  or _52342_ (_00652_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _52343_ (_00653_, \oc8051_gm_cxrom_1.cell14.valid );
  or _52344_ (_00654_, _00653_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _52345_ (_00655_, _00654_, _00652_);
  nand _52346_ (_00656_, _00655_, _43634_);
  or _52347_ (_00657_, \oc8051_gm_cxrom_1.cell14.data [7], _43634_);
  and _52348_ (_05822_, _00657_, _00656_);
  or _52349_ (_00658_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _52350_ (_00659_, \oc8051_gm_cxrom_1.cell14.data [0], _00653_);
  nand _52351_ (_00660_, _00659_, _00658_);
  nand _52352_ (_00661_, _00660_, _43634_);
  or _52353_ (_00662_, \oc8051_gm_cxrom_1.cell14.data [0], _43634_);
  and _52354_ (_05829_, _00662_, _00661_);
  or _52355_ (_00663_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _52356_ (_00664_, \oc8051_gm_cxrom_1.cell14.data [1], _00653_);
  nand _52357_ (_00665_, _00664_, _00663_);
  nand _52358_ (_00666_, _00665_, _43634_);
  or _52359_ (_00667_, \oc8051_gm_cxrom_1.cell14.data [1], _43634_);
  and _52360_ (_05833_, _00667_, _00666_);
  or _52361_ (_00668_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _52362_ (_00669_, \oc8051_gm_cxrom_1.cell14.data [2], _00653_);
  nand _52363_ (_00670_, _00669_, _00668_);
  nand _52364_ (_00671_, _00670_, _43634_);
  or _52365_ (_00672_, \oc8051_gm_cxrom_1.cell14.data [2], _43634_);
  and _52366_ (_05837_, _00672_, _00671_);
  or _52367_ (_00673_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _52368_ (_00674_, \oc8051_gm_cxrom_1.cell14.data [3], _00653_);
  nand _52369_ (_00675_, _00674_, _00673_);
  nand _52370_ (_00676_, _00675_, _43634_);
  or _52371_ (_00677_, \oc8051_gm_cxrom_1.cell14.data [3], _43634_);
  and _52372_ (_05841_, _00677_, _00676_);
  or _52373_ (_00678_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _52374_ (_00679_, \oc8051_gm_cxrom_1.cell14.data [4], _00653_);
  nand _52375_ (_00680_, _00679_, _00678_);
  nand _52376_ (_00681_, _00680_, _43634_);
  or _52377_ (_00682_, \oc8051_gm_cxrom_1.cell14.data [4], _43634_);
  and _52378_ (_05845_, _00682_, _00681_);
  nor _52379_ (_00683_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  nor _52380_ (_00684_, \oc8051_gm_cxrom_1.cell14.data [5], _00653_);
  or _52381_ (_00685_, _00684_, _00683_);
  nand _52382_ (_00686_, _00685_, _43634_);
  or _52383_ (_00687_, \oc8051_gm_cxrom_1.cell14.data [5], _43634_);
  and _52384_ (_05849_, _00687_, _00686_);
  or _52385_ (_00688_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _52386_ (_00689_, \oc8051_gm_cxrom_1.cell14.data [6], _00653_);
  nand _52387_ (_00690_, _00689_, _00688_);
  nand _52388_ (_00691_, _00690_, _43634_);
  or _52389_ (_00692_, \oc8051_gm_cxrom_1.cell14.data [6], _43634_);
  and _52390_ (_05853_, _00692_, _00691_);
  or _52391_ (_00693_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _52392_ (_00694_, \oc8051_gm_cxrom_1.cell15.valid );
  or _52393_ (_00695_, _00694_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand _52394_ (_00696_, _00695_, _00693_);
  nand _52395_ (_00697_, _00696_, _43634_);
  or _52396_ (_00698_, \oc8051_gm_cxrom_1.cell15.data [7], _43634_);
  and _52397_ (_05875_, _00698_, _00697_);
  or _52398_ (_00699_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _52399_ (_00700_, \oc8051_gm_cxrom_1.cell15.data [0], _00694_);
  nand _52400_ (_00701_, _00700_, _00699_);
  nand _52401_ (_00702_, _00701_, _43634_);
  or _52402_ (_00703_, \oc8051_gm_cxrom_1.cell15.data [0], _43634_);
  and _52403_ (_05882_, _00703_, _00702_);
  or _52404_ (_00704_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _52405_ (_00705_, \oc8051_gm_cxrom_1.cell15.data [1], _00694_);
  nand _52406_ (_00706_, _00705_, _00704_);
  nand _52407_ (_00707_, _00706_, _43634_);
  or _52408_ (_00708_, \oc8051_gm_cxrom_1.cell15.data [1], _43634_);
  and _52409_ (_05886_, _00708_, _00707_);
  or _52410_ (_00709_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _52411_ (_00710_, \oc8051_gm_cxrom_1.cell15.data [2], _00694_);
  nand _52412_ (_00711_, _00710_, _00709_);
  nand _52413_ (_00712_, _00711_, _43634_);
  or _52414_ (_00713_, \oc8051_gm_cxrom_1.cell15.data [2], _43634_);
  and _52415_ (_05890_, _00713_, _00712_);
  or _52416_ (_00714_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _52417_ (_00715_, \oc8051_gm_cxrom_1.cell15.data [3], _00694_);
  nand _52418_ (_00716_, _00715_, _00714_);
  nand _52419_ (_00717_, _00716_, _43634_);
  or _52420_ (_00718_, \oc8051_gm_cxrom_1.cell15.data [3], _43634_);
  and _52421_ (_05894_, _00718_, _00717_);
  or _52422_ (_00719_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _52423_ (_00720_, \oc8051_gm_cxrom_1.cell15.data [4], _00694_);
  nand _52424_ (_00721_, _00720_, _00719_);
  nand _52425_ (_00722_, _00721_, _43634_);
  or _52426_ (_00723_, \oc8051_gm_cxrom_1.cell15.data [4], _43634_);
  and _52427_ (_05898_, _00723_, _00722_);
  nor _52428_ (_00724_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  nor _52429_ (_00725_, \oc8051_gm_cxrom_1.cell15.data [5], _00694_);
  or _52430_ (_00726_, _00725_, _00724_);
  nand _52431_ (_00727_, _00726_, _43634_);
  or _52432_ (_00728_, \oc8051_gm_cxrom_1.cell15.data [5], _43634_);
  and _52433_ (_05902_, _00728_, _00727_);
  or _52434_ (_00729_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _52435_ (_00730_, \oc8051_gm_cxrom_1.cell15.data [6], _00694_);
  nand _52436_ (_00731_, _00730_, _00729_);
  nand _52437_ (_00732_, _00731_, _43634_);
  or _52438_ (_00733_, \oc8051_gm_cxrom_1.cell15.data [6], _43634_);
  and _52439_ (_05906_, _00733_, _00732_);
  nor _52440_ (_09681_, _39103_, rst);
  and _52441_ (_00734_, _37676_, _43634_);
  nand _52442_ (_00735_, _00734_, _39188_);
  nor _52443_ (_00736_, _39088_, _38854_);
  or _52444_ (_09684_, _00736_, _00735_);
  and _52445_ (_00737_, _39018_, _38994_);
  nor _52446_ (_00738_, _39064_, _39041_);
  and _52447_ (_00739_, _00738_, _00737_);
  not _52448_ (_00740_, _38058_);
  not _52449_ (_00741_, _38282_);
  not _52450_ (_00742_, _38788_);
  and _52451_ (_00743_, _00742_, _38535_);
  and _52452_ (_00744_, _00743_, _00741_);
  and _52453_ (_00745_, _00744_, _00740_);
  and _52454_ (_00746_, _00745_, _00739_);
  not _52455_ (_00747_, _39041_);
  and _52456_ (_00748_, _39064_, _00747_);
  not _52457_ (_00749_, _38994_);
  nor _52458_ (_00750_, _39018_, _00749_);
  and _52459_ (_00751_, _00750_, _00748_);
  not _52460_ (_00752_, _38535_);
  and _52461_ (_00753_, _38282_, _00742_);
  nor _52462_ (_00754_, _00753_, _00752_);
  not _52463_ (_00755_, _00754_);
  and _52464_ (_00756_, _00755_, _00751_);
  or _52465_ (_00757_, _00756_, _00746_);
  and _52466_ (_00758_, _38058_, _00741_);
  and _52467_ (_00759_, _38788_, _38535_);
  and _52468_ (_00760_, _00759_, _00758_);
  not _52469_ (_00761_, _39018_);
  and _52470_ (_00762_, _00738_, _00761_);
  and _52471_ (_00763_, _00762_, _00760_);
  and _52472_ (_00764_, _38282_, _38788_);
  and _52473_ (_00765_, _38058_, _38535_);
  and _52474_ (_00766_, _00765_, _00764_);
  and _52475_ (_00767_, _39064_, _39041_);
  and _52476_ (_00768_, _00767_, _39018_);
  and _52477_ (_00769_, _00768_, _00766_);
  or _52478_ (_00770_, _00769_, _00763_);
  or _52479_ (_00771_, _00770_, _00757_);
  and _52480_ (_00772_, _00739_, _00752_);
  nor _52481_ (_00773_, _39064_, _00747_);
  and _52482_ (_00774_, _00773_, _38994_);
  and _52483_ (_00775_, _00774_, _00760_);
  nor _52484_ (_00776_, _00775_, _00772_);
  and _52485_ (_00777_, _00773_, _00750_);
  and _52486_ (_00778_, _00764_, _38535_);
  and _52487_ (_00779_, _00778_, _00740_);
  and _52488_ (_00780_, _00779_, _00777_);
  and _52489_ (_00781_, _00751_, _00744_);
  nor _52490_ (_00782_, _00781_, _00780_);
  nand _52491_ (_00783_, _00782_, _00776_);
  and _52492_ (_00784_, _39018_, _00749_);
  and _52493_ (_00785_, _00784_, _00748_);
  and _52494_ (_00786_, _00785_, _00760_);
  and _52495_ (_00787_, _00758_, _00743_);
  and _52496_ (_00788_, _00787_, _00749_);
  and _52497_ (_00789_, _00788_, _00748_);
  or _52498_ (_00790_, _00789_, _00786_);
  or _52499_ (_00791_, _00790_, _00783_);
  or _52500_ (_00792_, _00791_, _00771_);
  nor _52501_ (_00793_, _39018_, _38994_);
  and _52502_ (_00794_, _00793_, _00773_);
  nor _52503_ (_00795_, _00794_, _00740_);
  and _52504_ (_00796_, _00759_, _00741_);
  not _52505_ (_00797_, _00796_);
  nor _52506_ (_00798_, _00797_, _00795_);
  not _52507_ (_00799_, _00798_);
  and _52508_ (_00800_, _00767_, _00750_);
  and _52509_ (_00801_, _00800_, _00760_);
  and _52510_ (_00802_, _00773_, _00784_);
  and _52511_ (_00803_, _00802_, _00760_);
  nor _52512_ (_00804_, _00803_, _00801_);
  and _52513_ (_00805_, _00804_, _00799_);
  and _52514_ (_00806_, _00748_, _39018_);
  and _52515_ (_00807_, _00806_, _00779_);
  and _52516_ (_00808_, _00767_, _00761_);
  and _52517_ (_00809_, _00808_, _00766_);
  or _52518_ (_00810_, _00809_, _00807_);
  and _52519_ (_00811_, _00778_, _00762_);
  and _52520_ (_00812_, _00811_, _00749_);
  or _52521_ (_00813_, _00812_, _00810_);
  and _52522_ (_00814_, _00811_, _38994_);
  or _52523_ (_00815_, _00793_, _00737_);
  and _52524_ (_00816_, _00767_, _00760_);
  and _52525_ (_00817_, _00816_, _00815_);
  or _52526_ (_00818_, _00817_, _00814_);
  nor _52527_ (_00819_, _00818_, _00813_);
  nand _52528_ (_00820_, _00819_, _00805_);
  or _52529_ (_00821_, _00820_, _00792_);
  and _52530_ (_00822_, _00821_, _37687_);
  not _52531_ (_00823_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _52532_ (_00824_, _37665_, _19459_);
  and _52533_ (_00825_, _00824_, _39089_);
  nor _52534_ (_00826_, _00825_, _00823_);
  or _52535_ (_00827_, _00826_, rst);
  or _52536_ (_09687_, _00827_, _00822_);
  nand _52537_ (_00828_, _39041_, _37611_);
  or _52538_ (_00829_, _37611_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _52539_ (_00830_, _00829_, _43634_);
  and _52540_ (_09690_, _00830_, _00828_);
  and _52541_ (_00831_, \oc8051_top_1.oc8051_sfr1.wait_data , _43634_);
  and _52542_ (_00832_, _00831_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _52543_ (_00833_, _39088_, _39086_);
  or _52544_ (_00834_, _00833_, _39124_);
  and _52545_ (_00835_, _39123_, _38865_);
  and _52546_ (_00836_, _39094_, _39088_);
  and _52547_ (_00837_, _38854_, _39112_);
  or _52548_ (_00838_, _00837_, _00836_);
  or _52549_ (_00839_, _00838_, _00835_);
  or _52550_ (_00840_, _00839_, _00834_);
  and _52551_ (_00841_, _39097_, _39189_);
  and _52552_ (_00842_, _39075_, _38865_);
  and _52553_ (_00843_, _00842_, _39000_);
  nor _52554_ (_00844_, _00843_, _00841_);
  nand _52555_ (_00845_, _00844_, _39182_);
  or _52556_ (_00846_, _00845_, _00840_);
  and _52557_ (_00847_, _00846_, _00734_);
  or _52558_ (_09693_, _00847_, _00832_);
  and _52559_ (_00848_, _39076_, _39088_);
  or _52560_ (_00849_, _00848_, _39072_);
  and _52561_ (_00850_, _39000_, _38590_);
  and _52562_ (_00851_, _00850_, _39111_);
  or _52563_ (_00852_, _00851_, _39209_);
  and _52564_ (_00853_, _39107_, _39096_);
  and _52565_ (_00854_, _00853_, _39123_);
  or _52566_ (_00855_, _00854_, _00852_);
  or _52567_ (_00856_, _00855_, _00849_);
  and _52568_ (_00857_, _00856_, _37676_);
  and _52569_ (_00858_, _39199_, _00823_);
  and _52570_ (_00859_, _39101_, _00858_);
  and _52571_ (_00860_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52572_ (_00861_, _00860_, _00859_);
  or _52573_ (_00862_, _00861_, _00857_);
  and _52574_ (_09696_, _00862_, _43634_);
  and _52575_ (_00863_, _00831_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _52576_ (_00864_, _38999_, _38590_);
  and _52577_ (_00865_, _00864_, _39070_);
  and _52578_ (_00866_, _39097_, _39162_);
  or _52579_ (_00867_, _39163_, _39113_);
  or _52580_ (_00868_, _00867_, _00866_);
  and _52581_ (_00869_, _00853_, _39133_);
  or _52582_ (_00870_, _00869_, _00868_);
  nor _52583_ (_00871_, _39162_, _39112_);
  nor _52584_ (_00872_, _00871_, _39095_);
  and _52585_ (_00873_, _00864_, _39132_);
  nor _52586_ (_00874_, _00873_, _00872_);
  not _52587_ (_00875_, _00874_);
  or _52588_ (_00876_, _00875_, _39216_);
  and _52589_ (_00877_, _39097_, _39076_);
  and _52590_ (_00878_, _39097_, _39125_);
  or _52591_ (_00879_, _00878_, _00877_);
  or _52592_ (_00880_, _00879_, _00849_);
  or _52593_ (_00881_, _00880_, _00876_);
  or _52594_ (_00882_, _00881_, _00870_);
  or _52595_ (_00883_, _00882_, _00865_);
  and _52596_ (_00884_, _00883_, _00734_);
  or _52597_ (_09699_, _00884_, _00863_);
  and _52598_ (_00885_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52599_ (_00886_, _39141_, _37676_);
  or _52600_ (_00887_, _00886_, _00885_);
  or _52601_ (_00888_, _00887_, _00859_);
  and _52602_ (_09702_, _00888_, _43634_);
  not _52603_ (_00889_, _39189_);
  nor _52604_ (_00890_, _00736_, _00889_);
  nor _52605_ (_00891_, _00890_, _00842_);
  not _52606_ (_00892_, _00891_);
  and _52607_ (_00893_, _00892_, _00858_);
  or _52608_ (_00894_, _00893_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52609_ (_00895_, _39133_, _39119_);
  and _52610_ (_00896_, _38843_, _39108_);
  and _52611_ (_00897_, _00896_, _38999_);
  or _52612_ (_00898_, _00897_, _00895_);
  and _52613_ (_00899_, _00898_, _39091_);
  or _52614_ (_00900_, _00899_, _37622_);
  and _52615_ (_00901_, _39094_, _38865_);
  or _52616_ (_00902_, _00898_, _00901_);
  and _52617_ (_00903_, _00902_, _00900_);
  or _52618_ (_00904_, _00903_, _00894_);
  or _52619_ (_00905_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _19459_);
  and _52620_ (_00906_, _00905_, _43634_);
  and _52621_ (_09705_, _00906_, _00904_);
  and _52622_ (_00907_, _00831_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _52623_ (_00908_, _00864_, _39111_);
  or _52624_ (_00909_, _00873_, _00908_);
  or _52625_ (_00910_, _39072_, _39113_);
  or _52626_ (_00911_, _00910_, _00909_);
  and _52627_ (_00912_, _39070_, _39119_);
  or _52628_ (_00913_, _00869_, _00837_);
  or _52629_ (_00914_, _00913_, _00912_);
  or _52630_ (_00915_, _00851_, _39168_);
  or _52631_ (_00916_, _39133_, _39123_);
  and _52632_ (_00917_, _00916_, _39184_);
  or _52633_ (_00918_, _00917_, _00915_);
  or _52634_ (_00919_, _00918_, _00914_);
  or _52635_ (_00920_, _00919_, _00911_);
  and _52636_ (_00921_, _00920_, _00734_);
  or _52637_ (_09708_, _00921_, _00907_);
  and _52638_ (_00922_, _00831_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or _52639_ (_00923_, _00854_, _39135_);
  and _52640_ (_00924_, _39131_, _38865_);
  and _52641_ (_00925_, _00853_, _39144_);
  or _52642_ (_00927_, _00925_, _00924_);
  nor _52643_ (_00928_, _00927_, _00923_);
  nand _52644_ (_00929_, _00928_, _00874_);
  nand _52645_ (_00930_, _39097_, _39116_);
  nand _52646_ (_00931_, _00930_, _39121_);
  and _52647_ (_00932_, _39211_, _39111_);
  or _52648_ (_00933_, _39226_, _39220_);
  or _52649_ (_00934_, _00933_, _00932_);
  or _52650_ (_00935_, _00934_, _00931_);
  or _52651_ (_00936_, _00935_, _00929_);
  and _52652_ (_00937_, _00850_, _39110_);
  and _52653_ (_00938_, _00850_, _39079_);
  or _52654_ (_00939_, _00938_, _00937_);
  nor _52655_ (_00940_, _39214_, _39145_);
  nand _52656_ (_00941_, _00940_, _39130_);
  or _52657_ (_00942_, _00941_, _00939_);
  or _52658_ (_00943_, _00942_, _00870_);
  or _52659_ (_00944_, _00943_, _00936_);
  and _52660_ (_00945_, _00944_, _00734_);
  or _52661_ (_09711_, _00945_, _00922_);
  and _52662_ (_00946_, _39184_, _39158_);
  and _52663_ (_00947_, _39076_, _38590_);
  or _52664_ (_00948_, _00947_, _00946_);
  and _52665_ (_00949_, _39184_, _39076_);
  and _52666_ (_00950_, _39158_, _38590_);
  and _52667_ (_00951_, _00853_, _39158_);
  or _52668_ (_00952_, _00951_, _00950_);
  or _52669_ (_00953_, _00952_, _00949_);
  or _52670_ (_00954_, _00953_, _00948_);
  and _52671_ (_00955_, _00853_, _39076_);
  or _52672_ (_00957_, _00955_, _39101_);
  or _52673_ (_00958_, _00957_, _00954_);
  and _52674_ (_00959_, _00958_, _00734_);
  nor _52675_ (_00960_, _39100_, _37622_);
  and _52676_ (_00961_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _52677_ (_00962_, _00961_, _00960_);
  and _52678_ (_00963_, _00962_, _43634_);
  or _52679_ (_09714_, _00963_, _00959_);
  or _52680_ (_00964_, _39170_, _39168_);
  not _52681_ (_00965_, _39146_);
  or _52682_ (_00966_, _00867_, _00965_);
  or _52683_ (_00967_, _00966_, _00964_);
  and _52684_ (_00968_, _39078_, _38999_);
  and _52685_ (_00969_, _00968_, _39109_);
  or _52686_ (_00970_, _00969_, _39134_);
  or _52687_ (_00971_, _00895_, _39117_);
  or _52688_ (_00972_, _00971_, _00970_);
  nand _52689_ (_00973_, _39142_, _39127_);
  or _52690_ (_00974_, _00973_, _00972_);
  or _52691_ (_00975_, _00974_, _00967_);
  and _52692_ (_00977_, _00968_, _39184_);
  or _52693_ (_00978_, _00977_, _39214_);
  or _52694_ (_00979_, _00978_, _39186_);
  and _52695_ (_00980_, _00864_, _39078_);
  or _52696_ (_00981_, _00980_, _39224_);
  or _52697_ (_00982_, _00852_, _39191_);
  or _52698_ (_00983_, _00982_, _00981_);
  or _52699_ (_00984_, _00983_, _00979_);
  and _52700_ (_00985_, _39094_, _38590_);
  or _52701_ (_00986_, _00897_, _39150_);
  or _52702_ (_00987_, _00986_, _00985_);
  or _52703_ (_00988_, _00987_, _00875_);
  or _52704_ (_00989_, _00988_, _00984_);
  or _52705_ (_00990_, _00989_, _00975_);
  and _52706_ (_00991_, _00990_, _37676_);
  and _52707_ (_00992_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52708_ (_00993_, _39091_, _39180_);
  or _52709_ (_00994_, _00899_, _00859_);
  or _52710_ (_00995_, _00994_, _00993_);
  or _52711_ (_00996_, _00995_, _00992_);
  or _52712_ (_00997_, _00996_, _00991_);
  and _52713_ (_09717_, _00997_, _43634_);
  and _52714_ (_09776_, _39235_, _43634_);
  nor _52715_ (_09778_, _39203_, rst);
  not _52716_ (_00998_, _00734_);
  or _52717_ (_09781_, _00891_, _00998_);
  and _52718_ (_00999_, _39188_, _39088_);
  nor _52719_ (_01000_, _00999_, _00842_);
  or _52720_ (_09784_, _01000_, _00998_);
  or _52721_ (_01001_, _00789_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _52722_ (_01002_, _01001_, _00810_);
  and _52723_ (_01003_, _01002_, _00825_);
  nor _52724_ (_01004_, _00824_, _39089_);
  or _52725_ (_01005_, _01004_, rst);
  or _52726_ (_09787_, _01005_, _01003_);
  nand _52727_ (_01006_, _38058_, _37611_);
  or _52728_ (_01007_, _37611_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _52729_ (_01008_, _01007_, _43634_);
  and _52730_ (_09790_, _01008_, _01006_);
  not _52731_ (_01009_, _37611_);
  or _52732_ (_01010_, _38282_, _01009_);
  or _52733_ (_01011_, _37611_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _52734_ (_01012_, _01011_, _43634_);
  and _52735_ (_09793_, _01012_, _01010_);
  nand _52736_ (_01013_, _38788_, _37611_);
  or _52737_ (_01014_, _37611_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _52738_ (_01015_, _01014_, _43634_);
  and _52739_ (_09796_, _01015_, _01013_);
  nand _52740_ (_01016_, _38535_, _37611_);
  or _52741_ (_01017_, _37611_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _52742_ (_01018_, _01017_, _43634_);
  and _52743_ (_09799_, _01018_, _01016_);
  or _52744_ (_01019_, _38994_, _01009_);
  or _52745_ (_01020_, _37611_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _52746_ (_01021_, _01020_, _43634_);
  and _52747_ (_09802_, _01021_, _01019_);
  nand _52748_ (_01022_, _39018_, _37611_);
  or _52749_ (_01023_, _37611_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _52750_ (_01024_, _01023_, _43634_);
  and _52751_ (_09805_, _01024_, _01022_);
  nand _52752_ (_01025_, _39064_, _37611_);
  or _52753_ (_01026_, _37611_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _52754_ (_01027_, _01026_, _43634_);
  and _52755_ (_09808_, _01027_, _01025_);
  and _52756_ (_01028_, _00853_, _39149_);
  and _52757_ (_01029_, _00850_, _39188_);
  and _52758_ (_01030_, _39097_, _39080_);
  or _52759_ (_01031_, _01030_, _01029_);
  or _52760_ (_01032_, _01031_, _01028_);
  and _52761_ (_01033_, _39188_, _38999_);
  and _52762_ (_01034_, _01033_, _39097_);
  or _52763_ (_01035_, _01034_, _00955_);
  or _52764_ (_01036_, _01035_, _00927_);
  or _52765_ (_01037_, _01036_, _01032_);
  or _52766_ (_01038_, _01037_, _39222_);
  and _52767_ (_01039_, _00853_, _39116_);
  or _52768_ (_01040_, _01039_, _00848_);
  or _52769_ (_01041_, _39132_, _39112_);
  and _52770_ (_01042_, _01041_, _39097_);
  or _52771_ (_01043_, _01042_, _01040_);
  and _52772_ (_01044_, _39211_, _39115_);
  nor _52773_ (_01045_, _00938_, _01044_);
  or _52774_ (_01046_, _39189_, _39158_);
  nand _52775_ (_01047_, _01046_, _00853_);
  nand _52776_ (_01048_, _01047_, _01045_);
  or _52777_ (_01049_, _01048_, _01043_);
  and _52778_ (_01050_, _00850_, _39115_);
  or _52779_ (_01051_, _01050_, _39072_);
  or _52780_ (_01052_, _39226_, _00949_);
  or _52781_ (_01053_, _01052_, _01051_);
  and _52782_ (_01054_, _00864_, _39115_);
  or _52783_ (_01055_, _01054_, _00950_);
  or _52784_ (_01056_, _01055_, _00948_);
  or _52785_ (_01057_, _01056_, _01053_);
  or _52786_ (_01058_, _01057_, _01049_);
  or _52787_ (_01059_, _01058_, _01038_);
  and _52788_ (_01060_, _01059_, _37676_);
  or _52789_ (_01061_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _19459_);
  and _52790_ (_01062_, _01061_, _00894_);
  or _52791_ (_01063_, _01062_, _01060_);
  and _52792_ (_09811_, _01063_, _43634_);
  and _52793_ (_01064_, _00831_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _52794_ (_01065_, _01040_, _00939_);
  or _52795_ (_01066_, _39144_, _39116_);
  nand _52796_ (_01067_, _01066_, _39119_);
  and _52797_ (_01068_, _39184_, _39125_);
  and _52798_ (_01069_, _39125_, _38590_);
  nor _52799_ (_01070_, _01069_, _01068_);
  nand _52800_ (_01071_, _01070_, _01067_);
  or _52801_ (_01072_, _01071_, _01065_);
  not _52802_ (_01073_, _39154_);
  nand _52803_ (_01074_, _39097_, _01073_);
  and _52804_ (_01075_, _01074_, _39169_);
  nand _52805_ (_01076_, _01075_, _00844_);
  not _52806_ (_01077_, _39144_);
  nand _52807_ (_01078_, _39159_, _01077_);
  and _52808_ (_01079_, _01078_, _39097_);
  or _52809_ (_01080_, _01079_, _00934_);
  or _52810_ (_01081_, _01080_, _01076_);
  or _52811_ (_01082_, _01081_, _01072_);
  and _52812_ (_01083_, _01082_, _00734_);
  or _52813_ (_34137_, _01083_, _01064_);
  or _52814_ (_01084_, _00987_, _39224_);
  or _52815_ (_01085_, _01084_, _00975_);
  and _52816_ (_01086_, _01085_, _37676_);
  and _52817_ (_01087_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52818_ (_01088_, _01087_, _00995_);
  or _52819_ (_01089_, _01088_, _01086_);
  and _52820_ (_34139_, _01089_, _43634_);
  and _52821_ (_01090_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52822_ (_01091_, _01090_, _00994_);
  and _52823_ (_01092_, _01091_, _43634_);
  and _52824_ (_01093_, _39132_, _39119_);
  nor _52825_ (_01094_, _01093_, _00896_);
  nor _52826_ (_01095_, _01094_, _39000_);
  and _52827_ (_01096_, _39143_, _39000_);
  or _52828_ (_01097_, _01096_, _39209_);
  or _52829_ (_01098_, _01097_, _00979_);
  or _52830_ (_01099_, _01098_, _01095_);
  and _52831_ (_01100_, _01099_, _00734_);
  or _52832_ (_34142_, _01100_, _01092_);
  and _52833_ (_01101_, _00853_, _39125_);
  or _52834_ (_01102_, _00955_, _00841_);
  or _52835_ (_01103_, _01102_, _01101_);
  and _52836_ (_01104_, _39097_, _39123_);
  or _52837_ (_01105_, _01034_, _39098_);
  or _52838_ (_01106_, _01105_, _01104_);
  or _52839_ (_01107_, _01106_, _01042_);
  or _52840_ (_01108_, _01107_, _01103_);
  or _52841_ (_01109_, _01055_, _00924_);
  or _52842_ (_01110_, _01066_, _39080_);
  and _52843_ (_01111_, _01110_, _39097_);
  or _52844_ (_01112_, _00947_, _39208_);
  or _52845_ (_01113_, _01112_, _01111_);
  or _52846_ (_01114_, _01113_, _01109_);
  and _52847_ (_01115_, _00951_, _39000_);
  or _52848_ (_01116_, _01115_, _39081_);
  or _52849_ (_01117_, _00980_, _00977_);
  or _52850_ (_01118_, _01117_, _00949_);
  and _52851_ (_01119_, _39149_, _39119_);
  and _52852_ (_01120_, _01033_, _39109_);
  or _52853_ (_01121_, _01120_, _01119_);
  or _52854_ (_01122_, _01121_, _01118_);
  or _52855_ (_01123_, _01122_, _01116_);
  or _52856_ (_01124_, _00842_, _39099_);
  and _52857_ (_01125_, _00951_, _38999_);
  or _52858_ (_01126_, _01125_, _01028_);
  or _52859_ (_01127_, _01126_, _01124_);
  or _52860_ (_01128_, _01127_, _01095_);
  or _52861_ (_01129_, _01128_, _01123_);
  or _52862_ (_01130_, _01129_, _01114_);
  or _52863_ (_01131_, _01130_, _01108_);
  and _52864_ (_01132_, _01131_, _37676_);
  and _52865_ (_01133_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52866_ (_01134_, _00893_, _00960_);
  or _52867_ (_01135_, _01134_, _01133_);
  or _52868_ (_01136_, _01135_, _01132_);
  and _52869_ (_34144_, _01136_, _43634_);
  nand _52870_ (_01137_, _39082_, _39161_);
  and _52871_ (_01138_, _39117_, _38124_);
  and _52872_ (_01139_, _39145_, _38124_);
  or _52873_ (_01140_, _01139_, _01138_);
  or _52874_ (_01141_, _01140_, _01137_);
  and _52875_ (_01142_, _00864_, _39188_);
  and _52876_ (_01143_, _01033_, _39184_);
  or _52877_ (_01144_, _01143_, _00848_);
  or _52878_ (_01145_, _01144_, _01142_);
  or _52879_ (_01146_, _00969_, _00949_);
  or _52880_ (_01147_, _39099_, _39150_);
  or _52881_ (_01148_, _01147_, _01146_);
  or _52882_ (_01149_, _01148_, _01145_);
  or _52883_ (_01150_, _01112_, _01109_);
  or _52884_ (_01151_, _01150_, _01149_);
  or _52885_ (_01152_, _01151_, _01141_);
  or _52886_ (_01153_, _01152_, _01108_);
  and _52887_ (_01154_, _01153_, _37676_);
  and _52888_ (_01155_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52889_ (_01156_, _01155_, _01134_);
  or _52890_ (_01157_, _01156_, _01154_);
  and _52891_ (_34146_, _01157_, _43634_);
  and _52892_ (_01158_, _00831_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _52893_ (_01159_, _00949_, _39140_);
  and _52894_ (_01160_, _00946_, _38999_);
  or _52895_ (_01161_, _01160_, _01125_);
  or _52896_ (_01162_, _01161_, _01159_);
  not _52897_ (_01163_, _43083_);
  or _52898_ (_01164_, _00917_, _01163_);
  or _52899_ (_01165_, _01164_, _01162_);
  nor _52900_ (_01166_, _39068_, _39074_);
  and _52901_ (_01167_, _00864_, _01166_);
  and _52902_ (_01168_, _01167_, _39047_);
  and _52903_ (_01169_, _39175_, _38865_);
  and _52904_ (_01170_, _39125_, _38865_);
  or _52905_ (_01171_, _01170_, _01169_);
  or _52906_ (_01172_, _01171_, _01168_);
  or _52907_ (_01173_, _01172_, _00911_);
  or _52908_ (_01174_, _01173_, _01165_);
  not _52909_ (_01175_, _43082_);
  or _52910_ (_01176_, _00955_, _01175_);
  and _52911_ (_01177_, _39132_, _38865_);
  and _52912_ (_01178_, _01177_, _38999_);
  and _52913_ (_01179_, _00837_, _38124_);
  or _52914_ (_01180_, _01179_, _01178_);
  or _52915_ (_01181_, _01180_, _01176_);
  and _52916_ (_01182_, _39097_, _39112_);
  or _52917_ (_01183_, _01182_, _00869_);
  or _52918_ (_01184_, _00947_, _00851_);
  or _52919_ (_01185_, _01184_, _00964_);
  or _52920_ (_01186_, _01185_, _01183_);
  or _52921_ (_01187_, _01186_, _01181_);
  or _52922_ (_01188_, _01187_, _01174_);
  and _52923_ (_01189_, _01188_, _00734_);
  or _52924_ (_34148_, _01189_, _01158_);
  and _52925_ (_01190_, _00831_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _52926_ (_01191_, _39220_, _39129_);
  or _52927_ (_01192_, _00854_, _00932_);
  or _52928_ (_01193_, _01192_, _01191_);
  or _52929_ (_01194_, _01193_, _00931_);
  or _52930_ (_01195_, _01194_, _01127_);
  or _52931_ (_01196_, _01182_, _01169_);
  or _52932_ (_01197_, _01178_, _01116_);
  or _52933_ (_01198_, _01197_, _01196_);
  or _52934_ (_01199_, _00937_, _37633_);
  or _52935_ (_01200_, _01199_, _39072_);
  or _52936_ (_01201_, _01200_, _39208_);
  or _52937_ (_01202_, _01055_, _39152_);
  or _52938_ (_01203_, _01202_, _01201_);
  or _52939_ (_01204_, _01203_, _01198_);
  or _52940_ (_01205_, _01204_, _01195_);
  or _52941_ (_01206_, _39099_, _37622_);
  nor _52942_ (_01207_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and _52943_ (_01208_, _01207_, _01206_);
  and _52944_ (_01209_, _01208_, _01205_);
  or _52945_ (_34150_, _01209_, _01190_);
  and _52946_ (_01210_, _00831_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or _52947_ (_01211_, _01028_, _39150_);
  nor _52948_ (_01212_, _01211_, _39148_);
  nor _52949_ (_01213_, _01103_, _00868_);
  nand _52950_ (_01214_, _01213_, _01212_);
  and _52951_ (_01215_, _39125_, _38854_);
  or _52952_ (_01216_, _01215_, _01034_);
  or _52953_ (_01217_, _01054_, _01044_);
  or _52954_ (_01219_, _01217_, _01184_);
  or _52955_ (_01221_, _01219_, _01216_);
  or _52956_ (_01223_, _01069_, _00854_);
  and _52957_ (_01225_, _39158_, _38865_);
  or _52958_ (_01227_, _01225_, _00869_);
  or _52959_ (_01229_, _01227_, _01223_);
  or _52960_ (_01231_, _39099_, _39128_);
  or _52961_ (_01233_, _01231_, _39213_);
  or _52962_ (_01235_, _01233_, _01229_);
  or _52963_ (_01237_, _01235_, _01221_);
  or _52964_ (_01239_, _01237_, _00876_);
  or _52965_ (_01241_, _01239_, _01214_);
  and _52966_ (_01243_, _01241_, _01208_);
  or _52967_ (_34152_, _01243_, _01210_);
  or _52968_ (_01246_, _01217_, _01216_);
  or _52969_ (_01248_, _01246_, _01211_);
  or _52970_ (_01250_, _39214_, _39209_);
  nor _52971_ (_01252_, _01250_, _01177_);
  nand _52972_ (_01254_, _01252_, _43082_);
  or _52973_ (_01256_, _01183_, _00915_);
  or _52974_ (_01258_, _01256_, _01254_);
  or _52975_ (_01260_, _00875_, _00868_);
  or _52976_ (_01262_, _01260_, _01258_);
  or _52977_ (_01264_, _01262_, _01248_);
  and _52978_ (_01266_, _01264_, _37676_);
  and _52979_ (_01268_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52980_ (_01270_, _39098_, _19459_);
  or _52981_ (_01272_, _01270_, _01268_);
  or _52982_ (_01274_, _01272_, _01266_);
  and _52983_ (_34154_, _01274_, _43634_);
  and _52984_ (_01277_, _00831_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor _52985_ (_01279_, _00835_, _39171_);
  nand _52986_ (_01281_, _01279_, _43083_);
  not _52987_ (_01283_, _38843_);
  or _52988_ (_01285_, _38865_, _01283_);
  and _52989_ (_01287_, _01285_, _39125_);
  or _52990_ (_01289_, _01287_, _01196_);
  or _52991_ (_01291_, _01289_, _01281_);
  or _52992_ (_01293_, _01291_, _00954_);
  or _52993_ (_01295_, _01293_, _01181_);
  and _52994_ (_01297_, _01295_, _00734_);
  or _52995_ (_34156_, _01297_, _01277_);
  nor _52996_ (_39695_, _39041_, rst);
  nor _52997_ (_39696_, _43238_, rst);
  and _52998_ (_01302_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _52999_ (_01304_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _53000_ (_01306_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _53001_ (_01308_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _53002_ (_01310_, _01308_, _01306_);
  and _53003_ (_01311_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _53004_ (_01312_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _53005_ (_01313_, _01312_, _01311_);
  and _53006_ (_01314_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _53007_ (_01315_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _53008_ (_01316_, _01315_, _01314_);
  and _53009_ (_01317_, _01316_, _01313_);
  and _53010_ (_01318_, _01317_, _01310_);
  nor _53011_ (_01319_, _01318_, _37742_);
  nor _53012_ (_01320_, _01319_, _01304_);
  nor _53013_ (_01321_, _01320_, _43140_);
  nor _53014_ (_01322_, _01321_, _01302_);
  nor _53015_ (_39698_, _01322_, rst);
  nor _53016_ (_39706_, _38058_, rst);
  and _53017_ (_39708_, _38282_, _43634_);
  nor _53018_ (_39709_, _38788_, rst);
  nor _53019_ (_39710_, _38535_, rst);
  and _53020_ (_39711_, _38994_, _43634_);
  nor _53021_ (_39712_, _39018_, rst);
  nor _53022_ (_39713_, _39064_, rst);
  nor _53023_ (_39714_, _43360_, rst);
  nor _53024_ (_39715_, _43276_, rst);
  nor _53025_ (_39717_, _43156_, rst);
  nor _53026_ (_39718_, _43399_, rst);
  nor _53027_ (_39719_, _43300_, rst);
  nor _53028_ (_39720_, _43184_, rst);
  nor _53029_ (_39721_, _43445_, rst);
  and _53030_ (_01323_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _53031_ (_01324_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _53032_ (_01325_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _53033_ (_01326_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _53034_ (_01327_, _01326_, _01325_);
  and _53035_ (_01328_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _53036_ (_01329_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _53037_ (_01330_, _01329_, _01328_);
  and _53038_ (_01331_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _53039_ (_01332_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _53040_ (_01333_, _01332_, _01331_);
  and _53041_ (_01334_, _01333_, _01330_);
  and _53042_ (_01335_, _01334_, _01327_);
  nor _53043_ (_01336_, _01335_, _37742_);
  nor _53044_ (_01337_, _01336_, _01324_);
  nor _53045_ (_01338_, _01337_, _43140_);
  nor _53046_ (_01339_, _01338_, _01323_);
  nor _53047_ (_39722_, _01339_, rst);
  and _53048_ (_01340_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _53049_ (_01341_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _53050_ (_01342_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _53051_ (_01343_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _53052_ (_01344_, _01343_, _01342_);
  and _53053_ (_01345_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _53054_ (_01346_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _53055_ (_01347_, _01346_, _01345_);
  and _53056_ (_01348_, _01347_, _01344_);
  and _53057_ (_01349_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _53058_ (_01350_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _53059_ (_01351_, _01350_, _01349_);
  and _53060_ (_01352_, _01351_, _01348_);
  nor _53061_ (_01353_, _01352_, _37742_);
  nor _53062_ (_01354_, _01353_, _01341_);
  nor _53063_ (_01355_, _01354_, _43140_);
  nor _53064_ (_01356_, _01355_, _01340_);
  nor _53065_ (_39723_, _01356_, rst);
  and _53066_ (_01357_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _53067_ (_01358_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _53068_ (_01359_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _53069_ (_01360_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _53070_ (_01361_, _01360_, _01359_);
  and _53071_ (_01362_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _53072_ (_01363_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _53073_ (_01364_, _01363_, _01362_);
  and _53074_ (_01365_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _53075_ (_01366_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _53076_ (_01367_, _01366_, _01365_);
  and _53077_ (_01368_, _01367_, _01364_);
  and _53078_ (_01369_, _01368_, _01361_);
  nor _53079_ (_01370_, _01369_, _37742_);
  nor _53080_ (_01371_, _01370_, _01358_);
  nor _53081_ (_01372_, _01371_, _43140_);
  nor _53082_ (_01373_, _01372_, _01357_);
  nor _53083_ (_39724_, _01373_, rst);
  and _53084_ (_01374_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _53085_ (_01375_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _53086_ (_01376_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _53087_ (_01377_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _53088_ (_01378_, _01377_, _01376_);
  and _53089_ (_01379_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _53090_ (_01380_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _53091_ (_01381_, _01380_, _01379_);
  and _53092_ (_01382_, _01381_, _01378_);
  and _53093_ (_01383_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _53094_ (_01384_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _53095_ (_01385_, _01384_, _01383_);
  and _53096_ (_01386_, _01385_, _01382_);
  nor _53097_ (_01387_, _01386_, _37742_);
  nor _53098_ (_01388_, _01387_, _01375_);
  nor _53099_ (_01389_, _01388_, _43140_);
  nor _53100_ (_01390_, _01389_, _01374_);
  nor _53101_ (_39725_, _01390_, rst);
  and _53102_ (_01391_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _53103_ (_01392_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _53104_ (_01393_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _53105_ (_01394_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _53106_ (_01395_, _01394_, _01393_);
  and _53107_ (_01396_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _53108_ (_01397_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _53109_ (_01398_, _01397_, _01396_);
  and _53110_ (_01399_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _53111_ (_01400_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _53112_ (_01401_, _01400_, _01399_);
  and _53113_ (_01402_, _01401_, _01398_);
  and _53114_ (_01403_, _01402_, _01395_);
  nor _53115_ (_01404_, _01403_, _37742_);
  nor _53116_ (_01405_, _01404_, _01392_);
  nor _53117_ (_01406_, _01405_, _43140_);
  nor _53118_ (_01407_, _01406_, _01391_);
  nor _53119_ (_39726_, _01407_, rst);
  and _53120_ (_01408_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _53121_ (_01409_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _53122_ (_01410_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _53123_ (_01411_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _53124_ (_01412_, _01411_, _01410_);
  and _53125_ (_01413_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _53126_ (_01414_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _53127_ (_01415_, _01414_, _01413_);
  and _53128_ (_01416_, _01415_, _01412_);
  and _53129_ (_01417_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _53130_ (_01418_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _53131_ (_01419_, _01418_, _01417_);
  and _53132_ (_01420_, _01419_, _01416_);
  nor _53133_ (_01421_, _01420_, _37742_);
  nor _53134_ (_01422_, _01421_, _01409_);
  nor _53135_ (_01423_, _01422_, _43140_);
  nor _53136_ (_01424_, _01423_, _01408_);
  nor _53137_ (_39728_, _01424_, rst);
  and _53138_ (_01425_, _43140_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _53139_ (_01426_, _37742_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _53140_ (_01427_, _37774_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _53141_ (_01428_, _37818_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _53142_ (_01429_, _01428_, _01427_);
  and _53143_ (_01430_, _37883_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _53144_ (_01431_, _37960_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _53145_ (_01432_, _01431_, _01430_);
  and _53146_ (_01433_, _01432_, _01429_);
  and _53147_ (_01434_, _37862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _53148_ (_01435_, _37916_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _53149_ (_01436_, _01435_, _01434_);
  and _53150_ (_01437_, _01436_, _01433_);
  nor _53151_ (_01438_, _01437_, _37742_);
  nor _53152_ (_01439_, _01438_, _01426_);
  nor _53153_ (_01440_, _01439_, _43140_);
  nor _53154_ (_01441_, _01440_, _01425_);
  nor _53155_ (_39729_, _01441_, rst);
  and _53156_ (_01442_, _37687_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _53157_ (_01443_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _53158_ (_01444_, _01442_, _39414_);
  and _53159_ (_01445_, _01444_, _43634_);
  and _53160_ (_39751_, _01445_, _01443_);
  not _53161_ (_01446_, _01442_);
  or _53162_ (_01447_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _53163_ (_01448_, _37687_, _43634_);
  and _53164_ (_00000_, _01448_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _53165_ (_01449_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _43634_);
  or _53166_ (_01450_, _01449_, _00000_);
  and _53167_ (_39752_, _01450_, _01447_);
  nor _53168_ (_39789_, _43243_, rst);
  nor _53169_ (_39791_, _43304_, rst);
  nor _53170_ (_39792_, _43221_, rst);
  nor _53171_ (_01451_, _43202_, _28611_);
  and _53172_ (_01452_, _43202_, _28611_);
  nor _53173_ (_01453_, _01452_, _01451_);
  nor _53174_ (_01454_, _43326_, _29061_);
  and _53175_ (_01455_, _43326_, _29061_);
  nor _53176_ (_01456_, _01455_, _01454_);
  nor _53177_ (_01457_, _01456_, _01453_);
  nor _53178_ (_01458_, _43404_, _28918_);
  and _53179_ (_01459_, _43404_, _28918_);
  nor _53180_ (_01460_, _01459_, _01458_);
  not _53181_ (_01461_, _01460_);
  not _53182_ (_01462_, _43555_);
  nor _53183_ (_01463_, _43450_, _28490_);
  and _53184_ (_01464_, _43450_, _28490_);
  nor _53185_ (_01465_, _01464_, _01463_);
  nor _53186_ (_01466_, _01465_, _01462_);
  and _53187_ (_01467_, _01466_, _01461_);
  and _53188_ (_01468_, _01467_, _01457_);
  nor _53189_ (_01469_, _43365_, _28250_);
  and _53190_ (_01470_, _43365_, _28250_);
  nor _53191_ (_01471_, _01470_, _01469_);
  nor _53192_ (_01472_, _01471_, _40057_);
  and _53193_ (_01473_, _43285_, _34487_);
  nor _53194_ (_01474_, _43285_, _34487_);
  or _53195_ (_01475_, _01474_, _01473_);
  nor _53196_ (_01476_, _43161_, _28008_);
  and _53197_ (_01477_, _43161_, _28008_);
  nor _53198_ (_01478_, _01477_, _01476_);
  nor _53199_ (_01479_, _01478_, _01475_);
  and _53200_ (_01480_, _01479_, _01472_);
  and _53201_ (_01481_, _01480_, _01468_);
  nor _53202_ (_01482_, _28765_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _53203_ (_01483_, _01482_, _01481_);
  not _53204_ (_01484_, _01483_);
  nor _53205_ (_01485_, _39182_, _39199_);
  nor _53206_ (_01486_, _32463_, _40695_);
  and _53207_ (_01487_, _01486_, _01468_);
  and _53208_ (_01488_, _01487_, _01485_);
  and _53209_ (_01489_, _39088_, _39079_);
  and _53210_ (_01490_, _01489_, _39091_);
  not _53211_ (_01491_, _39988_);
  and _53212_ (_01492_, _01491_, _01490_);
  not _53213_ (_01493_, _01492_);
  not _53214_ (_01494_, _39164_);
  nor _53215_ (_01495_, _00836_, _39081_);
  nor _53216_ (_01496_, _01101_, _39113_);
  and _53217_ (_01497_, _01496_, _01070_);
  not _53218_ (_01498_, _01497_);
  nor _53219_ (_01499_, _01498_, _00908_);
  nor _53220_ (_01500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _53221_ (_01501_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _53222_ (_01502_, _01501_, _01500_);
  nor _53223_ (_01503_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _53224_ (_01504_, _01503_, _01502_);
  and _53225_ (_01505_, _01504_, _39951_);
  nand _53226_ (_01506_, _01505_, _01490_);
  or _53227_ (_01507_, _01506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _53228_ (_01508_, _01485_, _30102_);
  not _53229_ (_01509_, _01508_);
  nand _53230_ (_01510_, _35042_, _30234_);
  nor _53231_ (_01511_, _01510_, _35390_);
  and _53232_ (_01512_, _01511_, _36217_);
  and _53233_ (_01513_, _01512_, _36903_);
  and _53234_ (_01514_, _01513_, _30397_);
  nor _53235_ (_01515_, _01485_, _39093_);
  and _53236_ (_01516_, _01515_, _32833_);
  and _53237_ (_01517_, _01516_, _01514_);
  and _53238_ (_01518_, _00833_, _39091_);
  and _53239_ (_01519_, _01518_, _39074_);
  and _53240_ (_01520_, _01519_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _53241_ (_01521_, _01520_, _01517_);
  and _53242_ (_01522_, _01521_, _01509_);
  and _53243_ (_01523_, _01522_, _01507_);
  not _53244_ (_01524_, _39088_);
  or _53245_ (_01525_, _39175_, _39080_);
  nor _53246_ (_01526_, _01525_, _39149_);
  nor _53247_ (_01527_, _01526_, _01524_);
  not _53248_ (_01528_, _01527_);
  and _53249_ (_01529_, _01528_, _01523_);
  and _53250_ (_01530_, _01529_, _01499_);
  and _53251_ (_01531_, _00833_, _39000_);
  or _53252_ (_01532_, _01531_, _39180_);
  or _53253_ (_01533_, _01532_, _01523_);
  nor _53254_ (_01534_, _01533_, _39179_);
  or _53255_ (_01535_, _01534_, _01530_);
  and _53256_ (_01536_, _01535_, _01495_);
  and _53257_ (_01537_, _01536_, _01494_);
  nor _53258_ (_01538_, _01537_, _43205_);
  nor _53259_ (_01539_, _01094_, _37633_);
  nor _53260_ (_01540_, _01539_, _39201_);
  not _53261_ (_01541_, _01540_);
  nor _53262_ (_01542_, _01541_, _01538_);
  nor _53263_ (_01543_, _39754_, _39744_);
  and _53264_ (_01544_, _01543_, _43107_);
  not _53265_ (_01545_, _01544_);
  and _53266_ (_01546_, _01545_, _01519_);
  nor _53267_ (_01547_, _01546_, _01542_);
  and _53268_ (_01548_, _01547_, _01493_);
  not _53269_ (_01549_, _01548_);
  nor _53270_ (_01550_, _01549_, _01488_);
  and _53271_ (_01551_, _01550_, _01484_);
  nor _53272_ (_01552_, _39201_, rst);
  and _53273_ (_39796_, _01552_, _01551_);
  and _53274_ (_39797_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _43634_);
  and _53275_ (_39798_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _43634_);
  not _53276_ (_01553_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _53277_ (_01554_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _53278_ (_01555_, _01554_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _53279_ (_01556_, _01555_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _53280_ (_01557_, _01556_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53281_ (_01558_, _01557_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _53282_ (_01559_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _53283_ (_01560_, _01559_, _01558_);
  and _53284_ (_01561_, _01560_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _53285_ (_01562_, _01561_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _53286_ (_01563_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _53287_ (_01564_, _37764_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _53288_ (_01565_, _01564_, _43140_);
  nor _53289_ (_01566_, _01565_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _53290_ (_01567_, _01566_);
  and _53291_ (_01568_, _01567_, _01563_);
  and _53292_ (_01569_, _01568_, _01562_);
  nand _53293_ (_01570_, _01569_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _53294_ (_01571_, _01570_, _01553_);
  or _53295_ (_01572_, _01570_, _01553_);
  and _53296_ (_01573_, _01572_, _01571_);
  or _53297_ (_01574_, _01573_, _01551_);
  and _53298_ (_01575_, _01574_, _43634_);
  not _53299_ (_01576_, _01322_);
  nor _53300_ (_01577_, _43205_, _39182_);
  not _53301_ (_01578_, _01577_);
  nor _53302_ (_01579_, _01497_, _43205_);
  and _53303_ (_01580_, _01093_, _37622_);
  not _53304_ (_01581_, _01580_);
  and _53305_ (_01582_, _39158_, _37622_);
  and _53306_ (_01583_, _01582_, _39088_);
  nor _53307_ (_01584_, _01583_, _39201_);
  and _53308_ (_01585_, _01584_, _01581_);
  not _53309_ (_01586_, _01585_);
  nor _53310_ (_01587_, _01586_, _01579_);
  and _53311_ (_01588_, _01587_, _01578_);
  nor _53312_ (_01589_, _01588_, _01576_);
  and _53313_ (_01590_, _01588_, _43238_);
  nor _53314_ (_01591_, _01590_, _01589_);
  and _53315_ (_01592_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _53316_ (_01593_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _53317_ (_01594_, _01441_);
  nor _53318_ (_01595_, _01588_, _01594_);
  and _53319_ (_01596_, _01588_, _43445_);
  nor _53320_ (_01597_, _01596_, _01595_);
  and _53321_ (_01598_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _53322_ (_01599_, _01597_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _53323_ (_01600_, _01599_, _01598_);
  not _53324_ (_01601_, _01424_);
  nor _53325_ (_01602_, _01588_, _01601_);
  and _53326_ (_01603_, _01588_, _43184_);
  nor _53327_ (_01604_, _01603_, _01602_);
  and _53328_ (_01605_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _53329_ (_01606_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _53330_ (_01607_, _01407_);
  nor _53331_ (_01608_, _01588_, _01607_);
  and _53332_ (_01609_, _01588_, _43300_);
  nor _53333_ (_01610_, _01609_, _01608_);
  nand _53334_ (_01611_, _01610_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _53335_ (_01612_, _01390_);
  nor _53336_ (_01613_, _01588_, _01612_);
  and _53337_ (_01614_, _01588_, _43399_);
  nor _53338_ (_01616_, _01614_, _01613_);
  and _53339_ (_01617_, _01616_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _53340_ (_01619_, _01616_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _53341_ (_01620_, _01373_);
  nor _53342_ (_01622_, _01588_, _01620_);
  and _53343_ (_01623_, _01588_, _43156_);
  nor _53344_ (_01625_, _01623_, _01622_);
  and _53345_ (_01626_, _01625_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _53346_ (_01628_, _01356_);
  nor _53347_ (_01629_, _01588_, _01628_);
  and _53348_ (_01631_, _01588_, _43276_);
  nor _53349_ (_01632_, _01631_, _01629_);
  and _53350_ (_01634_, _01632_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _53351_ (_01635_, _01339_);
  nor _53352_ (_01637_, _01588_, _01635_);
  and _53353_ (_01638_, _01588_, _43360_);
  nor _53354_ (_01640_, _01638_, _01637_);
  and _53355_ (_01641_, _01640_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _53356_ (_01643_, _01632_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _53357_ (_01644_, _01643_, _01634_);
  and _53358_ (_01646_, _01644_, _01641_);
  nor _53359_ (_01647_, _01646_, _01634_);
  not _53360_ (_01648_, _01647_);
  nor _53361_ (_01649_, _01625_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _53362_ (_01650_, _01649_, _01626_);
  and _53363_ (_01651_, _01650_, _01648_);
  nor _53364_ (_01652_, _01651_, _01626_);
  nor _53365_ (_01653_, _01652_, _01619_);
  or _53366_ (_01654_, _01653_, _01617_);
  or _53367_ (_01655_, _01610_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _53368_ (_01656_, _01655_, _01611_);
  nand _53369_ (_01657_, _01656_, _01654_);
  and _53370_ (_01658_, _01657_, _01611_);
  nor _53371_ (_01659_, _01658_, _01606_);
  or _53372_ (_01660_, _01659_, _01605_);
  and _53373_ (_01661_, _01660_, _01600_);
  nor _53374_ (_01662_, _01661_, _01598_);
  nor _53375_ (_01663_, _01662_, _01593_);
  or _53376_ (_01664_, _01663_, _01592_);
  and _53377_ (_01665_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53378_ (_01666_, _01665_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _53379_ (_01667_, _01666_, _01664_);
  and _53380_ (_01668_, _01667_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _53381_ (_01669_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53382_ (_01670_, _01669_, _01668_);
  nor _53383_ (_01671_, _01670_, _01591_);
  not _53384_ (_01672_, _01591_);
  nor _53385_ (_01673_, _01664_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53386_ (_01674_, _01673_, _39392_);
  and _53387_ (_01675_, _01674_, _39397_);
  and _53388_ (_01676_, _01675_, _39382_);
  and _53389_ (_01677_, _01676_, _39403_);
  and _53390_ (_01678_, _01677_, _39378_);
  nor _53391_ (_01679_, _01678_, _01672_);
  nor _53392_ (_01680_, _01679_, _01671_);
  or _53393_ (_01681_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _53394_ (_01682_, _01591_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53395_ (_01683_, _01682_, _01681_);
  and _53396_ (_01684_, _01683_, _01680_);
  or _53397_ (_01685_, _01684_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _53398_ (_01686_, _01684_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _53399_ (_01687_, _39088_, _37622_);
  and _53400_ (_01688_, _01687_, _39158_);
  not _53401_ (_01689_, _01688_);
  nor _53402_ (_01690_, _00908_, _00833_);
  and _53403_ (_01691_, _01690_, _01495_);
  nand _53404_ (_01692_, _01691_, _01497_);
  and _53405_ (_01693_, _01692_, _39091_);
  nor _53406_ (_01694_, _01693_, _01577_);
  and _53407_ (_01695_, _01694_, _01689_);
  not _53408_ (_01696_, _01588_);
  and _53409_ (_01697_, _39081_, _39091_);
  nor _53410_ (_01698_, _01697_, _01539_);
  nor _53411_ (_01699_, _01698_, _01696_);
  nor _53412_ (_01700_, _01699_, _01695_);
  and _53413_ (_01701_, _01700_, _01686_);
  and _53414_ (_01702_, _01701_, _01685_);
  and _53415_ (_01703_, _39201_, _31820_);
  not _53416_ (_01704_, _39463_);
  and _53417_ (_01705_, _01697_, _01704_);
  and _53418_ (_01706_, _01587_, _01539_);
  and _53419_ (_01707_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _53420_ (_01708_, _01707_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53421_ (_01709_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _53422_ (_01710_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _53423_ (_01711_, _01710_, _01709_);
  and _53424_ (_01712_, _01711_, _01708_);
  and _53425_ (_01713_, _01712_, _01666_);
  and _53426_ (_01714_, _01713_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _53427_ (_01715_, _01714_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53428_ (_01716_, _01715_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _53429_ (_01717_, _01716_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _53430_ (_01718_, _01717_, _39414_);
  or _53431_ (_01719_, _01717_, _39414_);
  and _53432_ (_01720_, _01719_, _01718_);
  and _53433_ (_01721_, _01720_, _01706_);
  and _53434_ (_01722_, _01580_, _43239_);
  and _53435_ (_01723_, _01698_, _01587_);
  and _53436_ (_01724_, _01723_, _01695_);
  and _53437_ (_01725_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _53438_ (_01726_, _01725_, _01722_);
  or _53439_ (_01727_, _01726_, _01721_);
  nor _53440_ (_01728_, _01727_, _01705_);
  nand _53441_ (_01729_, _01728_, _01551_);
  or _53442_ (_01730_, _01729_, _01703_);
  or _53443_ (_01731_, _01730_, _01702_);
  and _53444_ (_39799_, _01731_, _01575_);
  and _53445_ (_01732_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _43634_);
  and _53446_ (_01733_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _53447_ (_01734_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _53448_ (_01735_, _37676_, _01734_);
  not _53449_ (_01736_, _01735_);
  not _53450_ (_01737_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _53451_ (_01738_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _53452_ (_01739_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _53453_ (_01740_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _53454_ (_01741_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _53455_ (_01742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _53456_ (_01743_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _53457_ (_01744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _53458_ (_01745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53459_ (_01746_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _53460_ (_01747_, _01746_, _01745_);
  and _53461_ (_01748_, _01747_, _01744_);
  and _53462_ (_01749_, _01748_, _01743_);
  and _53463_ (_01750_, _01749_, _01742_);
  and _53464_ (_01751_, _01750_, _01741_);
  and _53465_ (_01752_, _01751_, _01740_);
  and _53466_ (_01753_, _01752_, _01739_);
  and _53467_ (_01754_, _01753_, _01738_);
  and _53468_ (_01755_, _01754_, _01737_);
  nor _53469_ (_01756_, _01755_, _01553_);
  and _53470_ (_01757_, _01755_, _01553_);
  nor _53471_ (_01758_, _01757_, _01756_);
  nor _53472_ (_01759_, _01754_, _01737_);
  nor _53473_ (_01760_, _01759_, _01755_);
  and _53474_ (_01761_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _53475_ (_01762_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _53476_ (_01763_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _53477_ (_01764_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _53478_ (_01765_, _01764_, _01762_);
  and _53479_ (_01766_, _01765_, _01763_);
  nor _53480_ (_01767_, _01766_, _01762_);
  nor _53481_ (_01768_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _53482_ (_01769_, _01768_, _01761_);
  not _53483_ (_01770_, _01769_);
  nor _53484_ (_01771_, _01770_, _01767_);
  nor _53485_ (_01772_, _01771_, _01761_);
  not _53486_ (_01773_, _01772_);
  and _53487_ (_01774_, _01773_, _01752_);
  and _53488_ (_01775_, _01774_, _01739_);
  and _53489_ (_01776_, _01775_, _01738_);
  not _53490_ (_01777_, _01776_);
  nor _53491_ (_01778_, _01777_, _01760_);
  and _53492_ (_01779_, _01777_, _01760_);
  or _53493_ (_01780_, _01779_, _01778_);
  not _53494_ (_01781_, _01780_);
  and _53495_ (_01782_, _01772_, _01754_);
  and _53496_ (_01783_, _01772_, _01753_);
  nor _53497_ (_01784_, _01783_, _01738_);
  nor _53498_ (_01785_, _01784_, _01782_);
  not _53499_ (_01786_, _01785_);
  and _53500_ (_01787_, _01772_, _01752_);
  nor _53501_ (_01788_, _01787_, _01739_);
  nor _53502_ (_01789_, _01788_, _01783_);
  not _53503_ (_01790_, _01789_);
  and _53504_ (_01791_, _01772_, _01750_);
  and _53505_ (_01792_, _01791_, _01741_);
  nor _53506_ (_01793_, _01792_, _01740_);
  nor _53507_ (_01794_, _01793_, _01787_);
  not _53508_ (_01795_, _01794_);
  nor _53509_ (_01796_, _01791_, _01741_);
  nor _53510_ (_01797_, _01796_, _01792_);
  not _53511_ (_01798_, _01797_);
  not _53512_ (_01799_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _53513_ (_01800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _53514_ (_01801_, _01772_, _01749_);
  and _53515_ (_01802_, _01801_, _01800_);
  nor _53516_ (_01803_, _01802_, _01799_);
  nor _53517_ (_01804_, _01803_, _01791_);
  not _53518_ (_01805_, _01804_);
  and _53519_ (_01806_, _01772_, _01747_);
  and _53520_ (_01807_, _01806_, _01744_);
  nor _53521_ (_01808_, _01807_, _01743_);
  nor _53522_ (_01809_, _01808_, _01801_);
  not _53523_ (_01810_, _01809_);
  nor _53524_ (_01811_, _01806_, _01744_);
  or _53525_ (_01812_, _01811_, _01807_);
  and _53526_ (_01813_, _01772_, _01746_);
  nor _53527_ (_01814_, _01813_, _01745_);
  nor _53528_ (_01815_, _01814_, _01806_);
  not _53529_ (_01816_, _01815_);
  not _53530_ (_01817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _53531_ (_01818_, _01772_, _01817_);
  nor _53532_ (_01819_, _01772_, _01817_);
  nor _53533_ (_01820_, _01819_, _01818_);
  not _53534_ (_01821_, _01820_);
  not _53535_ (_01822_, _00745_);
  and _53536_ (_01823_, _00750_, _00738_);
  or _53537_ (_01824_, _01823_, _00802_);
  not _53538_ (_01825_, _01824_);
  and _53539_ (_01826_, _00784_, _00738_);
  not _53540_ (_01827_, _01826_);
  and _53541_ (_01828_, _00793_, _00738_);
  nor _53542_ (_01829_, _01828_, _00767_);
  and _53543_ (_01830_, _01829_, _01827_);
  and _53544_ (_01831_, _01830_, _01825_);
  nor _53545_ (_01832_, _01831_, _01822_);
  not _53546_ (_01833_, _01832_);
  and _53547_ (_01834_, _01833_, _00805_);
  and _53548_ (_01835_, _00802_, _00787_);
  nor _53549_ (_01836_, _01835_, _00766_);
  not _53550_ (_01837_, _00802_);
  nor _53551_ (_01838_, _00777_, _00739_);
  and _53552_ (_01839_, _01838_, _01837_);
  nor _53553_ (_01840_, _01839_, _01836_);
  not _53554_ (_01841_, _01840_);
  and _53555_ (_01842_, _00787_, _00751_);
  not _53556_ (_01843_, _01842_);
  nor _53557_ (_01844_, _00817_, _00746_);
  and _53558_ (_01845_, _01844_, _01843_);
  and _53559_ (_01846_, _01845_, _01841_);
  and _53560_ (_01847_, _01846_, _01834_);
  not _53561_ (_01848_, _00766_);
  nor _53562_ (_01849_, _01826_, _00751_);
  nor _53563_ (_01850_, _01849_, _01848_);
  not _53564_ (_01851_, _01850_);
  nor _53565_ (_01852_, _00785_, _00777_);
  nor _53566_ (_01853_, _01852_, _01822_);
  and _53567_ (_01854_, _00751_, _00745_);
  and _53568_ (_01855_, _00773_, _00737_);
  and _53569_ (_01856_, _00779_, _01855_);
  or _53570_ (_01857_, _01856_, _01854_);
  nor _53571_ (_01858_, _01857_, _01853_);
  and _53572_ (_01859_, _01858_, _01851_);
  and _53573_ (_01860_, _00802_, _00779_);
  and _53574_ (_01861_, _00785_, _00766_);
  nor _53575_ (_01862_, _01861_, _01860_);
  not _53576_ (_01863_, _00760_);
  and _53577_ (_01864_, _00738_, _39018_);
  and _53578_ (_01865_, _00793_, _00748_);
  nor _53579_ (_01866_, _01865_, _01864_);
  nor _53580_ (_01867_, _01866_, _01863_);
  and _53581_ (_01868_, _00748_, _00737_);
  nor _53582_ (_01869_, _01868_, _00751_);
  nor _53583_ (_01870_, _01869_, _01863_);
  nor _53584_ (_01871_, _01870_, _01867_);
  and _53585_ (_01872_, _01871_, _01862_);
  nor _53586_ (_01873_, _00769_, _00756_);
  and _53587_ (_01874_, _00794_, _00778_);
  and _53588_ (_01875_, _00753_, _38535_);
  and _53589_ (_01876_, _00748_, _00749_);
  and _53590_ (_01877_, _01876_, _01875_);
  nor _53591_ (_01878_, _01877_, _01874_);
  and _53592_ (_01879_, _01878_, _01873_);
  not _53593_ (_01880_, _00786_);
  and _53594_ (_01881_, _01880_, _00776_);
  and _53595_ (_01882_, _01881_, _01879_);
  and _53596_ (_01883_, _01882_, _01872_);
  and _53597_ (_01884_, _00808_, _00788_);
  and _53598_ (_01885_, _00785_, _00752_);
  nor _53599_ (_01886_, _01885_, _01884_);
  and _53600_ (_01887_, _00800_, _00787_);
  not _53601_ (_01888_, _00777_);
  nor _53602_ (_01889_, _01875_, _00787_);
  nor _53603_ (_01890_, _01889_, _01888_);
  nor _53604_ (_01891_, _01890_, _01887_);
  and _53605_ (_01892_, _01891_, _01886_);
  nor _53606_ (_01893_, _01865_, _00777_);
  nor _53607_ (_01894_, _01893_, _38535_);
  not _53608_ (_01895_, _00744_);
  nor _53609_ (_01896_, _01868_, _00794_);
  nor _53610_ (_01897_, _01896_, _01895_);
  nor _53611_ (_01898_, _01897_, _01894_);
  nor _53612_ (_01899_, _01865_, _01868_);
  nor _53613_ (_01900_, _01899_, _01848_);
  not _53614_ (_01901_, _01855_);
  nor _53615_ (_01902_, _00766_, _00744_);
  nor _53616_ (_01903_, _01902_, _01901_);
  nor _53617_ (_01904_, _01903_, _01900_);
  and _53618_ (_01905_, _01904_, _01898_);
  and _53619_ (_01906_, _01905_, _01892_);
  and _53620_ (_01907_, _01906_, _01883_);
  and _53621_ (_01908_, _01907_, _01859_);
  and _53622_ (_01909_, _01908_, _01847_);
  not _53623_ (_01910_, _01909_);
  nor _53624_ (_01911_, _01765_, _01763_);
  nor _53625_ (_01912_, _01911_, _01766_);
  nand _53626_ (_01913_, _01912_, _01910_);
  or _53627_ (_01914_, _01860_, _00801_);
  and _53628_ (_01915_, _00794_, _00779_);
  and _53629_ (_01916_, _01868_, _00760_);
  nor _53630_ (_01917_, _01916_, _01915_);
  nand _53631_ (_01918_, _01917_, _01873_);
  nor _53632_ (_01919_, _01918_, _01914_);
  and _53633_ (_01920_, _01919_, _01858_);
  nand _53634_ (_01921_, _01920_, _01845_);
  nor _53635_ (_01922_, _01921_, _01909_);
  not _53636_ (_01923_, _01922_);
  nor _53637_ (_01924_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _53638_ (_01925_, _01924_, _01763_);
  and _53639_ (_01926_, _01925_, _01923_);
  or _53640_ (_01927_, _01912_, _01910_);
  and _53641_ (_01928_, _01927_, _01913_);
  nand _53642_ (_01929_, _01928_, _01926_);
  and _53643_ (_01930_, _01929_, _01913_);
  not _53644_ (_01931_, _01930_);
  and _53645_ (_01932_, _01770_, _01767_);
  nor _53646_ (_01933_, _01932_, _01771_);
  and _53647_ (_01934_, _01933_, _01931_);
  and _53648_ (_01935_, _01934_, _01821_);
  not _53649_ (_01936_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53650_ (_01937_, _01818_, _01936_);
  or _53651_ (_01938_, _01937_, _01813_);
  and _53652_ (_01939_, _01938_, _01935_);
  and _53653_ (_01940_, _01939_, _01816_);
  and _53654_ (_01941_, _01940_, _01812_);
  and _53655_ (_01942_, _01941_, _01810_);
  nor _53656_ (_01943_, _01801_, _01800_);
  or _53657_ (_01944_, _01943_, _01802_);
  and _53658_ (_01945_, _01944_, _01942_);
  and _53659_ (_01946_, _01945_, _01805_);
  and _53660_ (_01947_, _01946_, _01798_);
  and _53661_ (_01948_, _01947_, _01795_);
  and _53662_ (_01949_, _01948_, _01790_);
  and _53663_ (_01950_, _01949_, _01786_);
  and _53664_ (_01951_, _01950_, _01781_);
  nor _53665_ (_01952_, _01951_, _01778_);
  not _53666_ (_01953_, _01952_);
  nor _53667_ (_01954_, _01953_, _01758_);
  and _53668_ (_01955_, _01953_, _01758_);
  or _53669_ (_01956_, _01955_, _01954_);
  or _53670_ (_01957_, _01956_, _01736_);
  or _53671_ (_01958_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _53672_ (_01959_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _53673_ (_01960_, _01959_, _01958_);
  and _53674_ (_01961_, _01960_, _01957_);
  or _53675_ (_39801_, _01961_, _01733_);
  nor _53676_ (_01962_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _53677_ (_39802_, _01962_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _53678_ (_39803_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _43634_);
  nor _53679_ (_01963_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _53680_ (_01964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _53681_ (_01965_, _01964_, _01963_);
  nor _53682_ (_01966_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _53683_ (_01967_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _53684_ (_01968_, _01967_, _01966_);
  and _53685_ (_01969_, _01968_, _01965_);
  nor _53686_ (_01970_, _01969_, rst);
  and _53687_ (_01971_, \oc8051_top_1.oc8051_rom1.ea_int , _37644_);
  nand _53688_ (_01972_, _01971_, _37676_);
  and _53689_ (_01973_, _01972_, _39803_);
  or _53690_ (_39804_, _01973_, _01970_);
  and _53691_ (_01974_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _53692_ (_01975_, _01974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _53693_ (_39806_, _01975_, _43634_);
  nor _53694_ (_01976_, _01566_, _43140_);
  or _53695_ (_01977_, _01909_, _37796_);
  nor _53696_ (_01978_, _01922_, _37938_);
  nand _53697_ (_01979_, _01909_, _37796_);
  and _53698_ (_01980_, _01979_, _01977_);
  nand _53699_ (_01981_, _01980_, _01978_);
  and _53700_ (_01982_, _01981_, _01977_);
  nor _53701_ (_01983_, _01982_, _43140_);
  and _53702_ (_01984_, _01983_, _37753_);
  nor _53703_ (_01985_, _01983_, _37753_);
  nor _53704_ (_01986_, _01985_, _01984_);
  nor _53705_ (_01987_, _01986_, _01976_);
  and _53706_ (_01988_, _37807_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _53707_ (_01989_, _01988_, _01976_);
  and _53708_ (_01990_, _01989_, _01921_);
  or _53709_ (_01991_, _01990_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53710_ (_01992_, _01991_, _01987_);
  and _53711_ (_39807_, _01992_, _43634_);
  not _53712_ (_01993_, _38491_);
  nand _53713_ (_01994_, _39014_, _01993_);
  nor _53714_ (_01995_, _01994_, _39037_);
  nand _53715_ (_01996_, _39060_, _38744_);
  nor _53716_ (_01997_, _01996_, _38988_);
  not _53717_ (_01998_, _01448_);
  or _53718_ (_01999_, _01998_, _38228_);
  nor _53719_ (_02000_, _01999_, _38014_);
  and _53720_ (_02001_, _02000_, _01997_);
  and _53721_ (_39810_, _02001_, _01995_);
  nor _53722_ (_02002_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _53723_ (_02003_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _53724_ (_02004_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _53725_ (_39813_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _43634_);
  and _53726_ (_02005_, _39813_, _02004_);
  or _53727_ (_39811_, _02005_, _02003_);
  not _53728_ (_02006_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _53729_ (_02007_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53730_ (_02008_, _02007_, _02006_);
  and _53731_ (_02009_, _02007_, _02006_);
  nor _53732_ (_02010_, _02009_, _02008_);
  not _53733_ (_02011_, _02010_);
  and _53734_ (_02012_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _53735_ (_02013_, _02012_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53736_ (_02014_, _02012_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _53737_ (_02015_, _02014_, _02013_);
  or _53738_ (_02016_, _02015_, _02007_);
  and _53739_ (_02017_, _02016_, _02011_);
  nor _53740_ (_02018_, _02008_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _53741_ (_02019_, _02008_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _53742_ (_02020_, _02019_, _02018_);
  or _53743_ (_02021_, _02013_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _53744_ (_39815_, _02021_, _43634_);
  and _53745_ (_02022_, _39815_, _02020_);
  and _53746_ (_39814_, _02022_, _02017_);
  not _53747_ (_02023_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _53748_ (_02024_, _01566_, _02023_);
  and _53749_ (_02025_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _53750_ (_02026_, _02024_);
  and _53751_ (_02027_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _53752_ (_02028_, _02027_, _02025_);
  and _53753_ (_39816_, _02028_, _43634_);
  and _53754_ (_02029_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _53755_ (_02030_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _53756_ (_02031_, _02030_, _02029_);
  and _53757_ (_39817_, _02031_, _43634_);
  and _53758_ (_02032_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _53759_ (_02033_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53760_ (_02034_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _02033_);
  and _53761_ (_02035_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _53762_ (_02036_, _02035_, _02032_);
  and _53763_ (_39818_, _02036_, _43634_);
  and _53764_ (_02037_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53765_ (_02038_, _02037_, _02034_);
  and _53766_ (_39819_, _02038_, _43634_);
  or _53767_ (_02039_, _02033_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _53768_ (_39821_, _02039_, _43634_);
  not _53769_ (_02040_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _53770_ (_02041_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _53771_ (_02042_, _02041_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53772_ (_02043_, _02033_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _53773_ (_02044_, _02043_, _43634_);
  and _53774_ (_39822_, _02044_, _02042_);
  or _53775_ (_02045_, _02033_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _53776_ (_39823_, _02045_, _43634_);
  nor _53777_ (_02046_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _53778_ (_02047_, _02046_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53779_ (_02048_, _02047_, _43634_);
  and _53780_ (_02049_, _39813_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _53781_ (_39824_, _02049_, _02048_);
  and _53782_ (_02050_, _02023_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _53783_ (_02051_, _02050_, _02047_);
  and _53784_ (_39825_, _02051_, _43634_);
  nand _53785_ (_02052_, _02047_, _39463_);
  or _53786_ (_02053_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _53787_ (_02054_, _02053_, _43634_);
  and _53788_ (_39826_, _02054_, _02052_);
  nand _53789_ (_02055_, _39105_, _43634_);
  nor _53790_ (_39827_, _02055_, _39237_);
  or _53791_ (_02056_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _53792_ (_02057_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand _53793_ (_02058_, _01442_, _02057_);
  and _53794_ (_02059_, _02058_, _43634_);
  and _53795_ (_39863_, _02059_, _02056_);
  or _53796_ (_02060_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _53797_ (_02061_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _53798_ (_02062_, _01442_, _02061_);
  and _53799_ (_02063_, _02062_, _43634_);
  and _53800_ (_39864_, _02063_, _02060_);
  or _53801_ (_02064_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _53802_ (_02065_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _53803_ (_02066_, _01442_, _02065_);
  and _53804_ (_02067_, _02066_, _43634_);
  and _53805_ (_39865_, _02067_, _02064_);
  or _53806_ (_02068_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _53807_ (_02069_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _53808_ (_02070_, _01442_, _02069_);
  and _53809_ (_02071_, _02070_, _43634_);
  and _53810_ (_39866_, _02071_, _02068_);
  or _53811_ (_02072_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _53812_ (_02073_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _53813_ (_02074_, _01442_, _02073_);
  and _53814_ (_02075_, _02074_, _43634_);
  and _53815_ (_39867_, _02075_, _02072_);
  or _53816_ (_02076_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _53817_ (_02077_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _53818_ (_02078_, _01442_, _02077_);
  and _53819_ (_02079_, _02078_, _43634_);
  and _53820_ (_39869_, _02079_, _02076_);
  or _53821_ (_02080_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not _53822_ (_02081_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand _53823_ (_02082_, _01442_, _02081_);
  and _53824_ (_02083_, _02082_, _43634_);
  and _53825_ (_39870_, _02083_, _02080_);
  or _53826_ (_02084_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _53827_ (_02085_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _53828_ (_02086_, _01442_, _02085_);
  and _53829_ (_02087_, _02086_, _43634_);
  and _53830_ (_39871_, _02087_, _02084_);
  or _53831_ (_02088_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _53832_ (_02089_, _01442_, _39386_);
  and _53833_ (_02090_, _02089_, _43634_);
  and _53834_ (_39872_, _02090_, _02088_);
  or _53835_ (_02091_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _53836_ (_02092_, _01442_, _39392_);
  and _53837_ (_02093_, _02092_, _43634_);
  and _53838_ (_39873_, _02093_, _02091_);
  or _53839_ (_02094_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _53840_ (_02095_, _01442_, _39397_);
  and _53841_ (_02096_, _02095_, _43634_);
  and _53842_ (_39874_, _02096_, _02094_);
  or _53843_ (_02097_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _53844_ (_02098_, _01442_, _39382_);
  and _53845_ (_02099_, _02098_, _43634_);
  and _53846_ (_39875_, _02099_, _02097_);
  or _53847_ (_02100_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _53848_ (_02101_, _01442_, _39403_);
  and _53849_ (_02102_, _02101_, _43634_);
  and _53850_ (_39876_, _02102_, _02100_);
  or _53851_ (_02103_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _53852_ (_02104_, _01442_, _39378_);
  and _53853_ (_02105_, _02104_, _43634_);
  and _53854_ (_39877_, _02105_, _02103_);
  or _53855_ (_02106_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _53856_ (_02107_, _01442_, _39409_);
  and _53857_ (_02108_, _02107_, _43634_);
  and _53858_ (_39878_, _02108_, _02106_);
  and _53859_ (_02109_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _53860_ (_02110_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _53861_ (_02111_, _02110_, _02109_);
  and _53862_ (_39883_, _02111_, _43634_);
  and _53863_ (_02112_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53864_ (_02113_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _53865_ (_02114_, _02113_, _02112_);
  and _53866_ (_39884_, _02114_, _43634_);
  and _53867_ (_02115_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53868_ (_02116_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _53869_ (_02117_, _02116_, _02115_);
  and _53870_ (_39885_, _02117_, _43634_);
  and _53871_ (_02118_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53872_ (_02119_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53873_ (_02120_, _02119_, _02118_);
  and _53874_ (_39886_, _02120_, _43634_);
  and _53875_ (_02121_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _53876_ (_02122_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _53877_ (_02123_, _02122_, _02121_);
  and _53878_ (_39887_, _02123_, _43634_);
  and _53879_ (_02124_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _53880_ (_02125_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _53881_ (_02126_, _02125_, _02124_);
  and _53882_ (_39888_, _02126_, _43634_);
  and _53883_ (_02127_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _53884_ (_02128_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or _53885_ (_02129_, _02128_, _02127_);
  and _53886_ (_39889_, _02129_, _43634_);
  and _53887_ (_02130_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _53888_ (_02132_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or _53889_ (_02134_, _02132_, _02130_);
  and _53890_ (_39890_, _02134_, _43634_);
  and _53891_ (_02137_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _53892_ (_02139_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _53893_ (_02141_, _02139_, _02137_);
  and _53894_ (_39891_, _02141_, _43634_);
  and _53895_ (_02144_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _53896_ (_02146_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _53897_ (_02148_, _02146_, _02144_);
  and _53898_ (_39892_, _02148_, _43634_);
  and _53899_ (_02151_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _53900_ (_02153_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _53901_ (_02155_, _02153_, _02151_);
  and _53902_ (_39894_, _02155_, _43634_);
  and _53903_ (_02158_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _53904_ (_02160_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _53905_ (_02162_, _02160_, _02158_);
  and _53906_ (_39895_, _02162_, _43634_);
  and _53907_ (_02165_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _53908_ (_02167_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or _53909_ (_02169_, _02167_, _02165_);
  and _53910_ (_39896_, _02169_, _43634_);
  and _53911_ (_02172_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _53912_ (_02174_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _53913_ (_02176_, _02174_, _02172_);
  and _53914_ (_39897_, _02176_, _43634_);
  and _53915_ (_02179_, _01442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _53916_ (_02181_, _01446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _53917_ (_02183_, _02181_, _02179_);
  and _53918_ (_39898_, _02183_, _43634_);
  and _53919_ (_40076_, _38124_, _43634_);
  and _53920_ (_40077_, _38337_, _43634_);
  and _53921_ (_40078_, _38832_, _43634_);
  nor _53922_ (_40079_, _43109_, rst);
  and _53923_ (_02189_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _53924_ (_02190_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _53925_ (_02191_, _02190_, _02189_);
  and _53926_ (_40080_, _02191_, _43634_);
  and _53927_ (_02192_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _53928_ (_02193_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _53929_ (_02194_, _02193_, _02192_);
  and _53930_ (_40081_, _02194_, _43634_);
  and _53931_ (_02195_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _53932_ (_02196_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _53933_ (_02197_, _02196_, _02195_);
  and _53934_ (_40082_, _02197_, _43634_);
  and _53935_ (_02198_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _53936_ (_02199_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _53937_ (_02200_, _02199_, _02198_);
  and _53938_ (_40083_, _02200_, _43634_);
  and _53939_ (_02201_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _53940_ (_02202_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _53941_ (_02203_, _02202_, _02201_);
  and _53942_ (_40084_, _02203_, _43634_);
  and _53943_ (_02204_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _53944_ (_02205_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _53945_ (_02206_, _02205_, _02204_);
  and _53946_ (_40085_, _02206_, _43634_);
  and _53947_ (_02207_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _53948_ (_02208_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _53949_ (_02209_, _02208_, _02207_);
  and _53950_ (_40086_, _02209_, _43634_);
  and _53951_ (_02210_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _53952_ (_02211_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _53953_ (_02212_, _02211_, _02210_);
  and _53954_ (_40087_, _02212_, _43634_);
  and _53955_ (_02213_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _53956_ (_02214_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _53957_ (_02215_, _02214_, _02213_);
  and _53958_ (_40088_, _02215_, _43634_);
  and _53959_ (_02216_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _53960_ (_02217_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _53961_ (_02218_, _02217_, _02216_);
  and _53962_ (_40089_, _02218_, _43634_);
  and _53963_ (_02219_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _53964_ (_02220_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _53965_ (_02221_, _02220_, _02219_);
  and _53966_ (_40090_, _02221_, _43634_);
  and _53967_ (_02222_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _53968_ (_02223_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _53969_ (_02224_, _02223_, _02222_);
  and _53970_ (_40091_, _02224_, _43634_);
  and _53971_ (_02225_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _53972_ (_02226_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _53973_ (_02227_, _02226_, _02225_);
  and _53974_ (_40092_, _02227_, _43634_);
  and _53975_ (_02228_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _53976_ (_02229_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _53977_ (_02230_, _02229_, _02228_);
  and _53978_ (_40093_, _02230_, _43634_);
  and _53979_ (_02231_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _53980_ (_02232_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _53981_ (_02233_, _02232_, _02231_);
  and _53982_ (_40095_, _02233_, _43634_);
  and _53983_ (_02234_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _53984_ (_02235_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _53985_ (_02236_, _02235_, _02234_);
  and _53986_ (_40096_, _02236_, _43634_);
  and _53987_ (_02237_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _53988_ (_02238_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _53989_ (_02239_, _02238_, _02237_);
  and _53990_ (_40097_, _02239_, _43634_);
  and _53991_ (_02240_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _53992_ (_02241_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _53993_ (_02242_, _02241_, _02240_);
  and _53994_ (_40098_, _02242_, _43634_);
  and _53995_ (_02243_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _53996_ (_02244_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _53997_ (_02245_, _02244_, _02243_);
  and _53998_ (_40099_, _02245_, _43634_);
  and _53999_ (_02246_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _54000_ (_02247_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _54001_ (_02248_, _02247_, _02246_);
  and _54002_ (_40100_, _02248_, _43634_);
  and _54003_ (_02249_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _54004_ (_02250_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _54005_ (_02251_, _02250_, _02249_);
  and _54006_ (_40101_, _02251_, _43634_);
  and _54007_ (_02252_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _54008_ (_02253_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _54009_ (_02254_, _02253_, _02252_);
  and _54010_ (_40102_, _02254_, _43634_);
  and _54011_ (_02255_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _54012_ (_02256_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _54013_ (_02257_, _02256_, _02255_);
  and _54014_ (_40103_, _02257_, _43634_);
  and _54015_ (_02258_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _54016_ (_02259_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _54017_ (_02260_, _02259_, _02258_);
  and _54018_ (_40104_, _02260_, _43634_);
  and _54019_ (_02261_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _54020_ (_02262_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _54021_ (_02263_, _02262_, _02261_);
  and _54022_ (_40106_, _02263_, _43634_);
  and _54023_ (_02264_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _54024_ (_02265_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _54025_ (_02266_, _02265_, _02264_);
  and _54026_ (_40107_, _02266_, _43634_);
  and _54027_ (_02267_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _54028_ (_02268_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _54029_ (_02269_, _02268_, _02267_);
  and _54030_ (_40108_, _02269_, _43634_);
  and _54031_ (_02270_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _54032_ (_02271_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _54033_ (_02272_, _02271_, _02270_);
  and _54034_ (_40109_, _02272_, _43634_);
  and _54035_ (_02273_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _54036_ (_02274_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _54037_ (_02275_, _02274_, _02273_);
  and _54038_ (_40110_, _02275_, _43634_);
  and _54039_ (_02276_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _54040_ (_02277_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _54041_ (_02278_, _02277_, _02276_);
  and _54042_ (_40111_, _02278_, _43634_);
  and _54043_ (_02279_, _02024_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _54044_ (_02280_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _54045_ (_02281_, _02280_, _02279_);
  and _54046_ (_40112_, _02281_, _43634_);
  nor _54047_ (_40113_, _43339_, rst);
  nor _54048_ (_40115_, _43258_, rst);
  nor _54049_ (_40116_, _43128_, rst);
  nor _54050_ (_40117_, _43377_, rst);
  nor _54051_ (_40118_, _43318_, rst);
  nor _54052_ (_40119_, _43197_, rst);
  nor _54053_ (_40121_, _43427_, rst);
  and _54054_ (_40137_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _43634_);
  and _54055_ (_40138_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _43634_);
  and _54056_ (_40139_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _43634_);
  and _54057_ (_40140_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _43634_);
  and _54058_ (_40141_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _43634_);
  and _54059_ (_40143_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _43634_);
  and _54060_ (_40144_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _43634_);
  or _54061_ (_02282_, _01724_, _01697_);
  and _54062_ (_02283_, _02282_, _32964_);
  and _54063_ (_02284_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _54064_ (_02285_, _01580_, _01635_);
  and _54065_ (_02286_, _01706_, _43361_);
  or _54066_ (_02287_, _02286_, _02285_);
  or _54067_ (_02288_, _02287_, _02284_);
  nor _54068_ (_02289_, _01640_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _54069_ (_02290_, _02289_, _01641_);
  and _54070_ (_02291_, _02290_, _01700_);
  nor _54071_ (_02292_, _02291_, _02288_);
  nand _54072_ (_02293_, _02292_, _01551_);
  or _54073_ (_02294_, _02293_, _02283_);
  or _54074_ (_02295_, _01551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _54075_ (_02296_, _02295_, _43634_);
  and _54076_ (_40145_, _02296_, _02294_);
  or _54077_ (_02297_, _01551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _54078_ (_02298_, _02297_, _43634_);
  and _54079_ (_02299_, _02282_, _33650_);
  and _54080_ (_02300_, _01706_, _43277_);
  and _54081_ (_02301_, _01580_, _01628_);
  and _54082_ (_02302_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _54083_ (_02303_, _02302_, _02301_);
  or _54084_ (_02304_, _02303_, _02300_);
  or _54085_ (_02305_, _02304_, _02299_);
  nor _54086_ (_02306_, _01644_, _01641_);
  nor _54087_ (_02307_, _02306_, _01646_);
  nand _54088_ (_02308_, _02307_, _01700_);
  nand _54089_ (_02309_, _02308_, _01551_);
  or _54090_ (_02310_, _02309_, _02305_);
  and _54091_ (_40146_, _02310_, _02298_);
  not _54092_ (_02311_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _54093_ (_02312_, _01566_, _02311_);
  and _54094_ (_02313_, _01566_, _02311_);
  nor _54095_ (_02314_, _02313_, _02312_);
  or _54096_ (_02315_, _02314_, _01551_);
  and _54097_ (_02316_, _02315_, _43634_);
  and _54098_ (_02317_, _02282_, _34389_);
  or _54099_ (_02318_, _01650_, _01648_);
  not _54100_ (_02319_, _01651_);
  and _54101_ (_02320_, _01700_, _02319_);
  and _54102_ (_02321_, _02320_, _02318_);
  and _54103_ (_02322_, _01706_, _43157_);
  and _54104_ (_02323_, _01580_, _01620_);
  and _54105_ (_02324_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _54106_ (_02325_, _02324_, _02323_);
  or _54107_ (_02326_, _02325_, _02322_);
  nor _54108_ (_02327_, _02326_, _02321_);
  nand _54109_ (_02328_, _02327_, _01551_);
  or _54110_ (_02329_, _02328_, _02317_);
  and _54111_ (_40147_, _02329_, _02316_);
  and _54112_ (_02330_, _02312_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _54113_ (_02331_, _02312_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _54114_ (_02332_, _02331_, _02330_);
  or _54115_ (_02333_, _02332_, _01551_);
  and _54116_ (_02334_, _02333_, _43634_);
  and _54117_ (_02335_, _02282_, _35129_);
  and _54118_ (_02336_, _01706_, _43400_);
  and _54119_ (_02337_, _01580_, _01612_);
  and _54120_ (_02338_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _54121_ (_02339_, _02338_, _02337_);
  or _54122_ (_02340_, _02339_, _02336_);
  or _54123_ (_02341_, _01619_, _01617_);
  or _54124_ (_02342_, _02341_, _01652_);
  nand _54125_ (_02343_, _02341_, _01652_);
  and _54126_ (_02344_, _02343_, _01700_);
  and _54127_ (_02345_, _02344_, _02342_);
  nor _54128_ (_02346_, _02345_, _02340_);
  nand _54129_ (_02347_, _02346_, _01551_);
  or _54130_ (_02348_, _02347_, _02335_);
  and _54131_ (_40148_, _02348_, _02334_);
  and _54132_ (_02350_, _01555_, _01567_);
  nor _54133_ (_02351_, _02330_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _54134_ (_02352_, _02351_, _02350_);
  or _54135_ (_02353_, _02352_, _01551_);
  and _54136_ (_02354_, _02353_, _43634_);
  and _54137_ (_02355_, _02282_, _35891_);
  or _54138_ (_02356_, _01656_, _01654_);
  and _54139_ (_02357_, _01700_, _01657_);
  and _54140_ (_02358_, _02357_, _02356_);
  and _54141_ (_02359_, _01706_, _43301_);
  and _54142_ (_02360_, _01580_, _01607_);
  and _54143_ (_02361_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _54144_ (_02362_, _02361_, _02360_);
  or _54145_ (_02363_, _02362_, _02359_);
  nor _54146_ (_02364_, _02363_, _02358_);
  nand _54147_ (_02365_, _02364_, _01551_);
  or _54148_ (_02366_, _02365_, _02355_);
  and _54149_ (_40149_, _02366_, _02354_);
  and _54150_ (_02367_, _02282_, _36686_);
  or _54151_ (_02368_, _01606_, _01605_);
  nand _54152_ (_02369_, _02368_, _01658_);
  or _54153_ (_02370_, _02368_, _01658_);
  and _54154_ (_02371_, _02370_, _01700_);
  and _54155_ (_02372_, _02371_, _02369_);
  and _54156_ (_02373_, _01580_, _01601_);
  and _54157_ (_02374_, _01706_, _43185_);
  and _54158_ (_02375_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _54159_ (_02376_, _02375_, _02374_);
  or _54160_ (_02377_, _02376_, _02373_);
  nor _54161_ (_02378_, _02377_, _02372_);
  nand _54162_ (_02379_, _02378_, _01551_);
  or _54163_ (_02380_, _02379_, _02367_);
  and _54164_ (_02381_, _01556_, _01567_);
  nor _54165_ (_02382_, _02350_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _54166_ (_02383_, _02382_, _02381_);
  or _54167_ (_02384_, _02383_, _01551_);
  and _54168_ (_02385_, _02384_, _43634_);
  and _54169_ (_40150_, _02385_, _02380_);
  not _54170_ (_02386_, _01551_);
  nor _54171_ (_02387_, _01660_, _01600_);
  nor _54172_ (_02388_, _02387_, _01661_);
  and _54173_ (_02389_, _02388_, _01700_);
  and _54174_ (_02390_, _02282_, _37414_);
  and _54175_ (_02391_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _54176_ (_02392_, _01580_, _01594_);
  and _54177_ (_02393_, _01706_, _43446_);
  or _54178_ (_02394_, _02393_, _02392_);
  or _54179_ (_02395_, _02394_, _02391_);
  or _54180_ (_02396_, _02395_, _02390_);
  or _54181_ (_02397_, _02396_, _02389_);
  or _54182_ (_02398_, _02397_, _02386_);
  and _54183_ (_02399_, _02381_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _54184_ (_02400_, _02381_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _54185_ (_02401_, _02400_, _02399_);
  or _54186_ (_02402_, _02401_, _01551_);
  and _54187_ (_02403_, _02402_, _43634_);
  and _54188_ (_40151_, _02403_, _02398_);
  and _54189_ (_02404_, _02282_, _31820_);
  or _54190_ (_02405_, _01592_, _01593_);
  or _54191_ (_02406_, _02405_, _01662_);
  nand _54192_ (_02407_, _02405_, _01662_);
  and _54193_ (_02408_, _02407_, _01700_);
  and _54194_ (_02409_, _02408_, _02406_);
  and _54195_ (_02410_, _01580_, _01576_);
  and _54196_ (_02411_, _01706_, _43239_);
  and _54197_ (_02412_, _39201_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _54198_ (_02413_, _02412_, _02411_);
  nor _54199_ (_02414_, _02413_, _02410_);
  nand _54200_ (_02415_, _02414_, _01551_);
  or _54201_ (_02416_, _02415_, _02409_);
  or _54202_ (_02417_, _02416_, _02404_);
  and _54203_ (_02418_, _02399_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _54204_ (_02419_, _02399_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _54205_ (_02420_, _02419_, _02418_);
  or _54206_ (_02421_, _02420_, _01551_);
  and _54207_ (_02422_, _02421_, _43634_);
  and _54208_ (_40152_, _02422_, _02417_);
  and _54209_ (_02423_, _39201_, _32964_);
  not _54210_ (_02424_, _39507_);
  and _54211_ (_02425_, _01697_, _02424_);
  and _54212_ (_02426_, _01664_, _39386_);
  nor _54213_ (_02427_, _01664_, _39386_);
  nor _54214_ (_02428_, _02427_, _02426_);
  nor _54215_ (_02429_, _02428_, _01591_);
  and _54216_ (_02430_, _02428_, _01591_);
  or _54217_ (_02431_, _02430_, _02429_);
  and _54218_ (_02432_, _02431_, _01700_);
  and _54219_ (_02433_, _01580_, _43361_);
  and _54220_ (_02434_, _01706_, _00761_);
  and _54221_ (_02435_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _54222_ (_02436_, _02435_, _02434_);
  nor _54223_ (_02437_, _02436_, _02433_);
  nand _54224_ (_02438_, _02437_, _01551_);
  or _54225_ (_02439_, _02438_, _02432_);
  or _54226_ (_02440_, _02439_, _02425_);
  or _54227_ (_02441_, _02440_, _02423_);
  and _54228_ (_02442_, _02418_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _54229_ (_02443_, _02418_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _54230_ (_02444_, _02443_, _02442_);
  or _54231_ (_02445_, _02444_, _01551_);
  and _54232_ (_02446_, _02445_, _43634_);
  and _54233_ (_40154_, _02446_, _02441_);
  and _54234_ (_02447_, _01560_, _01567_);
  nor _54235_ (_02448_, _02442_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _54236_ (_02449_, _02448_, _02447_);
  or _54237_ (_02450_, _02449_, _01551_);
  and _54238_ (_02451_, _02450_, _43634_);
  and _54239_ (_02452_, _39201_, _33650_);
  and _54240_ (_02453_, _01664_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _54241_ (_02454_, _02453_, _01672_);
  and _54242_ (_02455_, _01673_, _01591_);
  nor _54243_ (_02456_, _02455_, _02454_);
  nand _54244_ (_02457_, _02456_, _39392_);
  or _54245_ (_02458_, _02456_, _39392_);
  and _54246_ (_02459_, _02458_, _02457_);
  and _54247_ (_02460_, _02459_, _01700_);
  not _54248_ (_02461_, _39539_);
  and _54249_ (_02462_, _01697_, _02461_);
  and _54250_ (_02463_, _01580_, _43277_);
  not _54251_ (_02464_, _39064_);
  and _54252_ (_02465_, _01706_, _02464_);
  and _54253_ (_02466_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _54254_ (_02467_, _02466_, _02465_);
  or _54255_ (_02468_, _02467_, _02463_);
  nor _54256_ (_02469_, _02468_, _02462_);
  nand _54257_ (_02470_, _02469_, _01551_);
  or _54258_ (_02471_, _02470_, _02460_);
  or _54259_ (_02472_, _02471_, _02452_);
  and _54260_ (_40155_, _02472_, _02451_);
  and _54261_ (_02473_, _39201_, _34389_);
  and _54262_ (_02474_, _01674_, _01591_);
  and _54263_ (_02475_, _02454_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _54264_ (_02476_, _02475_, _02474_);
  nor _54265_ (_02477_, _02476_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _54266_ (_02478_, _02476_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _54267_ (_02479_, _02478_, _02477_);
  and _54268_ (_02480_, _02479_, _01700_);
  not _54269_ (_02481_, _39569_);
  and _54270_ (_02482_, _01697_, _02481_);
  and _54271_ (_02483_, _01706_, _00747_);
  and _54272_ (_02484_, _01580_, _43157_);
  and _54273_ (_02485_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _54274_ (_02486_, _02485_, _02484_);
  or _54275_ (_02487_, _02486_, _02483_);
  nor _54276_ (_02488_, _02487_, _02482_);
  nand _54277_ (_02489_, _02488_, _01551_);
  or _54278_ (_02490_, _02489_, _02480_);
  or _54279_ (_02491_, _02490_, _02473_);
  and _54280_ (_02492_, _02447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _54281_ (_02493_, _02447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _54282_ (_02494_, _02493_, _02492_);
  or _54283_ (_02495_, _02494_, _01551_);
  and _54284_ (_02496_, _02495_, _43634_);
  and _54285_ (_40156_, _02496_, _02491_);
  and _54286_ (_02497_, _39201_, _35129_);
  and _54287_ (_02498_, _01667_, _01672_);
  and _54288_ (_02499_, _01675_, _01591_);
  nor _54289_ (_02500_, _02499_, _02498_);
  nor _54290_ (_02501_, _02500_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _54291_ (_02502_, _02500_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _54292_ (_02503_, _02502_, _02501_);
  and _54293_ (_02504_, _02503_, _01700_);
  not _54294_ (_02505_, _39600_);
  and _54295_ (_02506_, _01697_, _02505_);
  and _54296_ (_02507_, _01580_, _43400_);
  nor _54297_ (_02508_, _01713_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _54298_ (_02509_, _02508_, _01714_);
  and _54299_ (_02510_, _02509_, _01706_);
  and _54300_ (_02511_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _54301_ (_02512_, _02511_, _02510_);
  or _54302_ (_02513_, _02512_, _02507_);
  nor _54303_ (_02514_, _02513_, _02506_);
  nand _54304_ (_02515_, _02514_, _01551_);
  or _54305_ (_02516_, _02515_, _02504_);
  or _54306_ (_02517_, _02516_, _02497_);
  and _54307_ (_02518_, _02492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _54308_ (_02519_, _02492_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _54309_ (_02520_, _02519_, _02518_);
  or _54310_ (_02521_, _02520_, _01551_);
  and _54311_ (_02522_, _02521_, _43634_);
  and _54312_ (_40157_, _02522_, _02517_);
  and _54313_ (_02523_, _02518_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _54314_ (_02524_, _02518_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _54315_ (_02525_, _02524_, _02523_);
  or _54316_ (_02526_, _02525_, _01551_);
  and _54317_ (_02527_, _02526_, _43634_);
  and _54318_ (_02528_, _39201_, _35891_);
  and _54319_ (_02529_, _01668_, _01672_);
  and _54320_ (_02530_, _01676_, _01591_);
  nor _54321_ (_02531_, _02530_, _02529_);
  nand _54322_ (_02532_, _02531_, _39403_);
  or _54323_ (_02533_, _02531_, _39403_);
  and _54324_ (_02534_, _02533_, _01700_);
  and _54325_ (_02535_, _02534_, _02532_);
  not _54326_ (_02536_, _39631_);
  nand _54327_ (_02537_, _01697_, _02536_);
  and _54328_ (_02538_, _01580_, _43301_);
  nor _54329_ (_02539_, _01714_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _54330_ (_02540_, _02539_, _01715_);
  and _54331_ (_02542_, _02540_, _01706_);
  and _54332_ (_02543_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _54333_ (_02544_, _02543_, _02542_);
  nor _54334_ (_02545_, _02544_, _02538_);
  and _54335_ (_02546_, _02545_, _02537_);
  nand _54336_ (_02547_, _02546_, _01551_);
  or _54337_ (_02548_, _02547_, _02535_);
  or _54338_ (_02549_, _02548_, _02528_);
  and _54339_ (_40158_, _02549_, _02527_);
  and _54340_ (_02550_, _39201_, _36686_);
  and _54341_ (_02551_, _02529_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _54342_ (_02552_, _01677_, _01591_);
  nor _54343_ (_02553_, _02552_, _02551_);
  nand _54344_ (_02554_, _02553_, _39378_);
  or _54345_ (_02555_, _02553_, _39378_);
  and _54346_ (_02556_, _02555_, _01700_);
  and _54347_ (_02557_, _02556_, _02554_);
  not _54348_ (_02558_, _39664_);
  and _54349_ (_02559_, _01697_, _02558_);
  and _54350_ (_02560_, _01580_, _43185_);
  nor _54351_ (_02561_, _01715_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _54352_ (_02562_, _02561_, _01716_);
  and _54353_ (_02563_, _02562_, _01706_);
  and _54354_ (_02565_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _54355_ (_02566_, _02565_, _02563_);
  or _54356_ (_02567_, _02566_, _02560_);
  nor _54357_ (_02568_, _02567_, _02559_);
  nand _54358_ (_02569_, _02568_, _01551_);
  or _54359_ (_02570_, _02569_, _02557_);
  or _54360_ (_02571_, _02570_, _02550_);
  or _54361_ (_02572_, _02523_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _54362_ (_02573_, _02523_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _54363_ (_02574_, _02573_, _02572_);
  or _54364_ (_02575_, _02574_, _01551_);
  and _54365_ (_02577_, _02575_, _43634_);
  and _54366_ (_40159_, _02577_, _02571_);
  nand _54367_ (_02578_, _01680_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _54368_ (_02579_, _01680_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _54369_ (_02580_, _02579_, _01700_);
  and _54370_ (_02581_, _02580_, _02578_);
  and _54371_ (_02582_, _39201_, _37414_);
  not _54372_ (_02583_, _39693_);
  and _54373_ (_02584_, _01697_, _02583_);
  or _54374_ (_02585_, _01716_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _54375_ (_02586_, _02585_, _01717_);
  and _54376_ (_02587_, _02586_, _01706_);
  and _54377_ (_02588_, _01580_, _43446_);
  and _54378_ (_02589_, _01724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _54379_ (_02590_, _02589_, _02588_);
  or _54380_ (_02591_, _02590_, _02587_);
  nor _54381_ (_02592_, _02591_, _02584_);
  nand _54382_ (_02593_, _02592_, _01551_);
  or _54383_ (_02594_, _02593_, _02582_);
  or _54384_ (_02595_, _02594_, _02581_);
  or _54385_ (_02596_, _01569_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _54386_ (_02597_, _02596_, _01570_);
  or _54387_ (_02598_, _02597_, _01551_);
  and _54388_ (_02599_, _02598_, _43634_);
  and _54389_ (_40160_, _02599_, _02595_);
  or _54390_ (_02600_, _01925_, _01923_);
  nor _54391_ (_02601_, _01736_, _01926_);
  and _54392_ (_02602_, _02601_, _02600_);
  nor _54393_ (_02603_, _01735_, _02057_);
  or _54394_ (_02604_, _02603_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _54395_ (_02605_, _02604_, _02602_);
  or _54396_ (_02606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _37644_);
  and _54397_ (_02607_, _02606_, _43634_);
  and _54398_ (_40161_, _02607_, _02605_);
  or _54399_ (_02608_, _01928_, _01926_);
  and _54400_ (_02609_, _02608_, _01929_);
  or _54401_ (_02610_, _02609_, _01736_);
  or _54402_ (_02611_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _54403_ (_02612_, _02611_, _01959_);
  and _54404_ (_02613_, _02612_, _02610_);
  and _54405_ (_02614_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _54406_ (_40162_, _02614_, _02613_);
  and _54407_ (_02615_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _54408_ (_02616_, _01933_, _01931_);
  nor _54409_ (_02617_, _02616_, _01934_);
  or _54410_ (_02618_, _02617_, _01736_);
  or _54411_ (_02619_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _54412_ (_02620_, _02619_, _01959_);
  and _54413_ (_02621_, _02620_, _02618_);
  or _54414_ (_40163_, _02621_, _02615_);
  and _54415_ (_02622_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _54416_ (_02623_, _01934_, _01821_);
  nor _54417_ (_02624_, _02623_, _01935_);
  or _54418_ (_02625_, _02624_, _01736_);
  or _54419_ (_02626_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _54420_ (_02627_, _02626_, _01959_);
  and _54421_ (_02628_, _02627_, _02625_);
  or _54422_ (_40165_, _02628_, _02622_);
  and _54423_ (_02629_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _54424_ (_02630_, _01938_, _01935_);
  nor _54425_ (_02631_, _02630_, _01939_);
  or _54426_ (_02632_, _02631_, _01736_);
  or _54427_ (_02633_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _54428_ (_02634_, _02633_, _01959_);
  and _54429_ (_02635_, _02634_, _02632_);
  or _54430_ (_40166_, _02635_, _02629_);
  and _54431_ (_02636_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _54432_ (_02637_, _01939_, _01816_);
  nor _54433_ (_02638_, _02637_, _01940_);
  or _54434_ (_02639_, _02638_, _01736_);
  or _54435_ (_02640_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _54436_ (_02641_, _02640_, _01959_);
  and _54437_ (_02642_, _02641_, _02639_);
  or _54438_ (_40167_, _02642_, _02636_);
  nor _54439_ (_02643_, _01940_, _01812_);
  nor _54440_ (_02644_, _02643_, _01941_);
  or _54441_ (_02645_, _02644_, _01736_);
  or _54442_ (_02646_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _54443_ (_02647_, _02646_, _01959_);
  and _54444_ (_02648_, _02647_, _02645_);
  and _54445_ (_02649_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _54446_ (_40168_, _02649_, _02648_);
  nor _54447_ (_02650_, _01941_, _01810_);
  nor _54448_ (_02651_, _02650_, _01942_);
  or _54449_ (_02652_, _02651_, _01736_);
  or _54450_ (_02653_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _54451_ (_02654_, _02653_, _01959_);
  and _54452_ (_02655_, _02654_, _02652_);
  and _54453_ (_02656_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _54454_ (_40169_, _02656_, _02655_);
  and _54455_ (_02657_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _54456_ (_02658_, _01944_, _01942_);
  nor _54457_ (_02659_, _02658_, _01945_);
  or _54458_ (_02660_, _02659_, _01736_);
  or _54459_ (_02661_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _54460_ (_02662_, _02661_, _01959_);
  and _54461_ (_02663_, _02662_, _02660_);
  or _54462_ (_40170_, _02663_, _02657_);
  nor _54463_ (_02664_, _01945_, _01805_);
  nor _54464_ (_02665_, _02664_, _01946_);
  or _54465_ (_02666_, _02665_, _01736_);
  or _54466_ (_02667_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _54467_ (_02668_, _02667_, _01959_);
  and _54468_ (_02669_, _02668_, _02666_);
  and _54469_ (_02670_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _54470_ (_40171_, _02670_, _02669_);
  nor _54471_ (_02671_, _01946_, _01798_);
  nor _54472_ (_02672_, _02671_, _01947_);
  or _54473_ (_02673_, _02672_, _01736_);
  or _54474_ (_02674_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _54475_ (_02675_, _02674_, _01959_);
  and _54476_ (_02676_, _02675_, _02673_);
  and _54477_ (_02677_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _54478_ (_40172_, _02677_, _02676_);
  and _54479_ (_02678_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _54480_ (_02679_, _01947_, _01795_);
  nor _54481_ (_02680_, _02679_, _01948_);
  or _54482_ (_02681_, _02680_, _01736_);
  or _54483_ (_02682_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _54484_ (_02683_, _02682_, _01959_);
  and _54485_ (_02684_, _02683_, _02681_);
  or _54486_ (_40173_, _02684_, _02678_);
  and _54487_ (_02685_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _54488_ (_02686_, _01948_, _01790_);
  nor _54489_ (_02687_, _02686_, _01949_);
  or _54490_ (_02688_, _02687_, _01736_);
  or _54491_ (_02689_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _54492_ (_02690_, _02689_, _01959_);
  and _54493_ (_02691_, _02690_, _02688_);
  or _54494_ (_40174_, _02691_, _02685_);
  and _54495_ (_02692_, _01732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _54496_ (_02693_, _01949_, _01786_);
  nor _54497_ (_02694_, _02693_, _01950_);
  or _54498_ (_02695_, _02694_, _01736_);
  or _54499_ (_02696_, _01735_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _54500_ (_02697_, _02696_, _01959_);
  and _54501_ (_02698_, _02697_, _02695_);
  or _54502_ (_40176_, _02698_, _02692_);
  or _54503_ (_02699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _37644_);
  and _54504_ (_02700_, _02699_, _43634_);
  or _54505_ (_02701_, _01950_, _01781_);
  nor _54506_ (_02702_, _01736_, _01951_);
  and _54507_ (_02703_, _02702_, _02701_);
  nor _54508_ (_02704_, _01735_, _39409_);
  or _54509_ (_02705_, _02704_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _54510_ (_02706_, _02705_, _02703_);
  and _54511_ (_40177_, _02706_, _02700_);
  and _54512_ (_02707_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _54513_ (_02708_, _02707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _54514_ (_40178_, _02708_, _43634_);
  and _54515_ (_02709_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _54516_ (_02710_, _02709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _54517_ (_40179_, _02710_, _43634_);
  and _54518_ (_02711_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _54519_ (_02712_, _02711_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _54520_ (_40180_, _02712_, _43634_);
  and _54521_ (_02713_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _54522_ (_02714_, _02713_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _54523_ (_40181_, _02714_, _43634_);
  and _54524_ (_02715_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _54525_ (_02716_, _02715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _54526_ (_40182_, _02716_, _43634_);
  and _54527_ (_02717_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _54528_ (_02718_, _02717_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _54529_ (_40183_, _02718_, _43634_);
  and _54530_ (_02719_, _01969_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _54531_ (_02721_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _54532_ (_40184_, _02721_, _43634_);
  nor _54533_ (_02722_, _01922_, _43140_);
  or _54534_ (_02723_, _02722_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand _54535_ (_02724_, _02722_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _54536_ (_02725_, _02724_, _01959_);
  and _54537_ (_40185_, _02725_, _02723_);
  or _54538_ (_02726_, _01980_, _01978_);
  and _54539_ (_02727_, _02726_, _01981_);
  or _54540_ (_02728_, _02727_, _43140_);
  or _54541_ (_02729_, _37676_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _54542_ (_02730_, _02729_, _01959_);
  and _54543_ (_40187_, _02730_, _02728_);
  and _54544_ (_02731_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _54545_ (_02732_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _54546_ (_02733_, _02732_, _39813_);
  or _54547_ (_40203_, _02733_, _02731_);
  and _54548_ (_02734_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _54549_ (_02735_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _54550_ (_02736_, _02735_, _39813_);
  or _54551_ (_40204_, _02736_, _02734_);
  and _54552_ (_02737_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _54553_ (_02738_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _54554_ (_02739_, _02738_, _39813_);
  or _54555_ (_40205_, _02739_, _02737_);
  and _54556_ (_02740_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _54557_ (_02741_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _54558_ (_02742_, _02741_, _39813_);
  or _54559_ (_40206_, _02742_, _02740_);
  and _54560_ (_02743_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _54561_ (_02744_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _54562_ (_02745_, _02744_, _39813_);
  or _54563_ (_40207_, _02745_, _02743_);
  and _54564_ (_02746_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _54565_ (_02747_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _54566_ (_02748_, _02747_, _39813_);
  or _54567_ (_40209_, _02748_, _02746_);
  and _54568_ (_02749_, _02002_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _54569_ (_02750_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _54570_ (_02751_, _02750_, _39813_);
  or _54571_ (_40210_, _02751_, _02749_);
  and _54572_ (_40211_, _02010_, _43634_);
  nor _54573_ (_40212_, _02020_, rst);
  and _54574_ (_40213_, _02016_, _43634_);
  and _54575_ (_02752_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _54576_ (_02753_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _54577_ (_02754_, _02753_, _02752_);
  and _54578_ (_40214_, _02754_, _43634_);
  and _54579_ (_02755_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _54580_ (_02756_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _54581_ (_02757_, _02756_, _02755_);
  and _54582_ (_40215_, _02757_, _43634_);
  and _54583_ (_02758_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _54584_ (_02759_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _54585_ (_02760_, _02759_, _02758_);
  and _54586_ (_40216_, _02760_, _43634_);
  and _54587_ (_02761_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _54588_ (_02762_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _54589_ (_02763_, _02762_, _02761_);
  and _54590_ (_40217_, _02763_, _43634_);
  and _54591_ (_02764_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _54592_ (_02765_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _54593_ (_02766_, _02765_, _02764_);
  and _54594_ (_40218_, _02766_, _43634_);
  and _54595_ (_02767_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _54596_ (_02768_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _54597_ (_02769_, _02768_, _02767_);
  and _54598_ (_40220_, _02769_, _43634_);
  and _54599_ (_02770_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _54600_ (_02771_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _54601_ (_02772_, _02771_, _02770_);
  and _54602_ (_40221_, _02772_, _43634_);
  and _54603_ (_02773_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _54604_ (_02774_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _54605_ (_02775_, _02774_, _02773_);
  and _54606_ (_40222_, _02775_, _43634_);
  and _54607_ (_02776_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _54608_ (_02777_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _54609_ (_02778_, _02777_, _02776_);
  and _54610_ (_40223_, _02778_, _43634_);
  and _54611_ (_02779_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _54612_ (_02780_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _54613_ (_02781_, _02780_, _02779_);
  and _54614_ (_40224_, _02781_, _43634_);
  and _54615_ (_02782_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _54616_ (_02783_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _54617_ (_02784_, _02783_, _02782_);
  and _54618_ (_40225_, _02784_, _43634_);
  and _54619_ (_02785_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _54620_ (_02786_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _54621_ (_02787_, _02786_, _02785_);
  and _54622_ (_40226_, _02787_, _43634_);
  and _54623_ (_02788_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _54624_ (_02789_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _54625_ (_02790_, _02789_, _02788_);
  and _54626_ (_40227_, _02790_, _43634_);
  and _54627_ (_02791_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _54628_ (_02792_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _54629_ (_02793_, _02792_, _02791_);
  and _54630_ (_40228_, _02793_, _43634_);
  and _54631_ (_02794_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _54632_ (_02795_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _54633_ (_02796_, _02795_, _02794_);
  and _54634_ (_40229_, _02796_, _43634_);
  and _54635_ (_02797_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _54636_ (_02798_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _54637_ (_02799_, _02798_, _02797_);
  and _54638_ (_40231_, _02799_, _43634_);
  and _54639_ (_02800_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _54640_ (_02801_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _54641_ (_02802_, _02801_, _02800_);
  and _54642_ (_40232_, _02802_, _43634_);
  and _54643_ (_02803_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _54644_ (_02804_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _54645_ (_02805_, _02804_, _02803_);
  and _54646_ (_40233_, _02805_, _43634_);
  and _54647_ (_02806_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _54648_ (_02807_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _54649_ (_02808_, _02807_, _02806_);
  and _54650_ (_40234_, _02808_, _43634_);
  and _54651_ (_02809_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _54652_ (_02810_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _54653_ (_02811_, _02810_, _02809_);
  and _54654_ (_40235_, _02811_, _43634_);
  and _54655_ (_02813_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _54656_ (_02814_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _54657_ (_02815_, _02814_, _02813_);
  and _54658_ (_40236_, _02815_, _43634_);
  and _54659_ (_02817_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _54660_ (_02818_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _54661_ (_02819_, _02818_, _02817_);
  and _54662_ (_40237_, _02819_, _43634_);
  and _54663_ (_02820_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _54664_ (_02822_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _54665_ (_02823_, _02822_, _02820_);
  and _54666_ (_40238_, _02823_, _43634_);
  and _54667_ (_02824_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _54668_ (_02825_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _54669_ (_02827_, _02825_, _02824_);
  and _54670_ (_40239_, _02827_, _43634_);
  and _54671_ (_02828_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _54672_ (_02829_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _54673_ (_02830_, _02829_, _02828_);
  and _54674_ (_40240_, _02830_, _43634_);
  and _54675_ (_02832_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _54676_ (_02833_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _54677_ (_02834_, _02833_, _02832_);
  and _54678_ (_40242_, _02834_, _43634_);
  and _54679_ (_02836_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _54680_ (_02837_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _54681_ (_02838_, _02837_, _02836_);
  and _54682_ (_40243_, _02838_, _43634_);
  and _54683_ (_02839_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _54684_ (_02841_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _54685_ (_02842_, _02841_, _02839_);
  and _54686_ (_40244_, _02842_, _43634_);
  and _54687_ (_02844_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _54688_ (_02845_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _54689_ (_02846_, _02845_, _02844_);
  and _54690_ (_40245_, _02846_, _43634_);
  and _54691_ (_02848_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _54692_ (_02849_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _54693_ (_02851_, _02849_, _02848_);
  and _54694_ (_40246_, _02851_, _43634_);
  and _54695_ (_02852_, _02024_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _54696_ (_02854_, _02026_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _54697_ (_02855_, _02854_, _02852_);
  and _54698_ (_40247_, _02855_, _43634_);
  and _54699_ (_02857_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54700_ (_02858_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _54701_ (_02860_, _02858_, _02857_);
  and _54702_ (_40248_, _02860_, _43634_);
  and _54703_ (_02862_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54704_ (_02863_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _54705_ (_02865_, _02863_, _02862_);
  and _54706_ (_40249_, _02865_, _43634_);
  and _54707_ (_02866_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54708_ (_02868_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54709_ (_02869_, _02868_, _02866_);
  and _54710_ (_40250_, _02869_, _43634_);
  and _54711_ (_02871_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54712_ (_02872_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _54713_ (_02874_, _02872_, _02871_);
  and _54714_ (_40251_, _02874_, _43634_);
  and _54715_ (_02875_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54716_ (_02876_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _54717_ (_02877_, _02876_, _02875_);
  and _54718_ (_40253_, _02877_, _43634_);
  and _54719_ (_02878_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54720_ (_02880_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _54721_ (_02882_, _02880_, _02878_);
  and _54722_ (_40254_, _02882_, _43634_);
  and _54723_ (_02884_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _54724_ (_02885_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _54725_ (_02886_, _02885_, _02884_);
  and _54726_ (_40255_, _02886_, _43634_);
  and _54727_ (_02888_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54728_ (_02889_, _43339_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54729_ (_02891_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _54730_ (_02892_, _02891_, _02033_);
  and _54731_ (_02894_, _02892_, _02889_);
  or _54732_ (_02896_, _02894_, _02888_);
  and _54733_ (_40256_, _02896_, _43634_);
  and _54734_ (_02897_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54735_ (_02899_, _43258_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54736_ (_02900_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _54737_ (_02901_, _02900_, _02033_);
  and _54738_ (_02903_, _02901_, _02899_);
  or _54739_ (_02904_, _02903_, _02897_);
  and _54740_ (_40257_, _02904_, _43634_);
  and _54741_ (_02907_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54742_ (_02908_, _43128_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54743_ (_02909_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _54744_ (_02910_, _02909_, _02033_);
  and _54745_ (_02912_, _02910_, _02908_);
  or _54746_ (_02913_, _02912_, _02907_);
  and _54747_ (_40258_, _02913_, _43634_);
  and _54748_ (_02915_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54749_ (_02916_, _43377_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54750_ (_02917_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _54751_ (_02919_, _02917_, _02033_);
  and _54752_ (_02920_, _02919_, _02916_);
  or _54753_ (_02921_, _02920_, _02915_);
  and _54754_ (_40259_, _02921_, _43634_);
  and _54755_ (_02923_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54756_ (_02924_, _43318_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54757_ (_02926_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _54758_ (_02927_, _02926_, _02033_);
  and _54759_ (_02928_, _02927_, _02924_);
  or _54760_ (_02930_, _02928_, _02923_);
  and _54761_ (_40260_, _02930_, _43634_);
  and _54762_ (_02932_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54763_ (_02934_, _43197_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54764_ (_02935_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _54765_ (_02937_, _02935_, _02033_);
  and _54766_ (_02938_, _02937_, _02934_);
  or _54767_ (_02939_, _02938_, _02932_);
  and _54768_ (_40261_, _02939_, _43634_);
  and _54769_ (_02940_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54770_ (_02941_, _43427_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54771_ (_02943_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _54772_ (_02945_, _02943_, _02033_);
  and _54773_ (_02946_, _02945_, _02941_);
  or _54774_ (_02947_, _02946_, _02940_);
  and _54775_ (_40262_, _02947_, _43634_);
  and _54776_ (_02949_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _54777_ (_02950_, _43221_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _54778_ (_02952_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _54779_ (_02953_, _02952_, _02033_);
  and _54780_ (_02954_, _02953_, _02950_);
  or _54781_ (_02957_, _02954_, _02949_);
  and _54782_ (_40264_, _02957_, _43634_);
  and _54783_ (_02958_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _54784_ (_02960_, _02958_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54785_ (_02961_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _02033_);
  and _54786_ (_02962_, _02961_, _43634_);
  and _54787_ (_40265_, _02962_, _02960_);
  and _54788_ (_02964_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _54789_ (_02965_, _02964_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54790_ (_02967_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _02033_);
  and _54791_ (_02969_, _02967_, _43634_);
  and _54792_ (_40266_, _02969_, _02965_);
  and _54793_ (_02971_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _54794_ (_02972_, _02971_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54795_ (_02973_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _02033_);
  and _54796_ (_02975_, _02973_, _43634_);
  and _54797_ (_40267_, _02975_, _02972_);
  and _54798_ (_02976_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _54799_ (_02978_, _02976_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54800_ (_02979_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _02033_);
  and _54801_ (_02981_, _02979_, _43634_);
  and _54802_ (_40268_, _02981_, _02978_);
  and _54803_ (_02983_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _54804_ (_02984_, _02983_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54805_ (_02986_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _02033_);
  and _54806_ (_02987_, _02986_, _43634_);
  and _54807_ (_40269_, _02987_, _02984_);
  and _54808_ (_02989_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _54809_ (_02990_, _02989_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54810_ (_02991_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _02033_);
  and _54811_ (_02994_, _02991_, _43634_);
  and _54812_ (_40270_, _02994_, _02990_);
  and _54813_ (_02995_, _02040_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _54814_ (_02997_, _02995_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54815_ (_02998_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _02033_);
  and _54816_ (_03000_, _02998_, _43634_);
  and _54817_ (_40271_, _03000_, _02997_);
  nand _54818_ (_03001_, _02047_, _32953_);
  or _54819_ (_03002_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _54820_ (_03004_, _03002_, _43634_);
  and _54821_ (_40272_, _03004_, _03001_);
  nand _54822_ (_03006_, _02047_, _33639_);
  or _54823_ (_03008_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _54824_ (_03009_, _03008_, _43634_);
  and _54825_ (_40273_, _03009_, _03006_);
  nand _54826_ (_03011_, _02047_, _34378_);
  or _54827_ (_03012_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _54828_ (_03013_, _03012_, _43634_);
  and _54829_ (_40274_, _03013_, _03011_);
  nand _54830_ (_03015_, _02047_, _35118_);
  or _54831_ (_03017_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _54832_ (_03019_, _03017_, _43634_);
  and _54833_ (_40275_, _03019_, _03015_);
  nand _54834_ (_03020_, _02047_, _35880_);
  or _54835_ (_03022_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _54836_ (_03023_, _03022_, _43634_);
  and _54837_ (_40276_, _03023_, _03020_);
  nand _54838_ (_03025_, _02047_, _36675_);
  or _54839_ (_03026_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _54840_ (_03028_, _03026_, _43634_);
  and _54841_ (_40277_, _03028_, _03025_);
  nand _54842_ (_03030_, _02047_, _37403_);
  or _54843_ (_03031_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _54844_ (_03033_, _03031_, _43634_);
  and _54845_ (_40278_, _03033_, _03030_);
  nand _54846_ (_03034_, _02047_, _31809_);
  or _54847_ (_03036_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _54848_ (_03037_, _03036_, _43634_);
  and _54849_ (_40279_, _03037_, _03034_);
  nand _54850_ (_03039_, _02047_, _39507_);
  or _54851_ (_03040_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _54852_ (_03041_, _03040_, _43634_);
  and _54853_ (_40280_, _03041_, _03039_);
  nand _54854_ (_03043_, _02047_, _39539_);
  or _54855_ (_03044_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _54856_ (_03046_, _03044_, _43634_);
  and _54857_ (_40281_, _03046_, _03043_);
  nand _54858_ (_03047_, _02047_, _39569_);
  or _54859_ (_03049_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _54860_ (_03050_, _03049_, _43634_);
  and _54861_ (_40282_, _03050_, _03047_);
  nand _54862_ (_03052_, _02047_, _39600_);
  or _54863_ (_03053_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _54864_ (_03055_, _03053_, _43634_);
  and _54865_ (_40283_, _03055_, _03052_);
  nand _54866_ (_03056_, _02047_, _39631_);
  or _54867_ (_03057_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _54868_ (_03058_, _03057_, _43634_);
  and _54869_ (_40285_, _03058_, _03056_);
  nand _54870_ (_03059_, _02047_, _39664_);
  or _54871_ (_03061_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _54872_ (_03062_, _03061_, _43634_);
  and _54873_ (_40286_, _03062_, _03059_);
  nand _54874_ (_03064_, _02047_, _39693_);
  or _54875_ (_03065_, _02047_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _54876_ (_03066_, _03065_, _43634_);
  and _54877_ (_40287_, _03066_, _03064_);
  and _54878_ (_40499_, _43093_, _43634_);
  and _54879_ (_03068_, _39924_, _28765_);
  and _54880_ (_03070_, _03068_, _43100_);
  nand _54881_ (_03071_, _03070_, _39327_);
  or _54882_ (_03072_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _54883_ (_03074_, _03072_, _43634_);
  and _54884_ (_40500_, _03074_, _03071_);
  and _54885_ (_03075_, _40315_, _28765_);
  not _54886_ (_03077_, _03075_);
  nor _54887_ (_03078_, _03077_, _39327_);
  not _54888_ (_03079_, _43100_);
  and _54889_ (_03081_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _54890_ (_03082_, _03081_, _03079_);
  or _54891_ (_03084_, _03082_, _03078_);
  or _54892_ (_03085_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _54893_ (_03086_, _03085_, _43634_);
  and _54894_ (_40501_, _03086_, _03084_);
  and _54895_ (_03088_, _28271_, _28929_);
  and _54896_ (_03089_, _03088_, _28765_);
  not _54897_ (_03090_, _03089_);
  nor _54898_ (_03092_, _03090_, _39327_);
  and _54899_ (_03093_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _54900_ (_03094_, _03093_, _03079_);
  or _54901_ (_03096_, _03094_, _03092_);
  or _54902_ (_03097_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _54903_ (_03098_, _03097_, _43634_);
  and _54904_ (_40502_, _03098_, _03096_);
  and _54905_ (_03100_, _41351_, _28765_);
  and _54906_ (_03101_, _03100_, _43100_);
  not _54907_ (_03103_, _03101_);
  and _54908_ (_03104_, _03103_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _54909_ (_03105_, _03103_, _39327_);
  or _54910_ (_03107_, _03105_, _03104_);
  and _54911_ (_40504_, _03107_, _43634_);
  nand _54912_ (_03108_, _03070_, _39306_);
  or _54913_ (_03110_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _54914_ (_03111_, _03110_, _43634_);
  and _54915_ (_40531_, _03111_, _03108_);
  nand _54916_ (_03113_, _03070_, _39298_);
  or _54917_ (_03114_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _54918_ (_03115_, _03114_, _43634_);
  and _54919_ (_40532_, _03115_, _03113_);
  nand _54920_ (_03117_, _03070_, _39291_);
  or _54921_ (_03118_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _54922_ (_03120_, _03118_, _43634_);
  and _54923_ (_40533_, _03120_, _03117_);
  nand _54924_ (_03121_, _03070_, _39284_);
  or _54925_ (_03123_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _54926_ (_03124_, _03123_, _43634_);
  and _54927_ (_40534_, _03124_, _03121_);
  nand _54928_ (_03126_, _03070_, _39276_);
  or _54929_ (_03127_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _54930_ (_03128_, _03127_, _43634_);
  and _54931_ (_40535_, _03128_, _03126_);
  nand _54932_ (_03131_, _03070_, _39268_);
  or _54933_ (_03132_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _54934_ (_03134_, _03132_, _43634_);
  and _54935_ (_40536_, _03134_, _03131_);
  nand _54936_ (_03135_, _03070_, _39261_);
  or _54937_ (_03137_, _03070_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _54938_ (_03138_, _03137_, _43634_);
  and _54939_ (_40537_, _03138_, _03135_);
  nor _54940_ (_03140_, _03077_, _39306_);
  and _54941_ (_03141_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _54942_ (_03142_, _03141_, _03079_);
  or _54943_ (_03144_, _03142_, _03140_);
  or _54944_ (_03145_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _54945_ (_03146_, _03145_, _43634_);
  and _54946_ (_40539_, _03146_, _03144_);
  nor _54947_ (_03148_, _03077_, _39298_);
  and _54948_ (_03149_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _54949_ (_03151_, _03149_, _03079_);
  or _54950_ (_03152_, _03151_, _03148_);
  or _54951_ (_03153_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _54952_ (_03155_, _03153_, _43634_);
  and _54953_ (_40540_, _03155_, _03152_);
  nor _54954_ (_03156_, _03077_, _39291_);
  and _54955_ (_03158_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _54956_ (_03159_, _03158_, _03079_);
  or _54957_ (_03160_, _03159_, _03156_);
  or _54958_ (_03162_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _54959_ (_03163_, _03162_, _43634_);
  and _54960_ (_40541_, _03163_, _03160_);
  nor _54961_ (_03165_, _03077_, _39284_);
  and _54962_ (_03166_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _54963_ (_03168_, _03166_, _03079_);
  or _54964_ (_03169_, _03168_, _03165_);
  or _54965_ (_03170_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _54966_ (_03171_, _03170_, _43634_);
  and _54967_ (_40542_, _03171_, _03169_);
  nor _54968_ (_03173_, _03077_, _39276_);
  and _54969_ (_03174_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _54970_ (_03175_, _03174_, _03079_);
  or _54971_ (_03177_, _03175_, _03173_);
  or _54972_ (_03178_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _54973_ (_03179_, _03178_, _43634_);
  and _54974_ (_40543_, _03179_, _03177_);
  nor _54975_ (_03181_, _03077_, _39268_);
  and _54976_ (_03182_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _54977_ (_03184_, _03182_, _03079_);
  or _54978_ (_03185_, _03184_, _03181_);
  or _54979_ (_03186_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _54980_ (_03188_, _03186_, _43634_);
  and _54981_ (_40544_, _03188_, _03185_);
  nor _54982_ (_03189_, _03077_, _39261_);
  and _54983_ (_03191_, _03077_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _54984_ (_03192_, _03191_, _03079_);
  or _54985_ (_03193_, _03192_, _03189_);
  or _54986_ (_03195_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _54987_ (_03196_, _03195_, _43634_);
  and _54988_ (_40545_, _03196_, _03193_);
  nor _54989_ (_03198_, _03090_, _39306_);
  and _54990_ (_03199_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  or _54991_ (_03200_, _03199_, _03079_);
  or _54992_ (_03202_, _03200_, _03198_);
  or _54993_ (_03203_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _54994_ (_03204_, _03203_, _43634_);
  and _54995_ (_40546_, _03204_, _03202_);
  nor _54996_ (_03206_, _03090_, _39298_);
  and _54997_ (_03207_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _54998_ (_03209_, _03207_, _03079_);
  or _54999_ (_03210_, _03209_, _03206_);
  or _55000_ (_03211_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _55001_ (_03213_, _03211_, _43634_);
  and _55002_ (_40547_, _03213_, _03210_);
  nor _55003_ (_03214_, _03090_, _39291_);
  and _55004_ (_03216_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _55005_ (_03217_, _03216_, _03079_);
  or _55006_ (_03218_, _03217_, _03214_);
  or _55007_ (_03220_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _55008_ (_03221_, _03220_, _43634_);
  and _55009_ (_40548_, _03221_, _03218_);
  nor _55010_ (_03223_, _03090_, _39284_);
  and _55011_ (_03224_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _55012_ (_03226_, _03224_, _03079_);
  or _55013_ (_03227_, _03226_, _03223_);
  or _55014_ (_03228_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _55015_ (_03229_, _03228_, _43634_);
  and _55016_ (_40550_, _03229_, _03227_);
  nor _55017_ (_03231_, _03090_, _39276_);
  and _55018_ (_03232_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _55019_ (_03234_, _03232_, _03079_);
  or _55020_ (_03235_, _03234_, _03231_);
  or _55021_ (_03236_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _55022_ (_03238_, _03236_, _43634_);
  and _55023_ (_40551_, _03238_, _03235_);
  nor _55024_ (_03239_, _03090_, _39268_);
  and _55025_ (_03241_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _55026_ (_03242_, _03241_, _03079_);
  or _55027_ (_03243_, _03242_, _03239_);
  or _55028_ (_03245_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _55029_ (_03246_, _03245_, _43634_);
  and _55030_ (_40552_, _03246_, _03243_);
  nor _55031_ (_03248_, _03090_, _39261_);
  and _55032_ (_03249_, _03090_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _55033_ (_03250_, _03249_, _03079_);
  or _55034_ (_03252_, _03250_, _03248_);
  or _55035_ (_03253_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _55036_ (_03255_, _03253_, _43634_);
  and _55037_ (_40553_, _03255_, _03252_);
  not _55038_ (_03256_, _03100_);
  and _55039_ (_03257_, _03256_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _55040_ (_03259_, _03256_, _39306_);
  or _55041_ (_03260_, _03259_, _03079_);
  or _55042_ (_03261_, _03260_, _03257_);
  or _55043_ (_03263_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _55044_ (_03264_, _03263_, _43634_);
  and _55045_ (_40554_, _03264_, _03261_);
  nor _55046_ (_03266_, _03256_, _39298_);
  and _55047_ (_03267_, _03256_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _55048_ (_03268_, _03267_, _03079_);
  or _55049_ (_03270_, _03268_, _03266_);
  or _55050_ (_03271_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _55051_ (_03272_, _03271_, _43634_);
  and _55052_ (_40555_, _03272_, _03270_);
  and _55053_ (_03274_, _03103_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _55054_ (_03275_, _03103_, _39291_);
  or _55055_ (_03277_, _03275_, _03274_);
  and _55056_ (_40556_, _03277_, _43634_);
  nor _55057_ (_03278_, _03256_, _39284_);
  and _55058_ (_03280_, _03256_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _55059_ (_03281_, _03280_, _03079_);
  or _55060_ (_03282_, _03281_, _03278_);
  or _55061_ (_03283_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _55062_ (_03284_, _03283_, _43634_);
  and _55063_ (_40557_, _03284_, _03282_);
  nor _55064_ (_03285_, _03256_, _39276_);
  and _55065_ (_03286_, _03256_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _55066_ (_03287_, _03286_, _03079_);
  or _55067_ (_03288_, _03287_, _03285_);
  or _55068_ (_03289_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _55069_ (_03290_, _03289_, _43634_);
  and _55070_ (_40558_, _03290_, _03288_);
  and _55071_ (_03291_, _03103_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _55072_ (_03292_, _03103_, _39268_);
  or _55073_ (_03293_, _03292_, _03291_);
  and _55074_ (_40559_, _03293_, _43634_);
  nor _55075_ (_03294_, _03256_, _39261_);
  and _55076_ (_03295_, _03256_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _55077_ (_03296_, _03295_, _03079_);
  or _55078_ (_03297_, _03296_, _03294_);
  or _55079_ (_03298_, _43100_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _55080_ (_03299_, _03298_, _43634_);
  and _55081_ (_40561_, _03299_, _03297_);
  not _55082_ (_03300_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _55083_ (_03301_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _55084_ (_03302_, _03301_, _03300_);
  and _55085_ (_03303_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _43634_);
  and _55086_ (_40590_, _03303_, _03302_);
  nor _55087_ (_03304_, _03302_, rst);
  nand _55088_ (_03305_, _03301_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _55089_ (_03306_, _03301_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _55090_ (_03307_, _03306_, _03305_);
  and _55091_ (_40592_, _03307_, _03304_);
  nor _55092_ (_03308_, _43450_, _43203_);
  nor _55093_ (_03309_, _43326_, _43243_);
  and _55094_ (_03310_, _03309_, _43404_);
  and _55095_ (_03311_, _03310_, _03308_);
  not _55096_ (_03312_, _43161_);
  nor _55097_ (_03313_, _40033_, _40022_);
  and _55098_ (_03314_, _40033_, _40022_);
  nor _55099_ (_03315_, _03314_, _03313_);
  nor _55100_ (_03316_, _40044_, _39947_);
  and _55101_ (_03317_, _40044_, _39947_);
  nor _55102_ (_03318_, _03317_, _03316_);
  and _55103_ (_03319_, _03318_, _03315_);
  nor _55104_ (_03320_, _03318_, _03315_);
  or _55105_ (_03321_, _03320_, _03319_);
  and _55106_ (_03322_, _39985_, _39967_);
  nor _55107_ (_03323_, _39985_, _39967_);
  or _55108_ (_03324_, _03323_, _03322_);
  not _55109_ (_03325_, _03324_);
  nor _55110_ (_03326_, _40011_, _39999_);
  and _55111_ (_03327_, _40011_, _39999_);
  or _55112_ (_03328_, _03327_, _03326_);
  and _55113_ (_03329_, _03328_, _03325_);
  nor _55114_ (_03330_, _03328_, _03325_);
  nor _55115_ (_03331_, _03330_, _03329_);
  or _55116_ (_03332_, _03331_, _03321_);
  nand _55117_ (_03333_, _03331_, _03321_);
  and _55118_ (_03334_, _03333_, _03332_);
  or _55119_ (_03335_, _03334_, _03312_);
  and _55120_ (_03336_, _43365_, _43285_);
  or _55121_ (_03337_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _55122_ (_03338_, _03337_, _03336_);
  and _55123_ (_03339_, _03338_, _03335_);
  not _55124_ (_03340_, _43285_);
  nor _55125_ (_03341_, _43365_, _03340_);
  and _55126_ (_03342_, _03341_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor _55127_ (_03343_, _43365_, _43285_);
  and _55128_ (_03344_, _03343_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _55129_ (_03345_, _03344_, _03342_);
  and _55130_ (_03346_, _03345_, _03312_);
  and _55131_ (_03348_, _43365_, _03340_);
  nor _55132_ (_03349_, _43161_, _34781_);
  and _55133_ (_03350_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _55134_ (_03351_, _03350_, _03349_);
  and _55135_ (_03352_, _03351_, _03348_);
  and _55136_ (_03353_, _03341_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _55137_ (_03354_, _03343_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _55138_ (_03355_, _03354_, _03353_);
  and _55139_ (_03356_, _03355_, _43161_);
  or _55140_ (_03357_, _03356_, _03352_);
  or _55141_ (_03358_, _03357_, _03346_);
  or _55142_ (_03359_, _03358_, _03339_);
  and _55143_ (_03360_, _03359_, _03311_);
  not _55144_ (_03361_, _43243_);
  and _55145_ (_03362_, _43326_, _03361_);
  and _55146_ (_03363_, _43450_, _43202_);
  or _55147_ (_03364_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _55148_ (_03365_, _43161_, _41477_);
  and _55149_ (_03366_, _03365_, _03336_);
  and _55150_ (_03367_, _03366_, _03364_);
  or _55151_ (_03368_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _55152_ (_03369_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _55153_ (_03370_, _03369_, _03343_);
  and _55154_ (_03371_, _03370_, _03368_);
  or _55155_ (_03372_, _03371_, _03367_);
  and _55156_ (_03373_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _55157_ (_03374_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _55158_ (_03375_, _03374_, _03373_);
  and _55159_ (_03376_, _03375_, _03341_);
  or _55160_ (_03377_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _55161_ (_03378_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _55162_ (_03379_, _03378_, _03348_);
  and _55163_ (_03380_, _03379_, _03377_);
  or _55164_ (_03381_, _03380_, _03376_);
  or _55165_ (_03382_, _03381_, _03372_);
  and _55166_ (_03383_, _03382_, _03363_);
  and _55167_ (_03384_, _43450_, _43203_);
  and _55168_ (_03385_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _55169_ (_03386_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _55170_ (_03387_, _03386_, _03385_);
  and _55171_ (_03388_, _03387_, _03343_);
  or _55172_ (_03389_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _55173_ (_03390_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _55174_ (_03391_, _03390_, _03336_);
  and _55175_ (_03392_, _03391_, _03389_);
  or _55176_ (_03393_, _03392_, _03388_);
  and _55177_ (_03394_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _55178_ (_03395_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _55179_ (_03396_, _03395_, _03394_);
  and _55180_ (_03397_, _03396_, _03348_);
  or _55181_ (_03398_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _55182_ (_03399_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _55183_ (_03400_, _03399_, _03341_);
  and _55184_ (_03401_, _03400_, _03398_);
  or _55185_ (_03402_, _03401_, _03397_);
  or _55186_ (_03403_, _03402_, _03393_);
  and _55187_ (_03404_, _03403_, _03384_);
  or _55188_ (_03405_, _03404_, _03383_);
  and _55189_ (_03406_, _03405_, _03362_);
  or _55190_ (_03407_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _55191_ (_03408_, _43161_, _41654_);
  and _55192_ (_03409_, _03408_, _03343_);
  and _55193_ (_03410_, _03409_, _03407_);
  and _55194_ (_03411_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _55195_ (_03412_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _55196_ (_03413_, _03412_, _03411_);
  and _55197_ (_03414_, _03413_, _03348_);
  or _55198_ (_03415_, _03414_, _03410_);
  and _55199_ (_03416_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor _55200_ (_03417_, _43161_, _41639_);
  or _55201_ (_03418_, _03417_, _03416_);
  and _55202_ (_03419_, _03418_, _03336_);
  and _55203_ (_03420_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _55204_ (_03421_, _43161_, _41643_);
  or _55205_ (_03422_, _03421_, _03420_);
  and _55206_ (_03423_, _03422_, _03341_);
  or _55207_ (_03424_, _03423_, _03419_);
  or _55208_ (_03425_, _03424_, _03415_);
  and _55209_ (_03426_, _03425_, _03384_);
  and _55210_ (_03427_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _55211_ (_03428_, _43161_, _42096_);
  or _55212_ (_03429_, _03428_, _03427_);
  and _55213_ (_03430_, _03429_, _03343_);
  and _55214_ (_03431_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _55215_ (_03432_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _55216_ (_03433_, _03432_, _03431_);
  and _55217_ (_03434_, _03433_, _03348_);
  or _55218_ (_03435_, _03434_, _03430_);
  and _55219_ (_03436_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _55220_ (_03437_, _43161_, _42113_);
  or _55221_ (_03438_, _03437_, _03436_);
  and _55222_ (_03439_, _03438_, _03336_);
  and _55223_ (_03440_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _55224_ (_03441_, _43161_, _42520_);
  or _55225_ (_03442_, _03441_, _03440_);
  and _55226_ (_03443_, _03442_, _03341_);
  or _55227_ (_03444_, _03443_, _03439_);
  or _55228_ (_03445_, _03444_, _03435_);
  and _55229_ (_03446_, _03445_, _03363_);
  or _55230_ (_03447_, _03446_, _03426_);
  and _55231_ (_03448_, _03447_, _03309_);
  and _55232_ (_03449_, _03362_, _03308_);
  and _55233_ (_03450_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _55234_ (_03451_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _55235_ (_03452_, _03451_, _03450_);
  and _55236_ (_03453_, _03452_, _03312_);
  and _55237_ (_03454_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _55238_ (_03455_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _55239_ (_03456_, _03455_, _03454_);
  and _55240_ (_03457_, _03456_, _03343_);
  and _55241_ (_03458_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nor _55242_ (_03459_, _43161_, _42093_);
  or _55243_ (_03460_, _03459_, _03458_);
  and _55244_ (_03461_, _03460_, _03341_);
  or _55245_ (_03462_, _03461_, _03457_);
  and _55246_ (_03463_, _03336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _55247_ (_03464_, _03348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _55248_ (_03465_, _03464_, _03463_);
  and _55249_ (_03466_, _03465_, _43161_);
  or _55250_ (_03467_, _03466_, _03462_);
  or _55251_ (_03468_, _03467_, _03453_);
  and _55252_ (_03469_, _03468_, _03449_);
  or _55253_ (_03470_, _03469_, _03448_);
  or _55254_ (_03471_, _03470_, _03406_);
  and _55255_ (_03472_, _03471_, _43405_);
  and _55256_ (_03473_, _39115_, _38590_);
  nor _55257_ (_03474_, _03473_, _39167_);
  and _55258_ (_03475_, _03474_, _00940_);
  and _55259_ (_03476_, _03475_, _01045_);
  nor _55260_ (_03477_, _39170_, _39163_);
  and _55261_ (_03478_, _39185_, _39086_);
  not _55262_ (_03479_, _03478_);
  and _55263_ (_03480_, _03479_, _03477_);
  and _55264_ (_03481_, _03480_, _00874_);
  and _55265_ (_03482_, _03481_, _01212_);
  and _55266_ (_03483_, _03482_, _03476_);
  and _55267_ (_03484_, _03483_, _39139_);
  nor _55268_ (_03485_, _03484_, _37633_);
  and _55269_ (_03486_, _01446_, p1in_reg[0]);
  and _55270_ (_03487_, _01442_, p1_in[0]);
  or _55271_ (_03488_, _03487_, _03486_);
  or _55272_ (_03489_, _03488_, _03485_);
  not _55273_ (_03490_, _03485_);
  or _55274_ (_03491_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _55275_ (_03492_, _03491_, _03489_);
  or _55276_ (_03493_, _03492_, _03312_);
  and _55277_ (_03494_, _01446_, p1in_reg[4]);
  and _55278_ (_03495_, _01442_, p1_in[4]);
  or _55279_ (_03496_, _03495_, _03494_);
  or _55280_ (_03497_, _03496_, _03485_);
  or _55281_ (_03498_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _55282_ (_03499_, _03498_, _03497_);
  or _55283_ (_03500_, _03499_, _43161_);
  and _55284_ (_03501_, _03500_, _03336_);
  and _55285_ (_03502_, _03501_, _03493_);
  and _55286_ (_03503_, _01446_, p1in_reg[3]);
  and _55287_ (_03504_, _01442_, p1_in[3]);
  or _55288_ (_03505_, _03504_, _03503_);
  or _55289_ (_03506_, _03505_, _03485_);
  or _55290_ (_03507_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _55291_ (_03508_, _03507_, _03506_);
  or _55292_ (_03509_, _03508_, _03312_);
  and _55293_ (_03510_, _01446_, p1in_reg[7]);
  and _55294_ (_03511_, _01442_, p1_in[7]);
  or _55295_ (_03512_, _03511_, _03510_);
  or _55296_ (_03513_, _03512_, _03485_);
  or _55297_ (_03514_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _55298_ (_03515_, _03514_, _03513_);
  or _55299_ (_03516_, _03515_, _43161_);
  and _55300_ (_03517_, _03516_, _03343_);
  and _55301_ (_03518_, _03517_, _03509_);
  or _55302_ (_03519_, _03518_, _03502_);
  and _55303_ (_03520_, _01446_, p1in_reg[5]);
  and _55304_ (_03521_, _01442_, p1_in[5]);
  or _55305_ (_03522_, _03521_, _03520_);
  or _55306_ (_03523_, _03522_, _03485_);
  or _55307_ (_03524_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _55308_ (_03525_, _03524_, _03523_);
  and _55309_ (_03526_, _03525_, _03312_);
  and _55310_ (_03527_, _01446_, p1in_reg[1]);
  and _55311_ (_03528_, _01442_, p1_in[1]);
  or _55312_ (_03529_, _03528_, _03527_);
  or _55313_ (_03530_, _03529_, _03485_);
  or _55314_ (_03531_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _55315_ (_03532_, _03531_, _03530_);
  and _55316_ (_03533_, _03532_, _43161_);
  or _55317_ (_03534_, _03533_, _03526_);
  and _55318_ (_03535_, _03534_, _03341_);
  and _55319_ (_03536_, _01446_, p1in_reg[2]);
  and _55320_ (_03537_, _01442_, p1_in[2]);
  or _55321_ (_03538_, _03537_, _03536_);
  or _55322_ (_03539_, _03538_, _03485_);
  or _55323_ (_03540_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _55324_ (_03541_, _03540_, _03539_);
  or _55325_ (_03542_, _03541_, _03312_);
  and _55326_ (_03543_, _01446_, p1in_reg[6]);
  and _55327_ (_03544_, _01442_, p1_in[6]);
  or _55328_ (_03545_, _03544_, _03543_);
  or _55329_ (_03546_, _03545_, _03485_);
  or _55330_ (_03547_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _55331_ (_03549_, _03547_, _03546_);
  or _55332_ (_03550_, _03549_, _43161_);
  and _55333_ (_03551_, _03550_, _03348_);
  and _55334_ (_03552_, _03551_, _03542_);
  or _55335_ (_03553_, _03552_, _03535_);
  or _55336_ (_03554_, _03553_, _03519_);
  and _55337_ (_03555_, _03554_, _03310_);
  and _55338_ (_03556_, _03362_, _43404_);
  and _55339_ (_03557_, _01446_, p0in_reg[0]);
  and _55340_ (_03558_, _01442_, p0_in[0]);
  or _55341_ (_03559_, _03558_, _03557_);
  or _55342_ (_03560_, _03559_, _03485_);
  or _55343_ (_03561_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _55344_ (_03562_, _03561_, _03560_);
  or _55345_ (_03563_, _03562_, _03312_);
  and _55346_ (_03564_, _01446_, p0in_reg[4]);
  and _55347_ (_03565_, _01442_, p0_in[4]);
  or _55348_ (_03566_, _03565_, _03564_);
  or _55349_ (_03567_, _03566_, _03485_);
  or _55350_ (_03568_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _55351_ (_03569_, _03568_, _03567_);
  or _55352_ (_03570_, _03569_, _43161_);
  and _55353_ (_03571_, _03570_, _03336_);
  and _55354_ (_03572_, _03571_, _03563_);
  and _55355_ (_03573_, _01446_, p0in_reg[3]);
  and _55356_ (_03574_, _01442_, p0_in[3]);
  or _55357_ (_03575_, _03574_, _03573_);
  or _55358_ (_03576_, _03575_, _03485_);
  or _55359_ (_03577_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _55360_ (_03578_, _03577_, _03576_);
  or _55361_ (_03579_, _03578_, _03312_);
  and _55362_ (_03580_, _01446_, p0in_reg[7]);
  and _55363_ (_03581_, _01442_, p0_in[7]);
  or _55364_ (_03582_, _03581_, _03580_);
  or _55365_ (_03583_, _03582_, _03485_);
  or _55366_ (_03584_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _55367_ (_03585_, _03584_, _03583_);
  or _55368_ (_03586_, _03585_, _43161_);
  and _55369_ (_03587_, _03586_, _03343_);
  and _55370_ (_03588_, _03587_, _03579_);
  or _55371_ (_03589_, _03588_, _03572_);
  and _55372_ (_03590_, _01446_, p0in_reg[5]);
  and _55373_ (_03591_, _01442_, p0_in[5]);
  or _55374_ (_03592_, _03591_, _03590_);
  or _55375_ (_03593_, _03592_, _03485_);
  or _55376_ (_03594_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _55377_ (_03595_, _03594_, _03593_);
  and _55378_ (_03596_, _03595_, _03312_);
  and _55379_ (_03597_, _01446_, p0in_reg[1]);
  and _55380_ (_03598_, _01442_, p0_in[1]);
  or _55381_ (_03599_, _03598_, _03597_);
  or _55382_ (_03600_, _03599_, _03485_);
  or _55383_ (_03601_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _55384_ (_03602_, _03601_, _03600_);
  and _55385_ (_03603_, _03602_, _43161_);
  or _55386_ (_03604_, _03603_, _03596_);
  and _55387_ (_03605_, _03604_, _03341_);
  and _55388_ (_03606_, _01446_, p0in_reg[2]);
  and _55389_ (_03607_, _01442_, p0_in[2]);
  or _55390_ (_03608_, _03607_, _03606_);
  or _55391_ (_03609_, _03608_, _03485_);
  nand _55392_ (_03610_, _03485_, _40328_);
  and _55393_ (_03611_, _03610_, _03609_);
  or _55394_ (_03612_, _03611_, _03312_);
  and _55395_ (_03613_, _01446_, p0in_reg[6]);
  and _55396_ (_03614_, _01442_, p0_in[6]);
  or _55397_ (_03615_, _03614_, _03613_);
  or _55398_ (_03616_, _03615_, _03485_);
  or _55399_ (_03617_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _55400_ (_03618_, _03617_, _03616_);
  or _55401_ (_03619_, _03618_, _43161_);
  and _55402_ (_03620_, _03619_, _03348_);
  and _55403_ (_03621_, _03620_, _03612_);
  or _55404_ (_03622_, _03621_, _03605_);
  or _55405_ (_03623_, _03622_, _03589_);
  and _55406_ (_03624_, _03623_, _03556_);
  or _55407_ (_03625_, _03624_, _03555_);
  and _55408_ (_03626_, _03625_, _03363_);
  and _55409_ (_03627_, _01446_, p3in_reg[3]);
  and _55410_ (_03628_, _01442_, p3_in[3]);
  or _55411_ (_03629_, _03628_, _03627_);
  or _55412_ (_03630_, _03629_, _03485_);
  or _55413_ (_03631_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _55414_ (_03632_, _03631_, _03630_);
  or _55415_ (_03633_, _03632_, _03312_);
  and _55416_ (_03634_, _01446_, p3in_reg[7]);
  and _55417_ (_03635_, _01442_, p3_in[7]);
  or _55418_ (_03636_, _03635_, _03634_);
  or _55419_ (_03637_, _03636_, _03485_);
  or _55420_ (_03638_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _55421_ (_03639_, _03638_, _03637_);
  or _55422_ (_03640_, _03639_, _43161_);
  and _55423_ (_03641_, _03640_, _03343_);
  and _55424_ (_03642_, _03641_, _03633_);
  and _55425_ (_03643_, _01446_, p3in_reg[5]);
  and _55426_ (_03644_, _01442_, p3_in[5]);
  or _55427_ (_03645_, _03644_, _03643_);
  or _55428_ (_03646_, _03645_, _03485_);
  or _55429_ (_03647_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _55430_ (_03648_, _03647_, _03646_);
  and _55431_ (_03649_, _03648_, _03312_);
  and _55432_ (_03650_, _01446_, p3in_reg[1]);
  and _55433_ (_03651_, _01442_, p3_in[1]);
  or _55434_ (_03652_, _03651_, _03650_);
  or _55435_ (_03653_, _03652_, _03485_);
  or _55436_ (_03654_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _55437_ (_03655_, _03654_, _03653_);
  and _55438_ (_03656_, _03655_, _43161_);
  or _55439_ (_03657_, _03656_, _03649_);
  and _55440_ (_03658_, _03657_, _03341_);
  or _55441_ (_03659_, _03658_, _03642_);
  and _55442_ (_03660_, _01446_, p3in_reg[0]);
  and _55443_ (_03661_, _01442_, p3_in[0]);
  or _55444_ (_03662_, _03661_, _03660_);
  or _55445_ (_03663_, _03662_, _03485_);
  or _55446_ (_03664_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _55447_ (_03665_, _03664_, _03663_);
  or _55448_ (_03666_, _03665_, _03312_);
  and _55449_ (_03667_, _01446_, p3in_reg[4]);
  and _55450_ (_03668_, _01442_, p3_in[4]);
  or _55451_ (_03669_, _03668_, _03667_);
  or _55452_ (_03670_, _03669_, _03485_);
  or _55453_ (_03671_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _55454_ (_03672_, _03671_, _03670_);
  or _55455_ (_03673_, _03672_, _43161_);
  and _55456_ (_03674_, _03673_, _03336_);
  and _55457_ (_03675_, _03674_, _03666_);
  and _55458_ (_03676_, _01446_, p3in_reg[6]);
  and _55459_ (_03677_, _01442_, p3_in[6]);
  or _55460_ (_03678_, _03677_, _03676_);
  or _55461_ (_03679_, _03678_, _03485_);
  or _55462_ (_03680_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _55463_ (_03681_, _03680_, _03679_);
  and _55464_ (_03682_, _03681_, _03312_);
  and _55465_ (_03683_, _01446_, p3in_reg[2]);
  and _55466_ (_03684_, _01442_, p3_in[2]);
  or _55467_ (_03685_, _03684_, _03683_);
  or _55468_ (_03686_, _03685_, _03485_);
  or _55469_ (_03687_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _55470_ (_03688_, _03687_, _03686_);
  and _55471_ (_03689_, _03688_, _43161_);
  or _55472_ (_03690_, _03689_, _03682_);
  and _55473_ (_03691_, _03690_, _03348_);
  or _55474_ (_03692_, _03691_, _03675_);
  or _55475_ (_03693_, _03692_, _03659_);
  and _55476_ (_03694_, _03693_, _03384_);
  nor _55477_ (_03695_, _43450_, _43202_);
  and _55478_ (_03696_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _55479_ (_03697_, _43161_, _31897_);
  or _55480_ (_03698_, _03697_, _03696_);
  and _55481_ (_03699_, _03698_, _03343_);
  nor _55482_ (_03700_, _43161_, _37436_);
  and _55483_ (_03701_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _55484_ (_03702_, _03701_, _03700_);
  and _55485_ (_03703_, _03702_, _03348_);
  or _55486_ (_03704_, _03703_, _03699_);
  and _55487_ (_03705_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor _55488_ (_03706_, _43161_, _35913_);
  or _55489_ (_03707_, _03706_, _03705_);
  and _55490_ (_03708_, _03707_, _03336_);
  and _55491_ (_03709_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _55492_ (_03710_, _43161_, _36708_);
  or _55493_ (_03711_, _03710_, _03709_);
  and _55494_ (_03712_, _03711_, _03341_);
  or _55495_ (_03713_, _03712_, _03708_);
  or _55496_ (_03714_, _03713_, _03704_);
  and _55497_ (_03715_, _03714_, _03695_);
  or _55498_ (_03716_, _03715_, _03694_);
  and _55499_ (_03717_, _03716_, _03310_);
  and _55500_ (_03718_, _03695_, _03556_);
  or _55501_ (_03719_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _55502_ (_03720_, _43161_, _39970_);
  and _55503_ (_03721_, _03720_, _03341_);
  and _55504_ (_03722_, _03721_, _03719_);
  and _55505_ (_03723_, _03312_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _55506_ (_03724_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _55507_ (_03725_, _03724_, _03723_);
  and _55508_ (_03726_, _03725_, _03348_);
  or _55509_ (_03727_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _55510_ (_03728_, _43161_, _39951_);
  and _55511_ (_03729_, _03728_, _03336_);
  and _55512_ (_03730_, _03729_, _03727_);
  or _55513_ (_03731_, _43161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand _55514_ (_03732_, _43161_, _40002_);
  and _55515_ (_03733_, _03732_, _03343_);
  and _55516_ (_03734_, _03733_, _03731_);
  or _55517_ (_03735_, _03734_, _03730_);
  or _55518_ (_03736_, _03735_, _03726_);
  or _55519_ (_03737_, _03736_, _03722_);
  and _55520_ (_03738_, _03737_, _03718_);
  and _55521_ (_03739_, _01481_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _55522_ (_03740_, _43450_, _03361_);
  nand _55523_ (_03741_, _03740_, _43405_);
  nor _55524_ (_03742_, _03310_, _29785_);
  and _55525_ (_03743_, _03742_, _03741_);
  not _55526_ (_03744_, _03556_);
  or _55527_ (_03745_, _03744_, _03308_);
  nand _55528_ (_03746_, _03449_, _43405_);
  and _55529_ (_03747_, _03746_, _03745_);
  and _55530_ (_03748_, _03747_, _03743_);
  and _55531_ (_03750_, _03556_, _03384_);
  and _55532_ (_03751_, _01446_, p2in_reg[3]);
  and _55533_ (_03752_, _01442_, p2_in[3]);
  or _55534_ (_03753_, _03752_, _03751_);
  or _55535_ (_03754_, _03753_, _03485_);
  or _55536_ (_03755_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _55537_ (_03756_, _03755_, _03754_);
  or _55538_ (_03757_, _03756_, _03312_);
  and _55539_ (_03758_, _01446_, p2in_reg[7]);
  and _55540_ (_03759_, _01442_, p2_in[7]);
  or _55541_ (_03760_, _03759_, _03758_);
  or _55542_ (_03761_, _03760_, _03485_);
  or _55543_ (_03762_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _55544_ (_03763_, _03762_, _03761_);
  or _55545_ (_03764_, _03763_, _43161_);
  and _55546_ (_03765_, _03764_, _03343_);
  and _55547_ (_03766_, _03765_, _03757_);
  and _55548_ (_03767_, _01446_, p2in_reg[6]);
  and _55549_ (_03768_, _01442_, p2_in[6]);
  or _55550_ (_03769_, _03768_, _03767_);
  or _55551_ (_03770_, _03769_, _03485_);
  or _55552_ (_03771_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _55553_ (_03772_, _03771_, _03770_);
  and _55554_ (_03773_, _03772_, _03312_);
  and _55555_ (_03774_, _01446_, p2in_reg[2]);
  and _55556_ (_03775_, _01442_, p2_in[2]);
  or _55557_ (_03776_, _03775_, _03774_);
  or _55558_ (_03777_, _03776_, _03485_);
  or _55559_ (_03778_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _55560_ (_03779_, _03778_, _03777_);
  and _55561_ (_03780_, _03779_, _43161_);
  or _55562_ (_03781_, _03780_, _03773_);
  and _55563_ (_03782_, _03781_, _03348_);
  or _55564_ (_03783_, _03782_, _03766_);
  and _55565_ (_03784_, _01446_, p2in_reg[0]);
  and _55566_ (_03785_, _01442_, p2_in[0]);
  or _55567_ (_03786_, _03785_, _03784_);
  or _55568_ (_03787_, _03786_, _03485_);
  or _55569_ (_03788_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _55570_ (_03789_, _03788_, _03787_);
  or _55571_ (_03790_, _03789_, _03312_);
  and _55572_ (_03791_, _01446_, p2in_reg[4]);
  and _55573_ (_03792_, _01442_, p2_in[4]);
  or _55574_ (_03793_, _03792_, _03791_);
  or _55575_ (_03794_, _03793_, _03485_);
  or _55576_ (_03795_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _55577_ (_03796_, _03795_, _03794_);
  or _55578_ (_03797_, _03796_, _43161_);
  and _55579_ (_03798_, _03797_, _03336_);
  and _55580_ (_03799_, _03798_, _03790_);
  and _55581_ (_03800_, _01446_, p2in_reg[5]);
  and _55582_ (_03801_, _01442_, p2_in[5]);
  or _55583_ (_03802_, _03801_, _03800_);
  or _55584_ (_03803_, _03802_, _03485_);
  or _55585_ (_03804_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _55586_ (_03805_, _03804_, _03803_);
  and _55587_ (_03806_, _03805_, _03312_);
  and _55588_ (_03807_, _01446_, p2in_reg[1]);
  and _55589_ (_03808_, _01442_, p2_in[1]);
  or _55590_ (_03809_, _03808_, _03807_);
  or _55591_ (_03810_, _03809_, _03485_);
  or _55592_ (_03811_, _03490_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _55593_ (_03812_, _03811_, _03810_);
  and _55594_ (_03813_, _03812_, _43161_);
  or _55595_ (_03814_, _03813_, _03806_);
  and _55596_ (_03815_, _03814_, _03341_);
  or _55597_ (_03816_, _03815_, _03799_);
  or _55598_ (_03817_, _03816_, _03783_);
  and _55599_ (_03818_, _03817_, _03750_);
  or _55600_ (_03819_, _03818_, _03748_);
  or _55601_ (_03820_, _03819_, _03739_);
  or _55602_ (_03821_, _03820_, _03738_);
  or _55603_ (_03822_, _03821_, _03717_);
  or _55604_ (_03823_, _03822_, _03626_);
  or _55605_ (_03824_, _03823_, _03472_);
  or _55606_ (_03825_, _03824_, _03360_);
  and _55607_ (_03826_, _03718_, _39923_);
  nor _55608_ (_03827_, _03826_, _01487_);
  nand _55609_ (_03828_, _03739_, _32431_);
  and _55610_ (_03829_, _03828_, _03827_);
  and _55611_ (_03830_, _03829_, _03825_);
  nor _55612_ (_03831_, _43161_, _39268_);
  and _55613_ (_03832_, _43161_, _43256_);
  or _55614_ (_03833_, _03832_, _03831_);
  and _55615_ (_03834_, _03833_, _03341_);
  or _55616_ (_03835_, _43161_, _42899_);
  nand _55617_ (_03836_, _43161_, _39291_);
  and _55618_ (_03837_, _03836_, _03348_);
  and _55619_ (_03838_, _03837_, _03835_);
  nor _55620_ (_03839_, _43161_, _39327_);
  and _55621_ (_03840_, _43161_, _43367_);
  or _55622_ (_03841_, _03840_, _03839_);
  and _55623_ (_03842_, _03841_, _03343_);
  nand _55624_ (_03843_, _43161_, _39306_);
  or _55625_ (_03844_, _43161_, _43308_);
  and _55626_ (_03845_, _03844_, _03336_);
  and _55627_ (_03846_, _03845_, _03843_);
  or _55628_ (_03847_, _03846_, _03842_);
  or _55629_ (_03848_, _03847_, _03838_);
  nor _55630_ (_03849_, _03848_, _03834_);
  nor _55631_ (_03850_, _03849_, _03827_);
  or _55632_ (_03851_, _03850_, _03830_);
  and _55633_ (_40593_, _03851_, _43634_);
  and _55634_ (_03852_, _43326_, _43203_);
  nor _55635_ (_03853_, _43450_, _43243_);
  and _55636_ (_03854_, _43404_, _43161_);
  and _55637_ (_03855_, _03854_, _03336_);
  and _55638_ (_03856_, _03855_, _03853_);
  and _55639_ (_03857_, _03856_, _03852_);
  and _55640_ (_03858_, _03857_, _39923_);
  not _55641_ (_03859_, _39934_);
  and _55642_ (_03860_, _03343_, _03312_);
  nor _55643_ (_03861_, _03860_, _03859_);
  and _55644_ (_03862_, _03861_, _01468_);
  nor _55645_ (_03863_, _03862_, _03858_);
  and _55646_ (_03864_, _03863_, _01484_);
  and _55647_ (_03865_, _03363_, _03362_);
  and _55648_ (_03866_, _03854_, _03343_);
  and _55649_ (_03867_, _03866_, _03865_);
  and _55650_ (_03868_, _03867_, _39375_);
  not _55651_ (_03869_, _03868_);
  and _55652_ (_03870_, _03857_, _39920_);
  and _55653_ (_03871_, _43327_, _43202_);
  and _55654_ (_03872_, _03871_, _03856_);
  and _55655_ (_03873_, _03872_, _39754_);
  nor _55656_ (_03874_, _03873_, _03870_);
  and _55657_ (_03875_, _03874_, _03869_);
  nor _55658_ (_03876_, _03875_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _55659_ (_03877_, _03876_);
  and _55660_ (_03878_, _03877_, _03864_);
  and _55661_ (_03879_, _03865_, _03348_);
  and _55662_ (_03880_, _03879_, _03854_);
  and _55663_ (_03881_, _03880_, _39375_);
  or _55664_ (_03882_, _03881_, rst);
  nor _55665_ (_40594_, _03882_, _03878_);
  nand _55666_ (_03883_, _03881_, _31809_);
  and _55667_ (_03884_, _43405_, _43161_);
  and _55668_ (_03885_, _03884_, _03336_);
  and _55669_ (_03886_, _03885_, _03449_);
  and _55670_ (_03887_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _55671_ (_03888_, _43404_, _43161_);
  and _55672_ (_03889_, _03888_, _03336_);
  and _55673_ (_03890_, _03889_, _03449_);
  and _55674_ (_03891_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _55675_ (_03892_, _03891_, _03887_);
  and _55676_ (_03893_, _03884_, _03348_);
  and _55677_ (_03894_, _03893_, _03449_);
  and _55678_ (_03895_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _55679_ (_03896_, _03888_, _03341_);
  and _55680_ (_03897_, _03896_, _03449_);
  and _55681_ (_03898_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _55682_ (_03899_, _03898_, _03895_);
  or _55683_ (_03900_, _03899_, _03892_);
  and _55684_ (_03901_, _03884_, _03343_);
  and _55685_ (_03902_, _03901_, _03449_);
  and _55686_ (_03903_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _55687_ (_03904_, _03885_, _03865_);
  and _55688_ (_03905_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _55689_ (_03906_, _03905_, _03903_);
  and _55690_ (_03907_, _03384_, _03362_);
  and _55691_ (_03908_, _03907_, _03885_);
  and _55692_ (_03909_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _55693_ (_03910_, _03860_, _43404_);
  nor _55694_ (_03911_, _43326_, _43202_);
  and _55695_ (_03912_, _03911_, _03740_);
  and _55696_ (_03913_, _03912_, _03910_);
  and _55697_ (_03914_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _55698_ (_03915_, _03914_, _03909_);
  or _55699_ (_03916_, _03915_, _03906_);
  or _55700_ (_03917_, _03916_, _03900_);
  and _55701_ (_03918_, _03901_, _03865_);
  and _55702_ (_03919_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _55703_ (_03920_, _03884_, _03341_);
  and _55704_ (_03921_, _03920_, _03865_);
  and _55705_ (_03922_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _55706_ (_03923_, _03922_, _03919_);
  and _55707_ (_03924_, _03896_, _03865_);
  and _55708_ (_03925_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _55709_ (_03926_, _03893_, _03865_);
  and _55710_ (_03927_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _55711_ (_03928_, _03927_, _03925_);
  or _55712_ (_03929_, _03928_, _03923_);
  and _55713_ (_03930_, _03363_, _03309_);
  and _55714_ (_03931_, _03930_, _03920_);
  and _55715_ (_03932_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _55716_ (_03933_, _03885_, _03930_);
  and _55717_ (_03934_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _55718_ (_03935_, _03934_, _03932_);
  and _55719_ (_03936_, _03910_, _03865_);
  and _55720_ (_03937_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _55721_ (_03938_, _03889_, _03865_);
  and _55722_ (_03939_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _55723_ (_03940_, _03939_, _03937_);
  or _55724_ (_03941_, _03940_, _03935_);
  or _55725_ (_03942_, _03941_, _03929_);
  or _55726_ (_03943_, _03942_, _03917_);
  and _55727_ (_03944_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _55728_ (_03945_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _55729_ (_03946_, _03945_, _03944_);
  and _55730_ (_03947_, _03911_, _03856_);
  and _55731_ (_03949_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _55732_ (_03950_, _03854_, _03341_);
  and _55733_ (_03951_, _03950_, _03865_);
  and _55734_ (_03952_, _03951_, _39329_);
  or _55735_ (_03953_, _03952_, _03949_);
  or _55736_ (_03954_, _03953_, _03946_);
  and _55737_ (_03955_, _03912_, _03855_);
  and _55738_ (_03956_, _03955_, _03639_);
  and _55739_ (_03957_, _03907_, _03855_);
  and _55740_ (_03958_, _03957_, _03763_);
  or _55741_ (_03959_, _03958_, _03956_);
  and _55742_ (_03960_, _03865_, _03855_);
  and _55743_ (_03961_, _03960_, _03585_);
  and _55744_ (_03962_, _03930_, _03855_);
  and _55745_ (_03963_, _03962_, _03515_);
  or _55746_ (_03964_, _03963_, _03961_);
  or _55747_ (_03965_, _03964_, _03959_);
  or _55748_ (_03966_, _03965_, _03954_);
  and _55749_ (_03967_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _55750_ (_03968_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _55751_ (_03969_, _03968_, _03967_);
  or _55752_ (_03970_, _03969_, _03966_);
  or _55753_ (_03971_, _03970_, _03943_);
  and _55754_ (_03972_, _03971_, _03878_);
  not _55755_ (_03973_, _03878_);
  nor _55756_ (_03974_, _03890_, _03886_);
  nor _55757_ (_03975_, _03897_, _03894_);
  and _55758_ (_03976_, _03975_, _03974_);
  nor _55759_ (_03977_, _03904_, _03902_);
  nor _55760_ (_03978_, _03913_, _03908_);
  and _55761_ (_03979_, _03978_, _03977_);
  and _55762_ (_03980_, _03979_, _03976_);
  nor _55763_ (_03981_, _03921_, _03918_);
  nor _55764_ (_03982_, _03926_, _03924_);
  and _55765_ (_03983_, _03982_, _03981_);
  or _55766_ (_03984_, _03933_, _03931_);
  or _55767_ (_03985_, _03938_, _03936_);
  nor _55768_ (_03986_, _03985_, _03984_);
  and _55769_ (_03987_, _03986_, _03983_);
  and _55770_ (_03988_, _03987_, _03980_);
  nor _55771_ (_03989_, _03880_, _03867_);
  nor _55772_ (_03990_, _03951_, _03947_);
  and _55773_ (_03991_, _03990_, _03989_);
  nor _55774_ (_03992_, _03957_, _03955_);
  nor _55775_ (_03993_, _03962_, _03960_);
  and _55776_ (_03994_, _03993_, _03992_);
  and _55777_ (_03995_, _03994_, _03991_);
  nor _55778_ (_03996_, _03872_, _03857_);
  and _55779_ (_03997_, _03996_, _03995_);
  and _55780_ (_03998_, _03997_, _03988_);
  or _55781_ (_03999_, _03998_, _03973_);
  and _55782_ (_04000_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _55783_ (_04001_, _04000_, _03881_);
  or _55784_ (_04002_, _04001_, _03972_);
  and _55785_ (_04003_, _04002_, _43634_);
  and _55786_ (_40595_, _04003_, _03883_);
  nor _55787_ (_40672_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _55788_ (_04004_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _55789_ (_04005_, _03301_, rst);
  and _55790_ (_40673_, _04005_, _04004_);
  nor _55791_ (_04006_, _03301_, _03300_);
  or _55792_ (_04007_, _04006_, _03302_);
  and _55793_ (_04008_, _03305_, _43634_);
  and _55794_ (_40674_, _04008_, _04007_);
  and _55795_ (_04009_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _55796_ (_04010_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _55797_ (_04011_, _04010_, _04009_);
  and _55798_ (_04012_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _55799_ (_04013_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _55800_ (_04014_, _04013_, _04012_);
  or _55801_ (_04015_, _04014_, _04011_);
  and _55802_ (_04016_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _55803_ (_04017_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _55804_ (_04018_, _04017_, _04016_);
  and _55805_ (_04019_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _55806_ (_04020_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _55807_ (_04021_, _04020_, _04019_);
  or _55808_ (_04022_, _04021_, _04018_);
  or _55809_ (_04023_, _04022_, _04015_);
  and _55810_ (_04024_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _55811_ (_04025_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _55812_ (_04026_, _04025_, _04024_);
  and _55813_ (_04027_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _55814_ (_04028_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _55815_ (_04029_, _04028_, _04027_);
  or _55816_ (_04030_, _04029_, _04026_);
  and _55817_ (_04031_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _55818_ (_04032_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _55819_ (_04033_, _04032_, _04031_);
  and _55820_ (_04034_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _55821_ (_04035_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _55822_ (_04036_, _04035_, _04034_);
  or _55823_ (_04037_, _04036_, _04033_);
  or _55824_ (_04038_, _04037_, _04030_);
  or _55825_ (_04039_, _04038_, _04023_);
  and _55826_ (_04040_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _55827_ (_04041_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or _55828_ (_04042_, _04041_, _04040_);
  and _55829_ (_04043_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _55830_ (_04044_, _03951_, _43345_);
  or _55831_ (_04046_, _04044_, _04043_);
  or _55832_ (_04047_, _04046_, _04042_);
  and _55833_ (_04048_, _03955_, _03665_);
  and _55834_ (_04049_, _03957_, _03789_);
  or _55835_ (_04050_, _04049_, _04048_);
  and _55836_ (_04051_, _03962_, _03492_);
  and _55837_ (_04052_, _03960_, _03562_);
  or _55838_ (_04053_, _04052_, _04051_);
  or _55839_ (_04054_, _04053_, _04050_);
  or _55840_ (_04055_, _04054_, _04047_);
  and _55841_ (_04056_, _03872_, _03334_);
  and _55842_ (_04057_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _55843_ (_04058_, _04057_, _04056_);
  or _55844_ (_04059_, _04058_, _04055_);
  or _55845_ (_04060_, _04059_, _04039_);
  and _55846_ (_04061_, _04060_, _03878_);
  and _55847_ (_04062_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _55848_ (_04063_, _04062_, _03881_);
  or _55849_ (_04064_, _04063_, _04061_);
  nand _55850_ (_04065_, _03881_, _32953_);
  and _55851_ (_04066_, _04065_, _43634_);
  and _55852_ (_40675_, _04066_, _04064_);
  nand _55853_ (_04067_, _03881_, _33639_);
  and _55854_ (_04068_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _55855_ (_04069_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _55856_ (_04070_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _55857_ (_04071_, _04070_, _04069_);
  and _55858_ (_04072_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _55859_ (_04073_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _55860_ (_04074_, _04073_, _04072_);
  or _55861_ (_04075_, _04074_, _04071_);
  and _55862_ (_04076_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _55863_ (_04077_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _55864_ (_04078_, _04077_, _04076_);
  and _55865_ (_04079_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _55866_ (_04080_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _55867_ (_04081_, _04080_, _04079_);
  or _55868_ (_04082_, _04081_, _04078_);
  or _55869_ (_04083_, _04082_, _04075_);
  and _55870_ (_04084_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _55871_ (_04085_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _55872_ (_04086_, _04085_, _04084_);
  and _55873_ (_04087_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _55874_ (_04088_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _55875_ (_04089_, _04088_, _04087_);
  or _55876_ (_04090_, _04089_, _04086_);
  and _55877_ (_04091_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _55878_ (_04092_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _55879_ (_04093_, _04092_, _04091_);
  and _55880_ (_04094_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _55881_ (_04095_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _55882_ (_04096_, _04095_, _04094_);
  or _55883_ (_04097_, _04096_, _04093_);
  or _55884_ (_04098_, _04097_, _04090_);
  or _55885_ (_04099_, _04098_, _04083_);
  and _55886_ (_04100_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _55887_ (_04101_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _55888_ (_04102_, _04101_, _04100_);
  and _55889_ (_04103_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _55890_ (_04104_, _03951_, _43280_);
  or _55891_ (_04105_, _04104_, _04103_);
  or _55892_ (_04106_, _04105_, _04102_);
  and _55893_ (_04107_, _03955_, _03655_);
  and _55894_ (_04108_, _03957_, _03812_);
  or _55895_ (_04109_, _04108_, _04107_);
  and _55896_ (_04110_, _03962_, _03532_);
  and _55897_ (_04111_, _03960_, _03602_);
  or _55898_ (_04112_, _04111_, _04110_);
  or _55899_ (_04113_, _04112_, _04109_);
  or _55900_ (_04114_, _04113_, _04106_);
  and _55901_ (_04115_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _55902_ (_04116_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _55903_ (_04117_, _04116_, _04115_);
  or _55904_ (_04118_, _04117_, _04114_);
  or _55905_ (_04119_, _04118_, _04099_);
  and _55906_ (_04120_, _04119_, _03878_);
  or _55907_ (_04121_, _04120_, _04068_);
  or _55908_ (_04122_, _04121_, _03881_);
  and _55909_ (_04123_, _04122_, _43634_);
  and _55910_ (_40677_, _04123_, _04067_);
  nand _55911_ (_04124_, _03881_, _34378_);
  and _55912_ (_04125_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _55913_ (_04126_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _55914_ (_04127_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _55915_ (_04128_, _04127_, _04126_);
  and _55916_ (_04129_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _55917_ (_04130_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _55918_ (_04131_, _04130_, _04129_);
  or _55919_ (_04132_, _04131_, _04128_);
  and _55920_ (_04133_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _55921_ (_04134_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _55922_ (_04135_, _04134_, _04133_);
  and _55923_ (_04136_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _55924_ (_04137_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _55925_ (_04138_, _04137_, _04136_);
  or _55926_ (_04139_, _04138_, _04135_);
  or _55927_ (_04140_, _04139_, _04132_);
  and _55928_ (_04141_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _55929_ (_04142_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _55930_ (_04143_, _04142_, _04141_);
  and _55931_ (_04145_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _55932_ (_04146_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _55933_ (_04147_, _04146_, _04145_);
  or _55934_ (_04148_, _04147_, _04143_);
  and _55935_ (_04149_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _55936_ (_04150_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _55937_ (_04151_, _04150_, _04149_);
  and _55938_ (_04152_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _55939_ (_04153_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _55940_ (_04154_, _04153_, _04152_);
  or _55941_ (_04155_, _04154_, _04151_);
  or _55942_ (_04156_, _04155_, _04148_);
  or _55943_ (_04157_, _04156_, _04140_);
  and _55944_ (_04158_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _55945_ (_04159_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _55946_ (_04160_, _04159_, _04158_);
  and _55947_ (_04161_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _55948_ (_04162_, _03951_, _43132_);
  or _55949_ (_04163_, _04162_, _04161_);
  or _55950_ (_04164_, _04163_, _04160_);
  and _55951_ (_04165_, _03955_, _03688_);
  and _55952_ (_04166_, _03957_, _03779_);
  or _55953_ (_04167_, _04166_, _04165_);
  and _55954_ (_04168_, _03960_, _03611_);
  and _55955_ (_04169_, _03962_, _03541_);
  or _55956_ (_04170_, _04169_, _04168_);
  or _55957_ (_04171_, _04170_, _04167_);
  or _55958_ (_04172_, _04171_, _04164_);
  and _55959_ (_04173_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _55960_ (_04174_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _55961_ (_04175_, _04174_, _04173_);
  or _55962_ (_04176_, _04175_, _04172_);
  or _55963_ (_04177_, _04176_, _04157_);
  and _55964_ (_04178_, _04177_, _03878_);
  or _55965_ (_04179_, _04178_, _04125_);
  or _55966_ (_04180_, _04179_, _03881_);
  and _55967_ (_04181_, _04180_, _43634_);
  and _55968_ (_40678_, _04181_, _04124_);
  nand _55969_ (_04182_, _03881_, _35118_);
  and _55970_ (_04183_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _55971_ (_04184_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _55972_ (_04185_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _55973_ (_04186_, _04185_, _04184_);
  and _55974_ (_04187_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _55975_ (_04188_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _55976_ (_04189_, _04188_, _04187_);
  or _55977_ (_04190_, _04189_, _04186_);
  and _55978_ (_04191_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _55979_ (_04192_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _55980_ (_04193_, _04192_, _04191_);
  and _55981_ (_04194_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _55982_ (_04195_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _55983_ (_04196_, _04195_, _04194_);
  or _55984_ (_04197_, _04196_, _04193_);
  or _55985_ (_04198_, _04197_, _04190_);
  and _55986_ (_04199_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _55987_ (_04200_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _55988_ (_04201_, _04200_, _04199_);
  and _55989_ (_04202_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _55990_ (_04203_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _55991_ (_04204_, _04203_, _04202_);
  or _55992_ (_04205_, _04204_, _04201_);
  and _55993_ (_04206_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _55994_ (_04207_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _55995_ (_04208_, _04207_, _04206_);
  and _55996_ (_04209_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _55997_ (_04210_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _55998_ (_04211_, _04210_, _04209_);
  or _55999_ (_04212_, _04211_, _04208_);
  or _56000_ (_04213_, _04212_, _04205_);
  or _56001_ (_04214_, _04213_, _04198_);
  and _56002_ (_04215_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _56003_ (_04216_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or _56004_ (_04217_, _04216_, _04215_);
  and _56005_ (_04218_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _56006_ (_04219_, _03951_, _43381_);
  or _56007_ (_04220_, _04219_, _04218_);
  or _56008_ (_04221_, _04220_, _04217_);
  and _56009_ (_04222_, _03955_, _03632_);
  and _56010_ (_04223_, _03957_, _03756_);
  or _56011_ (_04224_, _04223_, _04222_);
  and _56012_ (_04225_, _03962_, _03508_);
  and _56013_ (_04226_, _03960_, _03578_);
  or _56014_ (_04227_, _04226_, _04225_);
  or _56015_ (_04228_, _04227_, _04224_);
  or _56016_ (_04229_, _04228_, _04221_);
  and _56017_ (_04230_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _56018_ (_04231_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _56019_ (_04232_, _04231_, _04230_);
  or _56020_ (_04233_, _04232_, _04229_);
  or _56021_ (_04234_, _04233_, _04214_);
  and _56022_ (_04235_, _04234_, _03878_);
  or _56023_ (_04236_, _04235_, _04183_);
  or _56024_ (_04237_, _04236_, _03881_);
  and _56025_ (_04238_, _04237_, _43634_);
  and _56026_ (_40679_, _04238_, _04182_);
  nand _56027_ (_04239_, _03881_, _35880_);
  and _56028_ (_04240_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _56029_ (_04241_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _56030_ (_04242_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _56031_ (_04244_, _04242_, _04241_);
  and _56032_ (_04245_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _56033_ (_04246_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _56034_ (_04247_, _04246_, _04245_);
  or _56035_ (_04248_, _04247_, _04244_);
  and _56036_ (_04249_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _56037_ (_04250_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _56038_ (_04251_, _04250_, _04249_);
  and _56039_ (_04252_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _56040_ (_04253_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _56041_ (_04254_, _04253_, _04252_);
  or _56042_ (_04255_, _04254_, _04251_);
  or _56043_ (_04256_, _04255_, _04248_);
  and _56044_ (_04257_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _56045_ (_04258_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _56046_ (_04259_, _04258_, _04257_);
  and _56047_ (_04260_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _56048_ (_04261_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _56049_ (_04262_, _04261_, _04260_);
  or _56050_ (_04263_, _04262_, _04259_);
  and _56051_ (_04264_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _56052_ (_04265_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _56053_ (_04266_, _04265_, _04264_);
  and _56054_ (_04267_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _56055_ (_04268_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _56056_ (_04269_, _04268_, _04267_);
  or _56057_ (_04270_, _04269_, _04266_);
  or _56058_ (_04271_, _04270_, _04263_);
  or _56059_ (_04272_, _04271_, _04256_);
  and _56060_ (_04273_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _56061_ (_04274_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _56062_ (_04275_, _04274_, _04273_);
  and _56063_ (_04276_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _56064_ (_04277_, _03951_, _43322_);
  or _56065_ (_04278_, _04277_, _04276_);
  or _56066_ (_04279_, _04278_, _04275_);
  and _56067_ (_04280_, _03955_, _03672_);
  and _56068_ (_04281_, _03957_, _03796_);
  or _56069_ (_04282_, _04281_, _04280_);
  and _56070_ (_04283_, _03962_, _03499_);
  and _56071_ (_04284_, _03960_, _03569_);
  or _56072_ (_04285_, _04284_, _04283_);
  or _56073_ (_04286_, _04285_, _04282_);
  or _56074_ (_04287_, _04286_, _04279_);
  and _56075_ (_04288_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _56076_ (_04289_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _56077_ (_04290_, _04289_, _04288_);
  or _56078_ (_04291_, _04290_, _04287_);
  or _56079_ (_04292_, _04291_, _04272_);
  and _56080_ (_04293_, _04292_, _03878_);
  or _56081_ (_04294_, _04293_, _04240_);
  or _56082_ (_04295_, _04294_, _03881_);
  and _56083_ (_04296_, _04295_, _43634_);
  and _56084_ (_40680_, _04296_, _04239_);
  and _56085_ (_04297_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _56086_ (_04298_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _56087_ (_04299_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _56088_ (_04300_, _04299_, _04298_);
  and _56089_ (_04301_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _56090_ (_04302_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _56091_ (_04303_, _04302_, _04301_);
  or _56092_ (_04304_, _04303_, _04300_);
  and _56093_ (_04305_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _56094_ (_04306_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _56095_ (_04307_, _04306_, _04305_);
  and _56096_ (_04308_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _56097_ (_04309_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _56098_ (_04310_, _04309_, _04308_);
  or _56099_ (_04311_, _04310_, _04307_);
  or _56100_ (_04312_, _04311_, _04304_);
  and _56101_ (_04313_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _56102_ (_04314_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _56103_ (_04315_, _04314_, _04313_);
  and _56104_ (_04316_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _56105_ (_04317_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _56106_ (_04318_, _04317_, _04316_);
  or _56107_ (_04319_, _04318_, _04315_);
  and _56108_ (_04320_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _56109_ (_04321_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _56110_ (_04322_, _04321_, _04320_);
  and _56111_ (_04323_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _56112_ (_04324_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _56113_ (_04325_, _04324_, _04323_);
  or _56114_ (_04326_, _04325_, _04322_);
  or _56115_ (_04327_, _04326_, _04319_);
  or _56116_ (_04328_, _04327_, _04312_);
  and _56117_ (_04329_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _56118_ (_04330_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _56119_ (_04331_, _04330_, _04329_);
  and _56120_ (_04332_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _56121_ (_04333_, _03951_, _43166_);
  or _56122_ (_04334_, _04333_, _04332_);
  or _56123_ (_04335_, _04334_, _04331_);
  and _56124_ (_04336_, _03955_, _03648_);
  and _56125_ (_04337_, _03957_, _03805_);
  or _56126_ (_04338_, _04337_, _04336_);
  and _56127_ (_04339_, _03960_, _03595_);
  and _56128_ (_04340_, _03962_, _03525_);
  or _56129_ (_04341_, _04340_, _04339_);
  or _56130_ (_04342_, _04341_, _04338_);
  or _56131_ (_04344_, _04342_, _04335_);
  and _56132_ (_04345_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _56133_ (_04346_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _56134_ (_04347_, _04346_, _04345_);
  or _56135_ (_04348_, _04347_, _04344_);
  or _56136_ (_04349_, _04348_, _04328_);
  or _56137_ (_04350_, _03864_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _56138_ (_04351_, _04350_, _03877_);
  and _56139_ (_04352_, _04351_, _04349_);
  or _56140_ (_04353_, _04352_, _04297_);
  or _56141_ (_04354_, _04353_, _03881_);
  nand _56142_ (_04355_, _03881_, _36675_);
  and _56143_ (_04356_, _04355_, _43634_);
  and _56144_ (_40681_, _04356_, _04354_);
  nand _56145_ (_04357_, _03881_, _37403_);
  and _56146_ (_04358_, _03999_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _56147_ (_04359_, _03886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _56148_ (_04360_, _03890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _56149_ (_04361_, _04360_, _04359_);
  and _56150_ (_04362_, _03897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _56151_ (_04363_, _03894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _56152_ (_04364_, _04363_, _04362_);
  or _56153_ (_04365_, _04364_, _04361_);
  and _56154_ (_04366_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _56155_ (_04367_, _03904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _56156_ (_04368_, _04367_, _04366_);
  and _56157_ (_04369_, _03908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _56158_ (_04370_, _03913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _56159_ (_04371_, _04370_, _04369_);
  or _56160_ (_04372_, _04371_, _04368_);
  or _56161_ (_04373_, _04372_, _04365_);
  and _56162_ (_04374_, _03926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _56163_ (_04375_, _03924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _56164_ (_04376_, _04375_, _04374_);
  and _56165_ (_04377_, _03921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _56166_ (_04378_, _03918_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _56167_ (_04379_, _04378_, _04377_);
  or _56168_ (_04380_, _04379_, _04376_);
  and _56169_ (_04381_, _03931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _56170_ (_04382_, _03933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _56171_ (_04383_, _04382_, _04381_);
  and _56172_ (_04384_, _03938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _56173_ (_04385_, _03936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _56174_ (_04386_, _04385_, _04384_);
  or _56175_ (_04387_, _04386_, _04383_);
  or _56176_ (_04388_, _04387_, _04380_);
  or _56177_ (_04389_, _04388_, _04373_);
  and _56178_ (_04390_, _03880_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _56179_ (_04391_, _03867_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _56180_ (_04392_, _04391_, _04390_);
  and _56181_ (_04393_, _03947_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _56182_ (_04394_, _03951_, _43415_);
  or _56183_ (_04395_, _04394_, _04393_);
  or _56184_ (_04396_, _04395_, _04392_);
  and _56185_ (_04397_, _03955_, _03681_);
  and _56186_ (_04398_, _03957_, _03772_);
  or _56187_ (_04399_, _04398_, _04397_);
  and _56188_ (_04400_, _03960_, _03618_);
  and _56189_ (_04401_, _03962_, _03549_);
  or _56190_ (_04402_, _04401_, _04400_);
  or _56191_ (_04403_, _04402_, _04399_);
  or _56192_ (_04404_, _04403_, _04396_);
  and _56193_ (_04405_, _03872_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _56194_ (_04406_, _03857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _56195_ (_04407_, _04406_, _04405_);
  or _56196_ (_04408_, _04407_, _04404_);
  or _56197_ (_04409_, _04408_, _04389_);
  and _56198_ (_04410_, _04409_, _03878_);
  or _56199_ (_04411_, _04410_, _04358_);
  or _56200_ (_04412_, _04411_, _03881_);
  and _56201_ (_04413_, _04412_, _43634_);
  and _56202_ (_40682_, _04413_, _04357_);
  and _56203_ (_40750_, _43564_, _43634_);
  nor _56204_ (_40754_, _43161_, rst);
  and _56205_ (_40776_, _43667_, _43634_);
  nor _56206_ (_40779_, _43365_, rst);
  nor _56207_ (_40780_, _43285_, rst);
  not _56208_ (_04414_, _00113_);
  nor _56209_ (_04415_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _56210_ (_04416_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _56211_ (_04417_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04416_);
  nor _56212_ (_04418_, _04417_, _04415_);
  nor _56213_ (_04419_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _56214_ (_04420_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04416_);
  nor _56215_ (_04421_, _04420_, _04419_);
  and _56216_ (_04422_, _04421_, _04418_);
  nor _56217_ (_04423_, _02314_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _56218_ (_04424_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04416_);
  nor _56219_ (_04425_, _04424_, _04423_);
  nor _56220_ (_04426_, _04425_, _04422_);
  and _56221_ (_04427_, _04425_, _04422_);
  or _56222_ (_04428_, _04427_, _04426_);
  not _56223_ (_04429_, _04427_);
  nor _56224_ (_04430_, _02332_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _56225_ (_04431_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04416_);
  or _56226_ (_04432_, _04431_, _04430_);
  and _56227_ (_04433_, _04432_, _04429_);
  nor _56228_ (_04434_, _04432_, _04429_);
  nor _56229_ (_04435_, _04434_, _04433_);
  not _56230_ (_04437_, _04435_);
  and _56231_ (_04438_, _04437_, _04428_);
  not _56232_ (_04439_, _04418_);
  nor _56233_ (_04440_, _04421_, _04439_);
  and _56234_ (_04441_, _04440_, _04438_);
  and _56235_ (_04442_, _04441_, _04414_);
  not _56236_ (_04443_, _00696_);
  nor _56237_ (_04444_, _04432_, _04428_);
  and _56238_ (_04445_, _04444_, _04440_);
  nor _56239_ (_04446_, _04421_, _04418_);
  and _56240_ (_04447_, _04446_, _04444_);
  nor _56241_ (_04448_, _04447_, _04445_);
  not _56242_ (_04449_, _04422_);
  and _56243_ (_04450_, _04444_, _04449_);
  and _56244_ (_04451_, _04450_, _04448_);
  and _56245_ (_04452_, _04451_, _04443_);
  not _56246_ (_04453_, _00072_);
  and _56247_ (_04454_, _04446_, _04438_);
  and _56248_ (_04455_, _04454_, _04453_);
  or _56249_ (_04456_, _04455_, _04452_);
  or _56250_ (_04457_, _04456_, _04442_);
  not _56251_ (_04458_, _00513_);
  and _56252_ (_04459_, _04421_, _04439_);
  and _56253_ (_04460_, _04435_, _04428_);
  and _56254_ (_04461_, _04460_, _04459_);
  and _56255_ (_04462_, _04461_, _04458_);
  not _56256_ (_04463_, _00472_);
  and _56257_ (_04464_, _04460_, _04440_);
  and _56258_ (_04465_, _04464_, _04463_);
  or _56259_ (_04466_, _04465_, _04462_);
  not _56260_ (_04467_, _00431_);
  and _56261_ (_04468_, _04460_, _04446_);
  and _56262_ (_04469_, _04468_, _04467_);
  not _56263_ (_04470_, _00175_);
  and _56264_ (_04471_, _04459_, _04438_);
  and _56265_ (_04472_, _04471_, _04470_);
  or _56266_ (_04473_, _04472_, _04469_);
  or _56267_ (_04474_, _04473_, _04466_);
  not _56268_ (_04475_, _00267_);
  nor _56269_ (_04476_, _04435_, _04428_);
  and _56270_ (_04477_, _04446_, _04476_);
  and _56271_ (_04478_, _04477_, _04475_);
  not _56272_ (_04479_, _00614_);
  and _56273_ (_04480_, _04447_, _04479_);
  not _56274_ (_04481_, _00308_);
  and _56275_ (_04482_, _04476_, _04440_);
  and _56276_ (_04483_, _04482_, _04481_);
  or _56277_ (_04484_, _04483_, _04480_);
  or _56278_ (_04485_, _04484_, _04478_);
  not _56279_ (_04486_, _00349_);
  and _56280_ (_04487_, _04459_, _04476_);
  and _56281_ (_04488_, _04487_, _04486_);
  not _56282_ (_04489_, _00226_);
  and _56283_ (_04490_, _04433_, _04422_);
  and _56284_ (_04491_, _04490_, _04489_);
  not _56285_ (_04492_, _00390_);
  and _56286_ (_04493_, _04432_, _04427_);
  and _56287_ (_04494_, _04493_, _04492_);
  not _56288_ (_04495_, _00031_);
  and _56289_ (_04496_, _04434_, _04495_);
  or _56290_ (_04497_, _04496_, _04494_);
  or _56291_ (_04498_, _04497_, _04491_);
  or _56292_ (_04499_, _04498_, _04488_);
  not _56293_ (_04500_, _00655_);
  and _56294_ (_04501_, _04445_, _04500_);
  not _56295_ (_04502_, _00557_);
  and _56296_ (_04503_, _04444_, _04422_);
  and _56297_ (_04504_, _04503_, _04502_);
  or _56298_ (_04505_, _04504_, _04501_);
  or _56299_ (_04506_, _04505_, _04499_);
  or _56300_ (_04507_, _04506_, _04485_);
  or _56301_ (_04508_, _04507_, _04474_);
  or _56302_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04508_, _04457_);
  and _56303_ (_04509_, _04451_, _04495_);
  and _56304_ (_04510_, _04441_, _04470_);
  and _56305_ (_04511_, _04454_, _04414_);
  or _56306_ (_04512_, _04511_, _04510_);
  or _56307_ (_04513_, _04512_, _04509_);
  and _56308_ (_04514_, _04461_, _04502_);
  and _56309_ (_04515_, _04464_, _04458_);
  or _56310_ (_04516_, _04515_, _04514_);
  and _56311_ (_04517_, _04468_, _04463_);
  and _56312_ (_04518_, _04471_, _04489_);
  or _56313_ (_04519_, _04518_, _04517_);
  or _56314_ (_04520_, _04519_, _04516_);
  and _56315_ (_04521_, _04477_, _04481_);
  and _56316_ (_04522_, _04445_, _04443_);
  and _56317_ (_04523_, _04503_, _04479_);
  or _56318_ (_04524_, _04523_, _04522_);
  or _56319_ (_04525_, _04524_, _04521_);
  and _56320_ (_04526_, _04487_, _04492_);
  and _56321_ (_04527_, _04490_, _04475_);
  and _56322_ (_04528_, _04493_, _04467_);
  and _56323_ (_04529_, _04434_, _04453_);
  or _56324_ (_04530_, _04529_, _04528_);
  or _56325_ (_04531_, _04530_, _04527_);
  or _56326_ (_04532_, _04531_, _04526_);
  and _56327_ (_04533_, _04447_, _04500_);
  and _56328_ (_04534_, _04482_, _04486_);
  or _56329_ (_04535_, _04534_, _04533_);
  or _56330_ (_04537_, _04535_, _04532_);
  or _56331_ (_04538_, _04537_, _04525_);
  or _56332_ (_04539_, _04538_, _04520_);
  or _56333_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04539_, _04513_);
  and _56334_ (_04540_, _04441_, _04489_);
  and _56335_ (_04541_, _04454_, _04470_);
  and _56336_ (_04542_, _04451_, _04453_);
  or _56337_ (_04543_, _04542_, _04541_);
  or _56338_ (_04544_, _04543_, _04540_);
  and _56339_ (_04545_, _04461_, _04479_);
  and _56340_ (_04546_, _04464_, _04502_);
  or _56341_ (_04547_, _04546_, _04545_);
  and _56342_ (_04548_, _04468_, _04458_);
  and _56343_ (_04549_, _04471_, _04475_);
  or _56344_ (_04550_, _04549_, _04548_);
  or _56345_ (_04551_, _04550_, _04547_);
  and _56346_ (_04552_, _04482_, _04492_);
  and _56347_ (_04553_, _04477_, _04486_);
  or _56348_ (_04554_, _04553_, _04552_);
  and _56349_ (_04555_, _04487_, _04467_);
  or _56350_ (_04556_, _04555_, _04554_);
  and _56351_ (_04557_, _04447_, _04443_);
  and _56352_ (_04558_, _04490_, _04481_);
  and _56353_ (_04559_, _04493_, _04463_);
  and _56354_ (_04560_, _04434_, _04414_);
  or _56355_ (_04561_, _04560_, _04559_);
  or _56356_ (_04562_, _04561_, _04558_);
  or _56357_ (_04563_, _04562_, _04557_);
  and _56358_ (_04564_, _04503_, _04500_);
  and _56359_ (_04565_, _04445_, _04495_);
  or _56360_ (_04566_, _04565_, _04564_);
  or _56361_ (_04567_, _04566_, _04563_);
  or _56362_ (_04568_, _04567_, _04556_);
  or _56363_ (_04569_, _04568_, _04551_);
  or _56364_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04569_, _04544_);
  and _56365_ (_04570_, _04441_, _04453_);
  and _56366_ (_04571_, _04451_, _04500_);
  and _56367_ (_04572_, _04454_, _04495_);
  or _56368_ (_04573_, _04572_, _04571_);
  or _56369_ (_04574_, _04573_, _04570_);
  and _56370_ (_04575_, _04464_, _04467_);
  and _56371_ (_04576_, _04471_, _04414_);
  or _56372_ (_04577_, _04576_, _04575_);
  and _56373_ (_04578_, _04461_, _04463_);
  and _56374_ (_04579_, _04468_, _04492_);
  or _56375_ (_04580_, _04579_, _04578_);
  or _56376_ (_04581_, _04580_, _04577_);
  and _56377_ (_04582_, _04503_, _04458_);
  and _56378_ (_04583_, _04447_, _04502_);
  and _56379_ (_04584_, _04482_, _04475_);
  or _56380_ (_04585_, _04584_, _04583_);
  or _56381_ (_04586_, _04585_, _04582_);
  and _56382_ (_04587_, _04487_, _04481_);
  and _56383_ (_04588_, _04490_, _04470_);
  and _56384_ (_04589_, _04434_, _04443_);
  and _56385_ (_04590_, _04493_, _04486_);
  or _56386_ (_04591_, _04590_, _04589_);
  or _56387_ (_04592_, _04591_, _04588_);
  or _56388_ (_04593_, _04592_, _04587_);
  and _56389_ (_04594_, _04445_, _04479_);
  and _56390_ (_04595_, _04477_, _04489_);
  or _56391_ (_04596_, _04595_, _04594_);
  or _56392_ (_04597_, _04596_, _04593_);
  or _56393_ (_04598_, _04597_, _04586_);
  or _56394_ (_04599_, _04598_, _04581_);
  or _56395_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04599_, _04574_);
  not _56396_ (_04600_, _00231_);
  and _56397_ (_04601_, _04441_, _04600_);
  not _56398_ (_04602_, _00186_);
  and _56399_ (_04603_, _04454_, _04602_);
  not _56400_ (_04604_, _00077_);
  and _56401_ (_04605_, _04451_, _04604_);
  or _56402_ (_04606_, _04605_, _04603_);
  or _56403_ (_04607_, _04606_, _04601_);
  not _56404_ (_04608_, _00565_);
  and _56405_ (_04609_, _04464_, _04608_);
  not _56406_ (_04610_, _00518_);
  and _56407_ (_04611_, _04468_, _04610_);
  or _56408_ (_04612_, _04611_, _04609_);
  not _56409_ (_04613_, _00619_);
  and _56410_ (_04614_, _04461_, _04613_);
  not _56411_ (_04615_, _00272_);
  and _56412_ (_04616_, _04471_, _04615_);
  or _56413_ (_04617_, _04616_, _04614_);
  or _56414_ (_04618_, _04617_, _04612_);
  not _56415_ (_04619_, _00354_);
  and _56416_ (_04620_, _04477_, _04619_);
  not _56417_ (_04621_, _00701_);
  and _56418_ (_04622_, _04447_, _04621_);
  not _56419_ (_04623_, _00660_);
  and _56420_ (_04624_, _04503_, _04623_);
  or _56421_ (_04625_, _04624_, _04622_);
  or _56422_ (_04626_, _04625_, _04620_);
  not _56423_ (_04627_, _00395_);
  and _56424_ (_04628_, _04482_, _04627_);
  not _56425_ (_04629_, _00313_);
  and _56426_ (_04630_, _04490_, _04629_);
  not _56427_ (_04631_, _00477_);
  and _56428_ (_04632_, _04493_, _04631_);
  not _56429_ (_04633_, _00118_);
  and _56430_ (_04635_, _04434_, _04633_);
  or _56431_ (_04636_, _04635_, _04632_);
  or _56432_ (_04637_, _04636_, _04630_);
  or _56433_ (_04638_, _04637_, _04628_);
  not _56434_ (_04639_, _00436_);
  and _56435_ (_04640_, _04487_, _04639_);
  not _56436_ (_04641_, _00036_);
  and _56437_ (_04642_, _04445_, _04641_);
  or _56438_ (_04643_, _04642_, _04640_);
  or _56439_ (_04644_, _04643_, _04638_);
  or _56440_ (_04645_, _04644_, _04626_);
  or _56441_ (_04646_, _04645_, _04618_);
  or _56442_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04646_, _04607_);
  not _56443_ (_04647_, _00236_);
  and _56444_ (_04648_, _04441_, _04647_);
  not _56445_ (_04649_, _00195_);
  and _56446_ (_04650_, _04454_, _04649_);
  not _56447_ (_04651_, _00082_);
  and _56448_ (_04652_, _04451_, _04651_);
  or _56449_ (_04653_, _04652_, _04650_);
  or _56450_ (_04654_, _04653_, _04648_);
  not _56451_ (_04655_, _00624_);
  and _56452_ (_04656_, _04461_, _04655_);
  not _56453_ (_04657_, _00573_);
  and _56454_ (_04658_, _04464_, _04657_);
  or _56455_ (_04659_, _04658_, _04656_);
  not _56456_ (_04660_, _00523_);
  and _56457_ (_04661_, _04468_, _04660_);
  not _56458_ (_04662_, _00277_);
  and _56459_ (_04663_, _04471_, _04662_);
  or _56460_ (_04664_, _04663_, _04661_);
  or _56461_ (_04665_, _04664_, _04659_);
  not _56462_ (_04666_, _00400_);
  and _56463_ (_04667_, _04482_, _04666_);
  not _56464_ (_04668_, _00359_);
  and _56465_ (_04669_, _04477_, _04668_);
  or _56466_ (_04670_, _04669_, _04667_);
  not _56467_ (_04671_, _00441_);
  and _56468_ (_04672_, _04487_, _04671_);
  or _56469_ (_04673_, _04672_, _04670_);
  not _56470_ (_04674_, _00706_);
  and _56471_ (_04675_, _04447_, _04674_);
  not _56472_ (_04676_, _00318_);
  and _56473_ (_04677_, _04490_, _04676_);
  not _56474_ (_04678_, _00482_);
  and _56475_ (_04679_, _04493_, _04678_);
  not _56476_ (_04680_, _00123_);
  and _56477_ (_04681_, _04434_, _04680_);
  or _56478_ (_04682_, _04681_, _04679_);
  or _56479_ (_04683_, _04682_, _04677_);
  or _56480_ (_04684_, _04683_, _04675_);
  not _56481_ (_04685_, _00665_);
  and _56482_ (_04686_, _04503_, _04685_);
  not _56483_ (_04687_, _00041_);
  and _56484_ (_04688_, _04445_, _04687_);
  or _56485_ (_04689_, _04688_, _04686_);
  or _56486_ (_04690_, _04689_, _04684_);
  or _56487_ (_04691_, _04690_, _04673_);
  or _56488_ (_04692_, _04691_, _04665_);
  or _56489_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04692_, _04654_);
  not _56490_ (_04693_, _00241_);
  and _56491_ (_04694_, _04441_, _04693_);
  not _56492_ (_04695_, _00200_);
  and _56493_ (_04696_, _04454_, _04695_);
  not _56494_ (_04697_, _00087_);
  and _56495_ (_04698_, _04451_, _04697_);
  or _56496_ (_04699_, _04698_, _04696_);
  or _56497_ (_04700_, _04699_, _04694_);
  not _56498_ (_04701_, _00581_);
  and _56499_ (_04702_, _04464_, _04701_);
  not _56500_ (_04703_, _00528_);
  and _56501_ (_04704_, _04468_, _04703_);
  or _56502_ (_04705_, _04704_, _04702_);
  not _56503_ (_04706_, _00629_);
  and _56504_ (_04707_, _04461_, _04706_);
  not _56505_ (_04708_, _00282_);
  and _56506_ (_04709_, _04471_, _04708_);
  or _56507_ (_04710_, _04709_, _04707_);
  or _56508_ (_04711_, _04710_, _04705_);
  not _56509_ (_04712_, _00364_);
  and _56510_ (_04713_, _04477_, _04712_);
  not _56511_ (_04714_, _00711_);
  and _56512_ (_04715_, _04447_, _04714_);
  not _56513_ (_04716_, _00670_);
  and _56514_ (_04717_, _04503_, _04716_);
  or _56515_ (_04718_, _04717_, _04715_);
  or _56516_ (_04719_, _04718_, _04713_);
  not _56517_ (_04720_, _00405_);
  and _56518_ (_04721_, _04482_, _04720_);
  not _56519_ (_04722_, _00323_);
  and _56520_ (_04723_, _04490_, _04722_);
  not _56521_ (_04724_, _00487_);
  and _56522_ (_04725_, _04493_, _04724_);
  not _56523_ (_04726_, _00128_);
  and _56524_ (_04727_, _04434_, _04726_);
  or _56525_ (_04728_, _04727_, _04725_);
  or _56526_ (_04729_, _04728_, _04723_);
  or _56527_ (_04730_, _04729_, _04721_);
  not _56528_ (_04731_, _00446_);
  and _56529_ (_04732_, _04487_, _04731_);
  not _56530_ (_04733_, _00046_);
  and _56531_ (_04734_, _04445_, _04733_);
  or _56532_ (_04735_, _04734_, _04732_);
  or _56533_ (_04736_, _04735_, _04730_);
  or _56534_ (_04737_, _04736_, _04719_);
  or _56535_ (_04738_, _04737_, _04711_);
  or _56536_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04738_, _04700_);
  not _56537_ (_04739_, _00246_);
  and _56538_ (_04740_, _04441_, _04739_);
  not _56539_ (_04741_, _00205_);
  and _56540_ (_04742_, _04454_, _04741_);
  not _56541_ (_04743_, _00092_);
  and _56542_ (_04744_, _04451_, _04743_);
  or _56543_ (_04745_, _04744_, _04742_);
  or _56544_ (_04746_, _04745_, _04740_);
  not _56545_ (_04747_, _00589_);
  and _56546_ (_04748_, _04464_, _04747_);
  not _56547_ (_04749_, _00533_);
  and _56548_ (_04750_, _04468_, _04749_);
  or _56549_ (_04751_, _04750_, _04748_);
  not _56550_ (_04752_, _00634_);
  and _56551_ (_04753_, _04461_, _04752_);
  not _56552_ (_04754_, _00287_);
  and _56553_ (_04755_, _04471_, _04754_);
  or _56554_ (_04756_, _04755_, _04753_);
  or _56555_ (_04757_, _04756_, _04751_);
  not _56556_ (_04758_, _00369_);
  and _56557_ (_04759_, _04477_, _04758_);
  not _56558_ (_04760_, _00716_);
  and _56559_ (_04761_, _04447_, _04760_);
  not _56560_ (_04762_, _00675_);
  and _56561_ (_04763_, _04503_, _04762_);
  or _56562_ (_04764_, _04763_, _04761_);
  or _56563_ (_04765_, _04764_, _04759_);
  not _56564_ (_04766_, _00451_);
  and _56565_ (_04767_, _04487_, _04766_);
  not _56566_ (_04768_, _00410_);
  and _56567_ (_04769_, _04482_, _04768_);
  or _56568_ (_04770_, _04769_, _04767_);
  not _56569_ (_04771_, _00051_);
  and _56570_ (_04772_, _04445_, _04771_);
  not _56571_ (_04773_, _00328_);
  and _56572_ (_04774_, _04490_, _04773_);
  not _56573_ (_04775_, _00492_);
  and _56574_ (_04776_, _04493_, _04775_);
  not _56575_ (_04777_, _00133_);
  and _56576_ (_04778_, _04434_, _04777_);
  or _56577_ (_04779_, _04778_, _04776_);
  or _56578_ (_04780_, _04779_, _04774_);
  or _56579_ (_04781_, _04780_, _04772_);
  or _56580_ (_04782_, _04781_, _04770_);
  or _56581_ (_04783_, _04782_, _04765_);
  or _56582_ (_04784_, _04783_, _04757_);
  or _56583_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04784_, _04746_);
  not _56584_ (_04785_, _00210_);
  and _56585_ (_04786_, _04454_, _04785_);
  not _56586_ (_04787_, _00251_);
  and _56587_ (_04788_, _04441_, _04787_);
  not _56588_ (_04789_, _00097_);
  and _56589_ (_04790_, _04451_, _04789_);
  or _56590_ (_04791_, _04790_, _04788_);
  or _56591_ (_04792_, _04791_, _04786_);
  not _56592_ (_04793_, _00639_);
  and _56593_ (_04794_, _04461_, _04793_);
  not _56594_ (_04795_, _00597_);
  and _56595_ (_04796_, _04464_, _04795_);
  or _56596_ (_04797_, _04796_, _04794_);
  not _56597_ (_04798_, _00538_);
  and _56598_ (_04799_, _04468_, _04798_);
  not _56599_ (_04800_, _00292_);
  and _56600_ (_04801_, _04471_, _04800_);
  or _56601_ (_04802_, _04801_, _04799_);
  or _56602_ (_04803_, _04802_, _04797_);
  not _56603_ (_04804_, _00374_);
  and _56604_ (_04805_, _04477_, _04804_);
  not _56605_ (_04806_, _00415_);
  and _56606_ (_04807_, _04482_, _04806_);
  or _56607_ (_04808_, _04807_, _04805_);
  not _56608_ (_04809_, _00056_);
  and _56609_ (_04810_, _04445_, _04809_);
  or _56610_ (_04811_, _04810_, _04808_);
  not _56611_ (_04812_, _00721_);
  and _56612_ (_04813_, _04447_, _04812_);
  not _56613_ (_04814_, _00333_);
  and _56614_ (_04815_, _04490_, _04814_);
  not _56615_ (_04816_, _00497_);
  and _56616_ (_04817_, _04493_, _04816_);
  not _56617_ (_04818_, _00140_);
  and _56618_ (_04819_, _04434_, _04818_);
  or _56619_ (_04820_, _04819_, _04817_);
  or _56620_ (_04821_, _04820_, _04815_);
  or _56621_ (_04822_, _04821_, _04813_);
  not _56622_ (_04823_, _00680_);
  and _56623_ (_04824_, _04503_, _04823_);
  not _56624_ (_04825_, _00456_);
  and _56625_ (_04826_, _04487_, _04825_);
  or _56626_ (_04827_, _04826_, _04824_);
  or _56627_ (_04828_, _04827_, _04822_);
  or _56628_ (_04829_, _04828_, _04811_);
  or _56629_ (_04830_, _04829_, _04803_);
  or _56630_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04830_, _04792_);
  not _56631_ (_04831_, _00215_);
  and _56632_ (_04832_, _04454_, _04831_);
  not _56633_ (_04833_, _00256_);
  and _56634_ (_04834_, _04441_, _04833_);
  not _56635_ (_04835_, _00102_);
  and _56636_ (_04836_, _04451_, _04835_);
  or _56637_ (_04837_, _04836_, _04834_);
  or _56638_ (_04838_, _04837_, _04832_);
  not _56639_ (_04839_, _00644_);
  and _56640_ (_04840_, _04461_, _04839_);
  not _56641_ (_04841_, _00603_);
  and _56642_ (_04842_, _04464_, _04841_);
  or _56643_ (_04843_, _04842_, _04840_);
  not _56644_ (_04844_, _00543_);
  and _56645_ (_04845_, _04468_, _04844_);
  not _56646_ (_04846_, _00297_);
  and _56647_ (_04847_, _04471_, _04846_);
  or _56648_ (_04848_, _04847_, _04845_);
  or _56649_ (_04849_, _04848_, _04843_);
  not _56650_ (_04850_, _00379_);
  and _56651_ (_04851_, _04477_, _04850_);
  not _56652_ (_04852_, _00420_);
  and _56653_ (_04853_, _04482_, _04852_);
  or _56654_ (_04854_, _04853_, _04851_);
  not _56655_ (_04855_, _00061_);
  and _56656_ (_04856_, _04445_, _04855_);
  or _56657_ (_04857_, _04856_, _04854_);
  not _56658_ (_04858_, _00726_);
  and _56659_ (_04859_, _04447_, _04858_);
  not _56660_ (_04860_, _00338_);
  and _56661_ (_04861_, _04490_, _04860_);
  not _56662_ (_04862_, _00502_);
  and _56663_ (_04863_, _04493_, _04862_);
  not _56664_ (_04864_, _00151_);
  and _56665_ (_04865_, _04434_, _04864_);
  or _56666_ (_04866_, _04865_, _04863_);
  or _56667_ (_04867_, _04866_, _04861_);
  or _56668_ (_04868_, _04867_, _04859_);
  not _56669_ (_04869_, _00685_);
  and _56670_ (_04870_, _04503_, _04869_);
  not _56671_ (_04871_, _00461_);
  and _56672_ (_04872_, _04487_, _04871_);
  or _56673_ (_04873_, _04872_, _04870_);
  or _56674_ (_04874_, _04873_, _04868_);
  or _56675_ (_04875_, _04874_, _04857_);
  or _56676_ (_04876_, _04875_, _04849_);
  or _56677_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04876_, _04838_);
  not _56678_ (_04877_, _00261_);
  and _56679_ (_04878_, _04441_, _04877_);
  not _56680_ (_04879_, _00220_);
  and _56681_ (_04880_, _04454_, _04879_);
  not _56682_ (_04881_, _00107_);
  and _56683_ (_04882_, _04451_, _04881_);
  or _56684_ (_04883_, _04882_, _04880_);
  or _56685_ (_04884_, _04883_, _04878_);
  not _56686_ (_04885_, _00608_);
  and _56687_ (_04886_, _04464_, _04885_);
  not _56688_ (_04887_, _00548_);
  and _56689_ (_04888_, _04468_, _04887_);
  or _56690_ (_04889_, _04888_, _04886_);
  not _56691_ (_04890_, _00649_);
  and _56692_ (_04891_, _04461_, _04890_);
  not _56693_ (_04892_, _00302_);
  and _56694_ (_04893_, _04471_, _04892_);
  or _56695_ (_04894_, _04893_, _04891_);
  or _56696_ (_04895_, _04894_, _04889_);
  not _56697_ (_04896_, _00384_);
  and _56698_ (_04897_, _04477_, _04896_);
  not _56699_ (_04898_, _00731_);
  and _56700_ (_04899_, _04447_, _04898_);
  not _56701_ (_04900_, _00690_);
  and _56702_ (_04901_, _04503_, _04900_);
  or _56703_ (_04902_, _04901_, _04899_);
  or _56704_ (_04903_, _04902_, _04897_);
  not _56705_ (_04904_, _00466_);
  and _56706_ (_04905_, _04487_, _04904_);
  not _56707_ (_04906_, _00425_);
  and _56708_ (_04907_, _04482_, _04906_);
  or _56709_ (_04908_, _04907_, _04905_);
  not _56710_ (_04909_, _00066_);
  and _56711_ (_04910_, _04445_, _04909_);
  not _56712_ (_04911_, _00343_);
  and _56713_ (_04912_, _04490_, _04911_);
  not _56714_ (_04913_, _00507_);
  and _56715_ (_04914_, _04493_, _04913_);
  not _56716_ (_04915_, _00162_);
  and _56717_ (_04916_, _04434_, _04915_);
  or _56718_ (_04917_, _04916_, _04914_);
  or _56719_ (_04918_, _04917_, _04912_);
  or _56720_ (_04919_, _04918_, _04910_);
  or _56721_ (_04920_, _04919_, _04908_);
  or _56722_ (_04921_, _04920_, _04903_);
  or _56723_ (_04922_, _04921_, _04895_);
  or _56724_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04922_, _04884_);
  and _56725_ (_04923_, _04454_, _04633_);
  and _56726_ (_04924_, _04441_, _04602_);
  and _56727_ (_04925_, _04451_, _04641_);
  or _56728_ (_04926_, _04925_, _04924_);
  or _56729_ (_04927_, _04926_, _04923_);
  and _56730_ (_04928_, _04461_, _04608_);
  and _56731_ (_04929_, _04464_, _04610_);
  or _56732_ (_04930_, _04929_, _04928_);
  and _56733_ (_04931_, _04468_, _04631_);
  and _56734_ (_04932_, _04471_, _04600_);
  or _56735_ (_04933_, _04932_, _04931_);
  or _56736_ (_04934_, _04933_, _04930_);
  and _56737_ (_04935_, _04503_, _04613_);
  and _56738_ (_04936_, _04445_, _04621_);
  and _56739_ (_04937_, _04447_, _04623_);
  or _56740_ (_04938_, _04937_, _04936_);
  or _56741_ (_04939_, _04938_, _04935_);
  and _56742_ (_04940_, _04482_, _04619_);
  and _56743_ (_04941_, _04490_, _04615_);
  and _56744_ (_04942_, _04493_, _04639_);
  and _56745_ (_04943_, _04434_, _04604_);
  or _56746_ (_04944_, _04943_, _04942_);
  or _56747_ (_04945_, _04944_, _04941_);
  or _56748_ (_04946_, _04945_, _04940_);
  and _56749_ (_04947_, _04487_, _04627_);
  and _56750_ (_04948_, _04477_, _04629_);
  or _56751_ (_04949_, _04948_, _04947_);
  or _56752_ (_04950_, _04949_, _04946_);
  or _56753_ (_04951_, _04950_, _04939_);
  or _56754_ (_04952_, _04951_, _04934_);
  or _56755_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04952_, _04927_);
  and _56756_ (_04953_, _04454_, _04680_);
  and _56757_ (_04954_, _04441_, _04649_);
  and _56758_ (_04955_, _04451_, _04687_);
  or _56759_ (_04956_, _04955_, _04954_);
  or _56760_ (_04957_, _04956_, _04953_);
  and _56761_ (_04958_, _04464_, _04660_);
  and _56762_ (_04959_, _04461_, _04657_);
  or _56763_ (_04960_, _04959_, _04958_);
  and _56764_ (_04961_, _04468_, _04678_);
  and _56765_ (_04962_, _04471_, _04647_);
  or _56766_ (_04963_, _04962_, _04961_);
  or _56767_ (_04964_, _04963_, _04960_);
  and _56768_ (_04965_, _04503_, _04655_);
  and _56769_ (_04966_, _04447_, _04685_);
  and _56770_ (_04967_, _04477_, _04676_);
  or _56771_ (_04968_, _04967_, _04966_);
  or _56772_ (_04969_, _04968_, _04965_);
  and _56773_ (_04970_, _04487_, _04666_);
  and _56774_ (_04971_, _04490_, _04662_);
  and _56775_ (_04972_, _04493_, _04671_);
  and _56776_ (_04973_, _04434_, _04651_);
  or _56777_ (_04974_, _04973_, _04972_);
  or _56778_ (_04975_, _04974_, _04971_);
  or _56779_ (_04976_, _04975_, _04970_);
  and _56780_ (_04977_, _04445_, _04674_);
  and _56781_ (_04978_, _04482_, _04668_);
  or _56782_ (_04979_, _04978_, _04977_);
  or _56783_ (_04980_, _04979_, _04976_);
  or _56784_ (_04981_, _04980_, _04969_);
  or _56785_ (_04982_, _04981_, _04964_);
  or _56786_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04982_, _04957_);
  and _56787_ (_04983_, _04454_, _04726_);
  and _56788_ (_04984_, _04441_, _04695_);
  and _56789_ (_04985_, _04451_, _04733_);
  or _56790_ (_04986_, _04985_, _04984_);
  or _56791_ (_04987_, _04986_, _04983_);
  and _56792_ (_04988_, _04461_, _04701_);
  and _56793_ (_04989_, _04464_, _04703_);
  or _56794_ (_04990_, _04989_, _04988_);
  and _56795_ (_04991_, _04468_, _04724_);
  and _56796_ (_04992_, _04471_, _04693_);
  or _56797_ (_04993_, _04992_, _04991_);
  or _56798_ (_04994_, _04993_, _04990_);
  and _56799_ (_04995_, _04503_, _04706_);
  and _56800_ (_04996_, _04445_, _04714_);
  and _56801_ (_04997_, _04447_, _04716_);
  or _56802_ (_04998_, _04997_, _04996_);
  or _56803_ (_04999_, _04998_, _04995_);
  and _56804_ (_05000_, _04482_, _04712_);
  and _56805_ (_05001_, _04490_, _04708_);
  and _56806_ (_05002_, _04493_, _04731_);
  and _56807_ (_05003_, _04434_, _04697_);
  or _56808_ (_05004_, _05003_, _05002_);
  or _56809_ (_05005_, _05004_, _05001_);
  or _56810_ (_05006_, _05005_, _05000_);
  and _56811_ (_05007_, _04487_, _04720_);
  and _56812_ (_05008_, _04477_, _04722_);
  or _56813_ (_05009_, _05008_, _05007_);
  or _56814_ (_05010_, _05009_, _05006_);
  or _56815_ (_05011_, _05010_, _04999_);
  or _56816_ (_05012_, _05011_, _04994_);
  or _56817_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _05012_, _04987_);
  and _56818_ (_05013_, _04441_, _04741_);
  and _56819_ (_05014_, _04451_, _04771_);
  and _56820_ (_05015_, _04454_, _04777_);
  or _56821_ (_05016_, _05015_, _05014_);
  or _56822_ (_05017_, _05016_, _05013_);
  and _56823_ (_05018_, _04461_, _04747_);
  and _56824_ (_05019_, _04471_, _04739_);
  or _56825_ (_05020_, _05019_, _05018_);
  and _56826_ (_05021_, _04464_, _04749_);
  and _56827_ (_05022_, _04468_, _04775_);
  or _56828_ (_05023_, _05022_, _05021_);
  or _56829_ (_05024_, _05023_, _05020_);
  and _56830_ (_05025_, _04477_, _04773_);
  and _56831_ (_05026_, _04503_, _04752_);
  and _56832_ (_05027_, _04482_, _04758_);
  or _56833_ (_05028_, _05027_, _05026_);
  or _56834_ (_05029_, _05028_, _05025_);
  and _56835_ (_05030_, _04487_, _04768_);
  and _56836_ (_05031_, _04490_, _04754_);
  and _56837_ (_05032_, _04493_, _04766_);
  and _56838_ (_05033_, _04434_, _04743_);
  or _56839_ (_05034_, _05033_, _05032_);
  or _56840_ (_05035_, _05034_, _05031_);
  or _56841_ (_05036_, _05035_, _05030_);
  and _56842_ (_05037_, _04445_, _04760_);
  and _56843_ (_05038_, _04447_, _04762_);
  or _56844_ (_05039_, _05038_, _05037_);
  or _56845_ (_05040_, _05039_, _05036_);
  or _56846_ (_05041_, _05040_, _05029_);
  or _56847_ (_05042_, _05041_, _05024_);
  or _56848_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _05042_, _05017_);
  and _56849_ (_05043_, _04451_, _04809_);
  and _56850_ (_05044_, _04441_, _04785_);
  and _56851_ (_05045_, _04454_, _04818_);
  or _56852_ (_05046_, _05045_, _05044_);
  or _56853_ (_05047_, _05046_, _05043_);
  and _56854_ (_05048_, _04461_, _04795_);
  and _56855_ (_05049_, _04464_, _04798_);
  or _56856_ (_05050_, _05049_, _05048_);
  and _56857_ (_05051_, _04468_, _04816_);
  and _56858_ (_05052_, _04471_, _04787_);
  or _56859_ (_05053_, _05052_, _05051_);
  or _56860_ (_05054_, _05053_, _05050_);
  and _56861_ (_05055_, _04487_, _04806_);
  and _56862_ (_05056_, _04447_, _04823_);
  and _56863_ (_05057_, _04477_, _04814_);
  or _56864_ (_05058_, _05057_, _05056_);
  or _56865_ (_05059_, _05058_, _05055_);
  and _56866_ (_05060_, _04482_, _04804_);
  and _56867_ (_05061_, _04490_, _04800_);
  and _56868_ (_05062_, _04493_, _04825_);
  and _56869_ (_05063_, _04434_, _04789_);
  or _56870_ (_05064_, _05063_, _05062_);
  or _56871_ (_05065_, _05064_, _05061_);
  or _56872_ (_05066_, _05065_, _05060_);
  and _56873_ (_05067_, _04445_, _04812_);
  and _56874_ (_05068_, _04503_, _04793_);
  or _56875_ (_05069_, _05068_, _05067_);
  or _56876_ (_05070_, _05069_, _05066_);
  or _56877_ (_05071_, _05070_, _05059_);
  or _56878_ (_05072_, _05071_, _05054_);
  or _56879_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _05072_, _05047_);
  and _56880_ (_05073_, _04451_, _04855_);
  and _56881_ (_05074_, _04441_, _04831_);
  and _56882_ (_05075_, _04454_, _04864_);
  or _56883_ (_05077_, _05075_, _05074_);
  or _56884_ (_05079_, _05077_, _05073_);
  and _56885_ (_05081_, _04461_, _04841_);
  and _56886_ (_05083_, _04468_, _04862_);
  or _56887_ (_05085_, _05083_, _05081_);
  and _56888_ (_05087_, _04464_, _04844_);
  and _56889_ (_05089_, _04471_, _04833_);
  or _56890_ (_05090_, _05089_, _05087_);
  or _56891_ (_05091_, _05090_, _05085_);
  and _56892_ (_05092_, _04487_, _04852_);
  and _56893_ (_05093_, _04447_, _04869_);
  and _56894_ (_05094_, _04477_, _04860_);
  or _56895_ (_05095_, _05094_, _05093_);
  or _56896_ (_05097_, _05095_, _05092_);
  and _56897_ (_05098_, _04482_, _04850_);
  and _56898_ (_05100_, _04490_, _04846_);
  and _56899_ (_05101_, _04493_, _04871_);
  and _56900_ (_05102_, _04434_, _04835_);
  or _56901_ (_05104_, _05102_, _05101_);
  or _56902_ (_05105_, _05104_, _05100_);
  or _56903_ (_05106_, _05105_, _05098_);
  and _56904_ (_05108_, _04445_, _04858_);
  and _56905_ (_05109_, _04503_, _04839_);
  or _56906_ (_05110_, _05109_, _05108_);
  or _56907_ (_05112_, _05110_, _05106_);
  or _56908_ (_05113_, _05112_, _05097_);
  or _56909_ (_05114_, _05113_, _05091_);
  or _56910_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _05114_, _05079_);
  and _56911_ (_05116_, _04454_, _04915_);
  and _56912_ (_05117_, _04441_, _04879_);
  and _56913_ (_05119_, _04451_, _04909_);
  or _56914_ (_05120_, _05119_, _05117_);
  or _56915_ (_05121_, _05120_, _05116_);
  and _56916_ (_05123_, _04461_, _04885_);
  and _56917_ (_05124_, _04464_, _04887_);
  or _56918_ (_05125_, _05124_, _05123_);
  and _56919_ (_05127_, _04468_, _04913_);
  and _56920_ (_05128_, _04471_, _04877_);
  or _56921_ (_05129_, _05128_, _05127_);
  or _56922_ (_05130_, _05129_, _05125_);
  and _56923_ (_05131_, _04503_, _04890_);
  and _56924_ (_05132_, _04445_, _04898_);
  and _56925_ (_05133_, _04447_, _04900_);
  or _56926_ (_05134_, _05133_, _05132_);
  or _56927_ (_05135_, _05134_, _05131_);
  and _56928_ (_05136_, _04482_, _04896_);
  and _56929_ (_05137_, _04490_, _04892_);
  and _56930_ (_05138_, _04493_, _04904_);
  and _56931_ (_05139_, _04434_, _04881_);
  or _56932_ (_05140_, _05139_, _05138_);
  or _56933_ (_05141_, _05140_, _05137_);
  or _56934_ (_05142_, _05141_, _05136_);
  and _56935_ (_05143_, _04487_, _04906_);
  and _56936_ (_05144_, _04477_, _04911_);
  or _56937_ (_05145_, _05144_, _05143_);
  or _56938_ (_05146_, _05145_, _05142_);
  or _56939_ (_05147_, _05146_, _05135_);
  or _56940_ (_05149_, _05147_, _05130_);
  or _56941_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _05149_, _05121_);
  and _56942_ (_05151_, _04441_, _04604_);
  and _56943_ (_05152_, _04451_, _04623_);
  and _56944_ (_05153_, _04454_, _04641_);
  or _56945_ (_05155_, _05153_, _05152_);
  or _56946_ (_05156_, _05155_, _05151_);
  and _56947_ (_05157_, _04464_, _04639_);
  and _56948_ (_05159_, _04461_, _04631_);
  or _56949_ (_05160_, _05159_, _05157_);
  and _56950_ (_05161_, _04468_, _04627_);
  and _56951_ (_05163_, _04471_, _04633_);
  or _56952_ (_05164_, _05163_, _05161_);
  or _56953_ (_05165_, _05164_, _05160_);
  and _56954_ (_05167_, _04503_, _04610_);
  and _56955_ (_05168_, _04447_, _04608_);
  and _56956_ (_05169_, _04482_, _04615_);
  or _56957_ (_05171_, _05169_, _05168_);
  or _56958_ (_05172_, _05171_, _05167_);
  and _56959_ (_05173_, _04487_, _04629_);
  and _56960_ (_05175_, _04490_, _04602_);
  and _56961_ (_05176_, _04434_, _04621_);
  and _56962_ (_05177_, _04493_, _04619_);
  or _56963_ (_05179_, _05177_, _05176_);
  or _56964_ (_05180_, _05179_, _05175_);
  or _56965_ (_05181_, _05180_, _05173_);
  and _56966_ (_05182_, _04445_, _04613_);
  and _56967_ (_05183_, _04477_, _04600_);
  or _56968_ (_05184_, _05183_, _05182_);
  or _56969_ (_05185_, _05184_, _05181_);
  or _56970_ (_05186_, _05185_, _05172_);
  or _56971_ (_05187_, _05186_, _05165_);
  or _56972_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _05187_, _05156_);
  and _56973_ (_05188_, _04441_, _04651_);
  and _56974_ (_05189_, _04451_, _04685_);
  and _56975_ (_05190_, _04454_, _04687_);
  or _56976_ (_05191_, _05190_, _05189_);
  or _56977_ (_05192_, _05191_, _05188_);
  and _56978_ (_05193_, _04464_, _04671_);
  and _56979_ (_05194_, _04471_, _04680_);
  or _56980_ (_05195_, _05194_, _05193_);
  and _56981_ (_05196_, _04461_, _04678_);
  and _56982_ (_05197_, _04468_, _04666_);
  or _56983_ (_05198_, _05197_, _05196_);
  or _56984_ (_05200_, _05198_, _05195_);
  and _56985_ (_05201_, _04503_, _04660_);
  and _56986_ (_05203_, _04447_, _04657_);
  and _56987_ (_05204_, _04482_, _04662_);
  or _56988_ (_05205_, _05204_, _05203_);
  or _56989_ (_05207_, _05205_, _05201_);
  and _56990_ (_05208_, _04487_, _04676_);
  and _56991_ (_05209_, _04490_, _04649_);
  and _56992_ (_05211_, _04434_, _04674_);
  and _56993_ (_05212_, _04493_, _04668_);
  or _56994_ (_05213_, _05212_, _05211_);
  or _56995_ (_05215_, _05213_, _05209_);
  or _56996_ (_05216_, _05215_, _05208_);
  and _56997_ (_05217_, _04445_, _04655_);
  and _56998_ (_05219_, _04477_, _04647_);
  or _56999_ (_05220_, _05219_, _05217_);
  or _57000_ (_05221_, _05220_, _05216_);
  or _57001_ (_05223_, _05221_, _05207_);
  or _57002_ (_05224_, _05223_, _05200_);
  or _57003_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _05224_, _05192_);
  and _57004_ (_05226_, _04441_, _04697_);
  and _57005_ (_05227_, _04451_, _04716_);
  and _57006_ (_05228_, _04454_, _04733_);
  or _57007_ (_05230_, _05228_, _05227_);
  or _57008_ (_05231_, _05230_, _05226_);
  and _57009_ (_05232_, _04464_, _04731_);
  and _57010_ (_05233_, _04471_, _04726_);
  or _57011_ (_05234_, _05233_, _05232_);
  and _57012_ (_05235_, _04461_, _04724_);
  and _57013_ (_05236_, _04468_, _04720_);
  or _57014_ (_05237_, _05236_, _05235_);
  or _57015_ (_05238_, _05237_, _05234_);
  and _57016_ (_05239_, _04503_, _04703_);
  and _57017_ (_05240_, _04447_, _04701_);
  and _57018_ (_05241_, _04482_, _04708_);
  or _57019_ (_05242_, _05241_, _05240_);
  or _57020_ (_05243_, _05242_, _05239_);
  and _57021_ (_05244_, _04487_, _04722_);
  and _57022_ (_05245_, _04490_, _04695_);
  and _57023_ (_05246_, _04434_, _04714_);
  and _57024_ (_05247_, _04493_, _04712_);
  or _57025_ (_05248_, _05247_, _05246_);
  or _57026_ (_05249_, _05248_, _05245_);
  or _57027_ (_05250_, _05249_, _05244_);
  and _57028_ (_05252_, _04445_, _04706_);
  and _57029_ (_05253_, _04477_, _04693_);
  or _57030_ (_05255_, _05253_, _05252_);
  or _57031_ (_05256_, _05255_, _05250_);
  or _57032_ (_05257_, _05256_, _05243_);
  or _57033_ (_05259_, _05257_, _05238_);
  or _57034_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _05259_, _05231_);
  and _57035_ (_05260_, _04441_, _04743_);
  and _57036_ (_05262_, _04451_, _04762_);
  and _57037_ (_05263_, _04454_, _04771_);
  or _57038_ (_05264_, _05263_, _05262_);
  or _57039_ (_05266_, _05264_, _05260_);
  and _57040_ (_05267_, _04464_, _04766_);
  and _57041_ (_05268_, _04461_, _04775_);
  or _57042_ (_05270_, _05268_, _05267_);
  and _57043_ (_05271_, _04468_, _04768_);
  and _57044_ (_05272_, _04471_, _04777_);
  or _57045_ (_05274_, _05272_, _05271_);
  or _57046_ (_05275_, _05274_, _05270_);
  and _57047_ (_05276_, _04503_, _04749_);
  and _57048_ (_05278_, _04447_, _04747_);
  and _57049_ (_05279_, _04482_, _04754_);
  or _57050_ (_05280_, _05279_, _05278_);
  or _57051_ (_05282_, _05280_, _05276_);
  and _57052_ (_05283_, _04487_, _04773_);
  and _57053_ (_05284_, _04490_, _04741_);
  and _57054_ (_05285_, _04434_, _04760_);
  and _57055_ (_05286_, _04493_, _04758_);
  or _57056_ (_05287_, _05286_, _05285_);
  or _57057_ (_05288_, _05287_, _05284_);
  or _57058_ (_05289_, _05288_, _05283_);
  and _57059_ (_05290_, _04445_, _04752_);
  and _57060_ (_05291_, _04477_, _04739_);
  or _57061_ (_05292_, _05291_, _05290_);
  or _57062_ (_05293_, _05292_, _05289_);
  or _57063_ (_05294_, _05293_, _05282_);
  or _57064_ (_05295_, _05294_, _05275_);
  or _57065_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _05295_, _05266_);
  and _57066_ (_05296_, _04454_, _04809_);
  and _57067_ (_05297_, _04471_, _04818_);
  or _57068_ (_05298_, _05297_, _05296_);
  and _57069_ (_05299_, _04441_, _04789_);
  and _57070_ (_05300_, _04487_, _04814_);
  and _57071_ (_05301_, _04482_, _04800_);
  or _57072_ (_05303_, _05301_, _05300_);
  and _57073_ (_05304_, _04490_, _04785_);
  and _57074_ (_05306_, _04477_, _04787_);
  or _57075_ (_05307_, _05306_, _05304_);
  or _57076_ (_05308_, _05307_, _05303_);
  or _57077_ (_05310_, _05308_, _05299_);
  or _57078_ (_05311_, _05310_, _05298_);
  and _57079_ (_05312_, _04451_, _04823_);
  and _57080_ (_05314_, _04468_, _04806_);
  and _57081_ (_05315_, _04461_, _04816_);
  and _57082_ (_05316_, _04503_, _04798_);
  or _57083_ (_05318_, _05316_, _05315_);
  or _57084_ (_05319_, _05318_, _05314_);
  and _57085_ (_05320_, _04464_, _04825_);
  and _57086_ (_05322_, _04447_, _04795_);
  and _57087_ (_05323_, _04434_, _04812_);
  and _57088_ (_05324_, _04493_, _04804_);
  or _57089_ (_05326_, _05324_, _05323_);
  and _57090_ (_05327_, _04445_, _04793_);
  or _57091_ (_05328_, _05327_, _05326_);
  or _57092_ (_05330_, _05328_, _05322_);
  or _57093_ (_05331_, _05330_, _05320_);
  or _57094_ (_05332_, _05331_, _05319_);
  or _57095_ (_05334_, _05332_, _05312_);
  or _57096_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _05334_, _05311_);
  and _57097_ (_05335_, _04454_, _04855_);
  and _57098_ (_05336_, _04471_, _04864_);
  or _57099_ (_05337_, _05336_, _05335_);
  and _57100_ (_05338_, _04441_, _04835_);
  and _57101_ (_05339_, _04487_, _04860_);
  and _57102_ (_05340_, _04482_, _04846_);
  or _57103_ (_05341_, _05340_, _05339_);
  and _57104_ (_05342_, _04490_, _04831_);
  and _57105_ (_05343_, _04477_, _04833_);
  or _57106_ (_05344_, _05343_, _05342_);
  or _57107_ (_05345_, _05344_, _05341_);
  or _57108_ (_05346_, _05345_, _05338_);
  or _57109_ (_05347_, _05346_, _05337_);
  and _57110_ (_05348_, _04451_, _04869_);
  and _57111_ (_05349_, _04468_, _04852_);
  and _57112_ (_05350_, _04461_, _04862_);
  and _57113_ (_05351_, _04503_, _04844_);
  or _57114_ (_05352_, _05351_, _05350_);
  or _57115_ (_05353_, _05352_, _05349_);
  and _57116_ (_05355_, _04464_, _04871_);
  and _57117_ (_05356_, _04447_, _04841_);
  and _57118_ (_05358_, _04434_, _04858_);
  and _57119_ (_05359_, _04493_, _04850_);
  or _57120_ (_05360_, _05359_, _05358_);
  and _57121_ (_05362_, _04445_, _04839_);
  or _57122_ (_05363_, _05362_, _05360_);
  or _57123_ (_05364_, _05363_, _05356_);
  or _57124_ (_05366_, _05364_, _05355_);
  or _57125_ (_05367_, _05366_, _05353_);
  or _57126_ (_05368_, _05367_, _05348_);
  or _57127_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05368_, _05347_);
  and _57128_ (_05370_, _04441_, _04881_);
  and _57129_ (_05371_, _04451_, _04900_);
  and _57130_ (_05373_, _04454_, _04909_);
  or _57131_ (_05374_, _05373_, _05371_);
  or _57132_ (_05375_, _05374_, _05370_);
  and _57133_ (_05377_, _04464_, _04904_);
  and _57134_ (_05378_, _04461_, _04913_);
  or _57135_ (_05379_, _05378_, _05377_);
  and _57136_ (_05381_, _04468_, _04906_);
  and _57137_ (_05382_, _04471_, _04915_);
  or _57138_ (_05383_, _05382_, _05381_);
  or _57139_ (_05385_, _05383_, _05379_);
  and _57140_ (_05386_, _04503_, _04887_);
  and _57141_ (_05387_, _04445_, _04890_);
  and _57142_ (_05388_, _04447_, _04885_);
  or _57143_ (_05389_, _05388_, _05387_);
  or _57144_ (_05390_, _05389_, _05386_);
  and _57145_ (_05391_, _04482_, _04892_);
  and _57146_ (_05392_, _04490_, _04879_);
  and _57147_ (_05393_, _04434_, _04898_);
  and _57148_ (_05394_, _04493_, _04896_);
  or _57149_ (_05395_, _05394_, _05393_);
  or _57150_ (_05396_, _05395_, _05392_);
  or _57151_ (_05397_, _05396_, _05391_);
  and _57152_ (_05398_, _04487_, _04911_);
  and _57153_ (_05399_, _04477_, _04877_);
  or _57154_ (_05400_, _05399_, _05398_);
  or _57155_ (_05401_, _05400_, _05397_);
  or _57156_ (_05402_, _05401_, _05390_);
  or _57157_ (_05403_, _05402_, _05385_);
  or _57158_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05403_, _05375_);
  and _57159_ (_05404_, _04451_, _04621_);
  and _57160_ (_05406_, _04441_, _04633_);
  and _57161_ (_05407_, _04454_, _04604_);
  or _57162_ (_05409_, _05407_, _05406_);
  or _57163_ (_05410_, _05409_, _05404_);
  and _57164_ (_05411_, _04461_, _04610_);
  and _57165_ (_05413_, _04468_, _04639_);
  or _57166_ (_05414_, _05413_, _05411_);
  and _57167_ (_05415_, _04464_, _04631_);
  and _57168_ (_05417_, _04471_, _04602_);
  or _57169_ (_05418_, _05417_, _05415_);
  or _57170_ (_05419_, _05418_, _05414_);
  and _57171_ (_05421_, _04487_, _04619_);
  and _57172_ (_05422_, _04447_, _04613_);
  and _57173_ (_05423_, _04477_, _04615_);
  or _57174_ (_05425_, _05423_, _05422_);
  or _57175_ (_05426_, _05425_, _05421_);
  and _57176_ (_05427_, _04482_, _04629_);
  and _57177_ (_05429_, _04490_, _04600_);
  and _57178_ (_05430_, _04493_, _04627_);
  and _57179_ (_05431_, _04434_, _04641_);
  or _57180_ (_05433_, _05431_, _05430_);
  or _57181_ (_05434_, _05433_, _05429_);
  or _57182_ (_05435_, _05434_, _05427_);
  and _57183_ (_05437_, _04445_, _04623_);
  and _57184_ (_05438_, _04503_, _04608_);
  or _57185_ (_05439_, _05438_, _05437_);
  or _57186_ (_05440_, _05439_, _05435_);
  or _57187_ (_05441_, _05440_, _05426_);
  or _57188_ (_05442_, _05441_, _05419_);
  or _57189_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05442_, _05410_);
  and _57190_ (_05443_, _04451_, _04674_);
  and _57191_ (_05444_, _04454_, _04651_);
  and _57192_ (_05445_, _04441_, _04680_);
  or _57193_ (_05446_, _05445_, _05444_);
  or _57194_ (_05447_, _05446_, _05443_);
  and _57195_ (_05448_, _04461_, _04660_);
  and _57196_ (_05449_, _04464_, _04678_);
  or _57197_ (_05450_, _05449_, _05448_);
  and _57198_ (_05451_, _04468_, _04671_);
  and _57199_ (_05452_, _04471_, _04649_);
  or _57200_ (_05453_, _05452_, _05451_);
  or _57201_ (_05454_, _05453_, _05450_);
  and _57202_ (_05455_, _04482_, _04676_);
  and _57203_ (_05456_, _04503_, _04657_);
  and _57204_ (_05458_, _04487_, _04668_);
  or _57205_ (_05459_, _05458_, _05456_);
  or _57206_ (_05461_, _05459_, _05455_);
  and _57207_ (_05462_, _04445_, _04685_);
  and _57208_ (_05463_, _04490_, _04647_);
  and _57209_ (_05465_, _04493_, _04666_);
  and _57210_ (_05466_, _04434_, _04687_);
  or _57211_ (_05467_, _05466_, _05465_);
  or _57212_ (_05469_, _05467_, _05463_);
  or _57213_ (_05470_, _05469_, _05462_);
  and _57214_ (_05471_, _04447_, _04655_);
  and _57215_ (_05473_, _04477_, _04662_);
  or _57216_ (_05474_, _05473_, _05471_);
  or _57217_ (_05475_, _05474_, _05470_);
  or _57218_ (_05477_, _05475_, _05461_);
  or _57219_ (_05478_, _05477_, _05454_);
  or _57220_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05478_, _05447_);
  and _57221_ (_05480_, _04451_, _04714_);
  and _57222_ (_05481_, _04441_, _04726_);
  and _57223_ (_05482_, _04454_, _04697_);
  or _57224_ (_05484_, _05482_, _05481_);
  or _57225_ (_05485_, _05484_, _05480_);
  and _57226_ (_05486_, _04461_, _04703_);
  and _57227_ (_05488_, _04468_, _04731_);
  or _57228_ (_05489_, _05488_, _05486_);
  and _57229_ (_05490_, _04464_, _04724_);
  and _57230_ (_05491_, _04471_, _04695_);
  or _57231_ (_05492_, _05491_, _05490_);
  or _57232_ (_05493_, _05492_, _05489_);
  and _57233_ (_05494_, _04487_, _04712_);
  and _57234_ (_05495_, _04447_, _04706_);
  and _57235_ (_05496_, _04477_, _04708_);
  or _57236_ (_05497_, _05496_, _05495_);
  or _57237_ (_05498_, _05497_, _05494_);
  and _57238_ (_05499_, _04482_, _04722_);
  and _57239_ (_05500_, _04490_, _04693_);
  and _57240_ (_05501_, _04493_, _04720_);
  and _57241_ (_05502_, _04434_, _04733_);
  or _57242_ (_05503_, _05502_, _05501_);
  or _57243_ (_05504_, _05503_, _05500_);
  or _57244_ (_05505_, _05504_, _05499_);
  and _57245_ (_05506_, _04445_, _04716_);
  and _57246_ (_05507_, _04503_, _04701_);
  or _57247_ (_05508_, _05507_, _05506_);
  or _57248_ (_05510_, _05508_, _05505_);
  or _57249_ (_05511_, _05510_, _05498_);
  or _57250_ (_05513_, _05511_, _05493_);
  or _57251_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05513_, _05485_);
  and _57252_ (_05514_, _04441_, _04777_);
  and _57253_ (_05516_, _04451_, _04760_);
  and _57254_ (_05517_, _04454_, _04743_);
  or _57255_ (_05518_, _05517_, _05516_);
  or _57256_ (_05520_, _05518_, _05514_);
  and _57257_ (_05521_, _04461_, _04749_);
  and _57258_ (_05522_, _04464_, _04775_);
  or _57259_ (_05524_, _05522_, _05521_);
  and _57260_ (_05525_, _04468_, _04766_);
  and _57261_ (_05526_, _04471_, _04741_);
  or _57262_ (_05528_, _05526_, _05525_);
  or _57263_ (_05529_, _05528_, _05524_);
  and _57264_ (_05530_, _04477_, _04754_);
  and _57265_ (_05532_, _04447_, _04752_);
  and _57266_ (_05533_, _04482_, _04773_);
  or _57267_ (_05534_, _05533_, _05532_);
  or _57268_ (_05536_, _05534_, _05530_);
  and _57269_ (_05537_, _04487_, _04758_);
  and _57270_ (_05538_, _04490_, _04739_);
  and _57271_ (_05540_, _04493_, _04768_);
  and _57272_ (_05541_, _04434_, _04771_);
  or _57273_ (_05542_, _05541_, _05540_);
  or _57274_ (_05543_, _05542_, _05538_);
  or _57275_ (_05544_, _05543_, _05537_);
  and _57276_ (_05545_, _04445_, _04762_);
  and _57277_ (_05546_, _04503_, _04747_);
  or _57278_ (_05547_, _05546_, _05545_);
  or _57279_ (_05548_, _05547_, _05544_);
  or _57280_ (_05549_, _05548_, _05536_);
  or _57281_ (_05550_, _05549_, _05529_);
  or _57282_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05550_, _05520_);
  and _57283_ (_05551_, _04451_, _04812_);
  and _57284_ (_05552_, _04441_, _04818_);
  and _57285_ (_05553_, _04454_, _04789_);
  or _57286_ (_05554_, _05553_, _05552_);
  or _57287_ (_05555_, _05554_, _05551_);
  and _57288_ (_05556_, _04461_, _04798_);
  and _57289_ (_05557_, _04464_, _04816_);
  or _57290_ (_05558_, _05557_, _05556_);
  and _57291_ (_05559_, _04468_, _04825_);
  and _57292_ (_05561_, _04471_, _04785_);
  or _57293_ (_05562_, _05561_, _05559_);
  or _57294_ (_05564_, _05562_, _05558_);
  and _57295_ (_05565_, _04487_, _04804_);
  and _57296_ (_05566_, _04447_, _04793_);
  and _57297_ (_05568_, _04477_, _04800_);
  or _57298_ (_05569_, _05568_, _05566_);
  or _57299_ (_05570_, _05569_, _05565_);
  and _57300_ (_05572_, _04482_, _04814_);
  and _57301_ (_05573_, _04490_, _04787_);
  and _57302_ (_05574_, _04493_, _04806_);
  and _57303_ (_05576_, _04434_, _04809_);
  or _57304_ (_05577_, _05576_, _05574_);
  or _57305_ (_05578_, _05577_, _05573_);
  or _57306_ (_05580_, _05578_, _05572_);
  and _57307_ (_05581_, _04445_, _04823_);
  and _57308_ (_05582_, _04503_, _04795_);
  or _57309_ (_05584_, _05582_, _05581_);
  or _57310_ (_05585_, _05584_, _05580_);
  or _57311_ (_05586_, _05585_, _05570_);
  or _57312_ (_05588_, _05586_, _05564_);
  or _57313_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05588_, _05555_);
  and _57314_ (_05589_, _04451_, _04858_);
  and _57315_ (_05591_, _04454_, _04835_);
  and _57316_ (_05592_, _04441_, _04864_);
  or _57317_ (_05593_, _05592_, _05591_);
  or _57318_ (_05594_, _05593_, _05589_);
  and _57319_ (_05595_, _04468_, _04871_);
  and _57320_ (_05596_, _04464_, _04862_);
  or _57321_ (_05597_, _05596_, _05595_);
  and _57322_ (_05598_, _04461_, _04844_);
  and _57323_ (_05599_, _04471_, _04831_);
  or _57324_ (_05600_, _05599_, _05598_);
  or _57325_ (_05601_, _05600_, _05597_);
  and _57326_ (_05602_, _04482_, _04860_);
  and _57327_ (_05603_, _04445_, _04869_);
  and _57328_ (_05604_, _04487_, _04850_);
  or _57329_ (_05605_, _05604_, _05603_);
  or _57330_ (_05606_, _05605_, _05602_);
  and _57331_ (_05607_, _04447_, _04839_);
  and _57332_ (_05608_, _04490_, _04833_);
  and _57333_ (_05609_, _04493_, _04852_);
  and _57334_ (_05610_, _04434_, _04855_);
  or _57335_ (_05611_, _05610_, _05609_);
  or _57336_ (_05613_, _05611_, _05608_);
  or _57337_ (_05614_, _05613_, _05607_);
  and _57338_ (_05616_, _04503_, _04841_);
  and _57339_ (_05617_, _04477_, _04846_);
  or _57340_ (_05618_, _05617_, _05616_);
  or _57341_ (_05620_, _05618_, _05614_);
  or _57342_ (_05621_, _05620_, _05606_);
  or _57343_ (_05622_, _05621_, _05601_);
  or _57344_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05622_, _05594_);
  and _57345_ (_05624_, _04451_, _04898_);
  and _57346_ (_05625_, _04454_, _04881_);
  and _57347_ (_05627_, _04441_, _04915_);
  or _57348_ (_05628_, _05627_, _05625_);
  or _57349_ (_05629_, _05628_, _05624_);
  and _57350_ (_05631_, _04468_, _04904_);
  and _57351_ (_05632_, _04464_, _04913_);
  or _57352_ (_05633_, _05632_, _05631_);
  and _57353_ (_05635_, _04461_, _04887_);
  and _57354_ (_05636_, _04471_, _04879_);
  or _57355_ (_05637_, _05636_, _05635_);
  or _57356_ (_05639_, _05637_, _05633_);
  and _57357_ (_05640_, _04482_, _04911_);
  and _57358_ (_05641_, _04445_, _04900_);
  and _57359_ (_05643_, _04487_, _04896_);
  or _57360_ (_05644_, _05643_, _05641_);
  or _57361_ (_05645_, _05644_, _05640_);
  and _57362_ (_05646_, _04447_, _04890_);
  and _57363_ (_05647_, _04490_, _04877_);
  and _57364_ (_05648_, _04493_, _04906_);
  and _57365_ (_05649_, _04434_, _04909_);
  or _57366_ (_05650_, _05649_, _05648_);
  or _57367_ (_05651_, _05650_, _05647_);
  or _57368_ (_05652_, _05651_, _05646_);
  and _57369_ (_05653_, _04503_, _04885_);
  and _57370_ (_05654_, _04477_, _04892_);
  or _57371_ (_05655_, _05654_, _05653_);
  or _57372_ (_05656_, _05655_, _05652_);
  or _57373_ (_05657_, _05656_, _05645_);
  or _57374_ (_05658_, _05657_, _05639_);
  or _57375_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05658_, _05629_);
  not _57376_ (_05659_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand _57377_ (_05660_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _57378_ (_05661_, \oc8051_golden_model_1.PC [3]);
  or _57379_ (_05662_, \oc8051_golden_model_1.PC [2], _05661_);
  or _57380_ (_05664_, _05662_, _05660_);
  or _57381_ (_05665_, _05664_, _00548_);
  not _57382_ (_05667_, \oc8051_golden_model_1.PC [1]);
  or _57383_ (_05668_, _05667_, \oc8051_golden_model_1.PC [0]);
  or _57384_ (_05669_, _05668_, _05662_);
  or _57385_ (_05671_, _05669_, _00507_);
  and _57386_ (_05672_, _05671_, _05665_);
  not _57387_ (_05673_, \oc8051_golden_model_1.PC [2]);
  or _57388_ (_05675_, _05673_, \oc8051_golden_model_1.PC [3]);
  or _57389_ (_05676_, _05675_, _05660_);
  or _57390_ (_05677_, _05676_, _00384_);
  or _57391_ (_05679_, _05675_, _05668_);
  or _57392_ (_05680_, _05679_, _00343_);
  and _57393_ (_05681_, _05680_, _05677_);
  and _57394_ (_05683_, _05681_, _05672_);
  nand _57395_ (_05684_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _57396_ (_05685_, _05684_, _05660_);
  or _57397_ (_05687_, _05685_, _00731_);
  or _57398_ (_05688_, _05684_, _05668_);
  or _57399_ (_05689_, _05688_, _00690_);
  and _57400_ (_05691_, _05689_, _05687_);
  or _57401_ (_05692_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _57402_ (_05693_, _05692_, _05660_);
  or _57403_ (_05695_, _05693_, _00220_);
  or _57404_ (_05696_, _05692_, _05668_);
  or _57405_ (_05697_, _05696_, _00162_);
  and _57406_ (_05698_, _05697_, _05695_);
  and _57407_ (_05699_, _05698_, _05691_);
  and _57408_ (_05700_, _05699_, _05683_);
  not _57409_ (_05701_, \oc8051_golden_model_1.PC [0]);
  or _57410_ (_05702_, \oc8051_golden_model_1.PC [1], _05701_);
  or _57411_ (_05703_, _05702_, _05684_);
  or _57412_ (_05704_, _05703_, _00649_);
  or _57413_ (_05705_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _57414_ (_05706_, _05705_, _05684_);
  or _57415_ (_05707_, _05706_, _00608_);
  and _57416_ (_05708_, _05707_, _05704_);
  or _57417_ (_05709_, _05692_, _05705_);
  or _57418_ (_05710_, _05709_, _00066_);
  or _57419_ (_05711_, _05692_, _05702_);
  or _57420_ (_05712_, _05711_, _00107_);
  and _57421_ (_05713_, _05712_, _05710_);
  and _57422_ (_05714_, _05713_, _05708_);
  or _57423_ (_05715_, _05702_, _05662_);
  or _57424_ (_05717_, _05715_, _00466_);
  or _57425_ (_05718_, _05705_, _05662_);
  or _57426_ (_05720_, _05718_, _00425_);
  and _57427_ (_05721_, _05720_, _05717_);
  or _57428_ (_05722_, _05702_, _05675_);
  or _57429_ (_05724_, _05722_, _00302_);
  or _57430_ (_05725_, _05705_, _05675_);
  or _57431_ (_05726_, _05725_, _00261_);
  and _57432_ (_05728_, _05726_, _05724_);
  and _57433_ (_05729_, _05728_, _05721_);
  and _57434_ (_05730_, _05729_, _05714_);
  nand _57435_ (_05732_, _05730_, _05700_);
  or _57436_ (_05733_, _05664_, _00513_);
  or _57437_ (_05734_, _05669_, _00472_);
  and _57438_ (_05736_, _05734_, _05733_);
  or _57439_ (_05737_, _05676_, _00349_);
  or _57440_ (_05738_, _05679_, _00308_);
  and _57441_ (_05740_, _05738_, _05737_);
  and _57442_ (_05741_, _05740_, _05736_);
  or _57443_ (_05742_, _05685_, _00696_);
  or _57444_ (_05744_, _05688_, _00655_);
  and _57445_ (_05745_, _05744_, _05742_);
  or _57446_ (_05746_, _05693_, _00175_);
  or _57447_ (_05748_, _05696_, _00113_);
  and _57448_ (_05749_, _05748_, _05746_);
  and _57449_ (_05750_, _05749_, _05745_);
  and _57450_ (_05751_, _05750_, _05741_);
  or _57451_ (_05752_, _05703_, _00614_);
  or _57452_ (_05753_, _05706_, _00557_);
  and _57453_ (_05754_, _05753_, _05752_);
  or _57454_ (_05755_, _05709_, _00031_);
  or _57455_ (_05756_, _05711_, _00072_);
  and _57456_ (_05757_, _05756_, _05755_);
  and _57457_ (_05758_, _05757_, _05754_);
  or _57458_ (_05759_, _05715_, _00431_);
  or _57459_ (_05760_, _05718_, _00390_);
  and _57460_ (_05761_, _05760_, _05759_);
  or _57461_ (_05762_, _05722_, _00267_);
  or _57462_ (_05763_, _05725_, _00226_);
  and _57463_ (_05764_, _05763_, _05762_);
  and _57464_ (_05765_, _05764_, _05761_);
  and _57465_ (_05766_, _05765_, _05758_);
  nand _57466_ (_05767_, _05766_, _05751_);
  or _57467_ (_05768_, _05767_, _05732_);
  or _57468_ (_05770_, _05664_, _00538_);
  or _57469_ (_05771_, _05669_, _00497_);
  and _57470_ (_05773_, _05771_, _05770_);
  or _57471_ (_05774_, _05676_, _00374_);
  or _57472_ (_05775_, _05679_, _00333_);
  and _57473_ (_05777_, _05775_, _05774_);
  and _57474_ (_05778_, _05777_, _05773_);
  or _57475_ (_05779_, _05685_, _00721_);
  or _57476_ (_05781_, _05688_, _00680_);
  and _57477_ (_05782_, _05781_, _05779_);
  or _57478_ (_05783_, _05693_, _00210_);
  or _57479_ (_05785_, _05696_, _00140_);
  and _57480_ (_05786_, _05785_, _05783_);
  and _57481_ (_05787_, _05786_, _05782_);
  and _57482_ (_05789_, _05787_, _05778_);
  or _57483_ (_05790_, _05703_, _00639_);
  or _57484_ (_05791_, _05706_, _00597_);
  and _57485_ (_05793_, _05791_, _05790_);
  or _57486_ (_05794_, _05709_, _00056_);
  or _57487_ (_05795_, _05711_, _00097_);
  and _57488_ (_05797_, _05795_, _05794_);
  and _57489_ (_05798_, _05797_, _05793_);
  or _57490_ (_05799_, _05715_, _00456_);
  or _57491_ (_05801_, _05718_, _00415_);
  and _57492_ (_05802_, _05801_, _05799_);
  or _57493_ (_05803_, _05722_, _00292_);
  or _57494_ (_05804_, _05725_, _00251_);
  and _57495_ (_05805_, _05804_, _05803_);
  and _57496_ (_05806_, _05805_, _05802_);
  and _57497_ (_05807_, _05806_, _05798_);
  nand _57498_ (_05808_, _05807_, _05789_);
  or _57499_ (_05809_, _05664_, _00543_);
  or _57500_ (_05810_, _05669_, _00502_);
  and _57501_ (_05811_, _05810_, _05809_);
  or _57502_ (_05812_, _05676_, _00379_);
  or _57503_ (_05813_, _05679_, _00338_);
  and _57504_ (_05814_, _05813_, _05812_);
  and _57505_ (_05815_, _05814_, _05811_);
  or _57506_ (_05816_, _05685_, _00726_);
  or _57507_ (_05817_, _05688_, _00685_);
  and _57508_ (_05818_, _05817_, _05816_);
  or _57509_ (_05819_, _05693_, _00215_);
  or _57510_ (_05820_, _05696_, _00151_);
  and _57511_ (_05821_, _05820_, _05819_);
  and _57512_ (_05823_, _05821_, _05818_);
  and _57513_ (_05824_, _05823_, _05815_);
  or _57514_ (_05826_, _05703_, _00644_);
  or _57515_ (_05827_, _05706_, _00603_);
  and _57516_ (_05828_, _05827_, _05826_);
  or _57517_ (_05830_, _05709_, _00061_);
  or _57518_ (_05831_, _05711_, _00102_);
  and _57519_ (_05832_, _05831_, _05830_);
  and _57520_ (_05834_, _05832_, _05828_);
  or _57521_ (_05835_, _05715_, _00461_);
  or _57522_ (_05836_, _05718_, _00420_);
  and _57523_ (_05838_, _05836_, _05835_);
  or _57524_ (_05839_, _05722_, _00297_);
  or _57525_ (_05840_, _05725_, _00256_);
  and _57526_ (_05842_, _05840_, _05839_);
  and _57527_ (_05843_, _05842_, _05838_);
  and _57528_ (_05844_, _05843_, _05834_);
  and _57529_ (_05846_, _05844_, _05824_);
  nand _57530_ (_05847_, _05846_, _05808_);
  nor _57531_ (_05848_, _05847_, _05768_);
  or _57532_ (_05850_, _05664_, _00518_);
  or _57533_ (_05851_, _05669_, _00477_);
  and _57534_ (_05852_, _05851_, _05850_);
  or _57535_ (_05854_, _05676_, _00354_);
  or _57536_ (_05855_, _05679_, _00313_);
  and _57537_ (_05856_, _05855_, _05854_);
  and _57538_ (_05857_, _05856_, _05852_);
  or _57539_ (_05858_, _05685_, _00701_);
  or _57540_ (_05859_, _05688_, _00660_);
  and _57541_ (_05860_, _05859_, _05858_);
  or _57542_ (_05861_, _05693_, _00186_);
  or _57543_ (_05862_, _05696_, _00118_);
  and _57544_ (_05863_, _05862_, _05861_);
  and _57545_ (_05864_, _05863_, _05860_);
  and _57546_ (_05865_, _05864_, _05857_);
  or _57547_ (_05866_, _05703_, _00619_);
  or _57548_ (_05867_, _05706_, _00565_);
  and _57549_ (_05868_, _05867_, _05866_);
  or _57550_ (_05869_, _05709_, _00036_);
  or _57551_ (_05870_, _05711_, _00077_);
  and _57552_ (_05871_, _05870_, _05869_);
  and _57553_ (_05872_, _05871_, _05868_);
  or _57554_ (_05873_, _05715_, _00436_);
  or _57555_ (_05874_, _05718_, _00395_);
  and _57556_ (_05876_, _05874_, _05873_);
  or _57557_ (_05877_, _05722_, _00272_);
  or _57558_ (_05879_, _05725_, _00231_);
  and _57559_ (_05880_, _05879_, _05877_);
  and _57560_ (_05881_, _05880_, _05876_);
  and _57561_ (_05883_, _05881_, _05872_);
  and _57562_ (_05884_, _05883_, _05865_);
  or _57563_ (_05885_, _05664_, _00523_);
  or _57564_ (_05887_, _05669_, _00482_);
  and _57565_ (_05888_, _05887_, _05885_);
  or _57566_ (_05889_, _05676_, _00359_);
  or _57567_ (_05891_, _05679_, _00318_);
  and _57568_ (_05892_, _05891_, _05889_);
  and _57569_ (_05893_, _05892_, _05888_);
  or _57570_ (_05895_, _05685_, _00706_);
  or _57571_ (_05896_, _05688_, _00665_);
  and _57572_ (_05897_, _05896_, _05895_);
  or _57573_ (_05899_, _05693_, _00195_);
  or _57574_ (_05900_, _05696_, _00123_);
  and _57575_ (_05901_, _05900_, _05899_);
  and _57576_ (_05903_, _05901_, _05897_);
  and _57577_ (_05904_, _05903_, _05893_);
  or _57578_ (_05905_, _05703_, _00624_);
  or _57579_ (_05907_, _05706_, _00573_);
  and _57580_ (_05908_, _05907_, _05905_);
  or _57581_ (_05909_, _05709_, _00041_);
  or _57582_ (_05910_, _05711_, _00082_);
  and _57583_ (_05911_, _05910_, _05909_);
  and _57584_ (_05912_, _05911_, _05908_);
  or _57585_ (_05913_, _05715_, _00441_);
  or _57586_ (_05914_, _05718_, _00400_);
  and _57587_ (_05915_, _05914_, _05913_);
  or _57588_ (_05916_, _05722_, _00277_);
  or _57589_ (_05917_, _05725_, _00236_);
  and _57590_ (_05918_, _05917_, _05916_);
  and _57591_ (_05919_, _05918_, _05915_);
  and _57592_ (_05920_, _05919_, _05912_);
  nand _57593_ (_05921_, _05920_, _05904_);
  not _57594_ (_05922_, _05921_);
  and _57595_ (_05923_, _05922_, _05884_);
  or _57596_ (_05924_, _05664_, _00528_);
  or _57597_ (_05925_, _05669_, _00487_);
  and _57598_ (_05926_, _05925_, _05924_);
  or _57599_ (_05927_, _05676_, _00364_);
  or _57600_ (_05928_, _05679_, _00323_);
  and _57601_ (_05929_, _05928_, _05927_);
  and _57602_ (_05930_, _05929_, _05926_);
  or _57603_ (_05931_, _05685_, _00711_);
  or _57604_ (_05932_, _05688_, _00670_);
  and _57605_ (_05933_, _05932_, _05931_);
  or _57606_ (_05934_, _05693_, _00200_);
  or _57607_ (_05935_, _05696_, _00128_);
  and _57608_ (_05936_, _05935_, _05934_);
  and _57609_ (_05937_, _05936_, _05933_);
  and _57610_ (_05938_, _05937_, _05930_);
  or _57611_ (_05939_, _05703_, _00629_);
  or _57612_ (_05940_, _05706_, _00581_);
  and _57613_ (_05941_, _05940_, _05939_);
  or _57614_ (_05942_, _05709_, _00046_);
  or _57615_ (_05943_, _05711_, _00087_);
  and _57616_ (_05944_, _05943_, _05942_);
  and _57617_ (_05945_, _05944_, _05941_);
  or _57618_ (_05946_, _05715_, _00446_);
  or _57619_ (_05947_, _05718_, _00405_);
  and _57620_ (_05948_, _05947_, _05946_);
  or _57621_ (_05949_, _05722_, _00282_);
  or _57622_ (_05950_, _05725_, _00241_);
  and _57623_ (_05951_, _05950_, _05949_);
  and _57624_ (_05952_, _05951_, _05948_);
  and _57625_ (_05953_, _05952_, _05945_);
  nand _57626_ (_05954_, _05953_, _05938_);
  or _57627_ (_05955_, _05664_, _00533_);
  or _57628_ (_05956_, _05669_, _00492_);
  and _57629_ (_05957_, _05956_, _05955_);
  or _57630_ (_05958_, _05676_, _00369_);
  or _57631_ (_05959_, _05679_, _00328_);
  and _57632_ (_05960_, _05959_, _05958_);
  and _57633_ (_05961_, _05960_, _05957_);
  or _57634_ (_05962_, _05685_, _00716_);
  or _57635_ (_05963_, _05688_, _00675_);
  and _57636_ (_05964_, _05963_, _05962_);
  or _57637_ (_05965_, _05693_, _00205_);
  or _57638_ (_05966_, _05696_, _00133_);
  and _57639_ (_05967_, _05966_, _05965_);
  and _57640_ (_05968_, _05967_, _05964_);
  and _57641_ (_05969_, _05968_, _05961_);
  or _57642_ (_05970_, _05703_, _00634_);
  or _57643_ (_05971_, _05706_, _00589_);
  and _57644_ (_05972_, _05971_, _05970_);
  or _57645_ (_05973_, _05709_, _00051_);
  or _57646_ (_05974_, _05711_, _00092_);
  and _57647_ (_05975_, _05974_, _05973_);
  and _57648_ (_05976_, _05975_, _05972_);
  or _57649_ (_05977_, _05715_, _00451_);
  or _57650_ (_05978_, _05718_, _00410_);
  and _57651_ (_05979_, _05978_, _05977_);
  or _57652_ (_05980_, _05722_, _00287_);
  or _57653_ (_05981_, _05725_, _00246_);
  and _57654_ (_05982_, _05981_, _05980_);
  and _57655_ (_05983_, _05982_, _05979_);
  and _57656_ (_05984_, _05983_, _05976_);
  nand _57657_ (_05985_, _05984_, _05969_);
  or _57658_ (_05986_, _05985_, _05954_);
  not _57659_ (_05987_, _05986_);
  and _57660_ (_05988_, _05987_, _05923_);
  and _57661_ (_05989_, _05988_, _05848_);
  not _57662_ (_05990_, _05989_);
  or _57663_ (_05991_, _05921_, _05884_);
  or _57664_ (_05992_, _05991_, _05986_);
  not _57665_ (_05993_, _05992_);
  and _57666_ (_05994_, _05807_, _05789_);
  nand _57667_ (_05995_, _05846_, _05994_);
  nor _57668_ (_05996_, _05995_, _05768_);
  and _57669_ (_05997_, _05996_, _05993_);
  and _57670_ (_05998_, _05993_, _05848_);
  nor _57671_ (_05999_, _05998_, _05997_);
  and _57672_ (_06000_, _05766_, _05751_);
  or _57673_ (_06001_, _06000_, _05732_);
  nor _57674_ (_06002_, _06001_, _05995_);
  not _57675_ (_06003_, _06002_);
  or _57676_ (_06004_, _06003_, _05992_);
  and _57677_ (_06005_, _05730_, _05700_);
  or _57678_ (_06006_, _05767_, _06005_);
  or _57679_ (_06007_, _05846_, _05994_);
  or _57680_ (_06008_, _06007_, _06006_);
  or _57681_ (_06009_, _06008_, _05992_);
  or _57682_ (_06010_, _05846_, _05808_);
  or _57683_ (_06011_, _06006_, _06010_);
  or _57684_ (_06012_, _06011_, _05992_);
  and _57685_ (_06013_, _06012_, _06009_);
  and _57686_ (_06014_, _06013_, _06004_);
  or _57687_ (_06015_, _06007_, _05768_);
  or _57688_ (_06016_, _06015_, _05992_);
  or _57689_ (_06017_, _06006_, _05847_);
  or _57690_ (_06018_, _06017_, _05992_);
  and _57691_ (_06019_, _06018_, _06016_);
  or _57692_ (_06020_, _06010_, _05768_);
  or _57693_ (_06021_, _06020_, _05992_);
  or _57694_ (_06022_, _06006_, _05995_);
  or _57695_ (_06023_, _06022_, _05992_);
  and _57696_ (_06024_, _06023_, _06021_);
  and _57697_ (_06025_, _06024_, _06019_);
  and _57698_ (_06026_, _06025_, _06014_);
  and _57699_ (_06027_, _06026_, _05999_);
  not _57700_ (_06028_, _05884_);
  and _57701_ (_06029_, _05921_, _06028_);
  and _57702_ (_06030_, _06029_, _05987_);
  and _57703_ (_06031_, _06030_, _06002_);
  not _57704_ (_06032_, _06031_);
  not _57705_ (_06033_, _05991_);
  not _57706_ (_06034_, _05985_);
  and _57707_ (_06035_, _06034_, _05954_);
  and _57708_ (_06036_, _06035_, _06033_);
  and _57709_ (_06037_, _06036_, _06002_);
  nor _57710_ (_06038_, _06001_, _05847_);
  and _57711_ (_06039_, _06038_, _05993_);
  nor _57712_ (_06040_, _06039_, _06037_);
  and _57713_ (_06041_, _06040_, _06032_);
  and _57714_ (_06042_, _06038_, _06030_);
  not _57715_ (_06043_, _06042_);
  and _57716_ (_06044_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _57717_ (_06045_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _57718_ (_06046_, _06045_, _06044_);
  or _57719_ (_06047_, _06046_, _06043_);
  or _57720_ (_06048_, _06001_, _06007_);
  or _57721_ (_06049_, _06048_, _05992_);
  or _57722_ (_06050_, _06000_, _06005_);
  or _57723_ (_06051_, _06050_, _05847_);
  or _57724_ (_06052_, _06051_, _05992_);
  and _57725_ (_06053_, _06052_, _06049_);
  or _57726_ (_06054_, _06001_, _06010_);
  or _57727_ (_06055_, _06054_, _05992_);
  or _57728_ (_06056_, _06050_, _05995_);
  or _57729_ (_06057_, _06056_, _05992_);
  and _57730_ (_06058_, _06057_, _06055_);
  or _57731_ (_06059_, _06050_, _06007_);
  or _57732_ (_06060_, _06059_, _05992_);
  or _57733_ (_06061_, _06050_, _06010_);
  or _57734_ (_06062_, _06061_, _05992_);
  and _57735_ (_06063_, _06062_, _06060_);
  and _57736_ (_06064_, _06063_, _06058_);
  and _57737_ (_06065_, _06064_, _06053_);
  nor _57738_ (_06066_, _06042_, _05701_);
  nand _57739_ (_06067_, _06066_, _06065_);
  nand _57740_ (_06068_, _06067_, _06047_);
  and _57741_ (_06069_, _06068_, _06041_);
  and _57742_ (_06070_, \oc8051_golden_model_1.ACC [0], _05701_);
  not _57743_ (_06071_, \oc8051_golden_model_1.ACC [0]);
  and _57744_ (_06072_, _06071_, \oc8051_golden_model_1.PC [0]);
  nor _57745_ (_06073_, _06072_, _06070_);
  nor _57746_ (_06074_, _06073_, _06032_);
  or _57747_ (_06075_, _06074_, _06069_);
  nand _57748_ (_06076_, _06075_, _06027_);
  and _57749_ (_06077_, _06065_, _06040_);
  and _57750_ (_06078_, _06077_, _06027_);
  or _57751_ (_06079_, _06078_, \oc8051_golden_model_1.PC [0]);
  nand _57752_ (_06080_, _06079_, _06076_);
  or _57753_ (_06081_, _06077_, \oc8051_golden_model_1.PC [1]);
  and _57754_ (_06082_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _57755_ (_06083_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _57756_ (_06084_, _06083_, _06082_);
  and _57757_ (_06085_, _06084_, _06044_);
  nor _57758_ (_06086_, _06084_, _06044_);
  nor _57759_ (_06087_, _06086_, _06085_);
  nand _57760_ (_06088_, _06087_, _06042_);
  and _57761_ (_06089_, _05702_, _05668_);
  nor _57762_ (_06090_, _06089_, _06042_);
  nand _57763_ (_06091_, _06090_, _06065_);
  nand _57764_ (_06092_, _06091_, _06088_);
  and _57765_ (_06093_, _06040_, _06027_);
  nand _57766_ (_06094_, _06093_, _06092_);
  nand _57767_ (_06095_, _06094_, _06081_);
  nand _57768_ (_06096_, _06095_, _06032_);
  not _57769_ (_06097_, \oc8051_golden_model_1.ACC [1]);
  nor _57770_ (_06098_, _06089_, _06097_);
  and _57771_ (_06099_, _06089_, _06097_);
  nor _57772_ (_06100_, _06099_, _06098_);
  and _57773_ (_06101_, _06100_, _06070_);
  nor _57774_ (_06102_, _06100_, _06070_);
  nor _57775_ (_06103_, _06102_, _06101_);
  and _57776_ (_06104_, _06103_, _06031_);
  nor _57777_ (_06105_, _06027_, \oc8051_golden_model_1.PC [1]);
  nor _57778_ (_06106_, _06105_, _06104_);
  and _57779_ (_06107_, _06106_, _06096_);
  or _57780_ (_06108_, _06107_, _06080_);
  and _57781_ (_06109_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _57782_ (_06110_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _57783_ (_06111_, _06110_, _06109_);
  or _57784_ (_06112_, _06111_, _06027_);
  not _57785_ (_06113_, _06111_);
  or _57786_ (_06114_, _06113_, _06077_);
  nor _57787_ (_06115_, _06085_, _06082_);
  and _57788_ (_06116_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _57789_ (_06117_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _57790_ (_06118_, _06117_, _06116_);
  not _57791_ (_06119_, _06118_);
  nor _57792_ (_06120_, _06119_, _06115_);
  and _57793_ (_06121_, _06119_, _06115_);
  nor _57794_ (_06122_, _06121_, _06120_);
  nand _57795_ (_06123_, _06122_, _06042_);
  nand _57796_ (_06124_, _06064_, _06053_);
  nor _57797_ (_06125_, _05660_, _05673_);
  and _57798_ (_06126_, _05660_, _05673_);
  nor _57799_ (_06127_, _06126_, _06125_);
  not _57800_ (_06128_, _06127_);
  or _57801_ (_06129_, _06128_, _06042_);
  or _57802_ (_06130_, _06129_, _06124_);
  nand _57803_ (_06131_, _06130_, _06123_);
  nand _57804_ (_06132_, _06131_, _06040_);
  and _57805_ (_06133_, _06132_, _06114_);
  or _57806_ (_06134_, _06133_, _06031_);
  nor _57807_ (_06135_, _06101_, _06098_);
  and _57808_ (_06136_, _06127_, \oc8051_golden_model_1.ACC [2]);
  nor _57809_ (_06137_, _06127_, \oc8051_golden_model_1.ACC [2]);
  nor _57810_ (_06138_, _06137_, _06136_);
  not _57811_ (_06139_, _06138_);
  and _57812_ (_06140_, _06139_, _06135_);
  nor _57813_ (_06141_, _06139_, _06135_);
  nor _57814_ (_06142_, _06141_, _06140_);
  and _57815_ (_06143_, _06142_, _06031_);
  not _57816_ (_06144_, _06143_);
  and _57817_ (_06145_, _06144_, _06027_);
  nand _57818_ (_06146_, _06145_, _06134_);
  nand _57819_ (_06147_, _06146_, _06112_);
  nor _57820_ (_06148_, _05684_, _05667_);
  nor _57821_ (_06149_, _06109_, \oc8051_golden_model_1.PC [3]);
  nor _57822_ (_06150_, _06149_, _06148_);
  or _57823_ (_06151_, _06150_, _06078_);
  nor _57824_ (_06152_, _06141_, _06136_);
  not _57825_ (_06153_, _05676_);
  nor _57826_ (_06154_, _06125_, _05661_);
  nor _57827_ (_06155_, _06154_, _06153_);
  nor _57828_ (_06156_, _06155_, \oc8051_golden_model_1.ACC [3]);
  and _57829_ (_06157_, _06155_, \oc8051_golden_model_1.ACC [3]);
  nor _57830_ (_06158_, _06157_, _06156_);
  and _57831_ (_06159_, _06158_, _06152_);
  nor _57832_ (_06160_, _06158_, _06152_);
  nor _57833_ (_06161_, _06160_, _06159_);
  nor _57834_ (_06162_, _06161_, _06032_);
  nor _57835_ (_06163_, _06120_, _06116_);
  and _57836_ (_06164_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _57837_ (_06165_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _57838_ (_06166_, _06165_, _06164_);
  not _57839_ (_06167_, _06166_);
  nor _57840_ (_06168_, _06167_, _06163_);
  and _57841_ (_06169_, _06167_, _06163_);
  nor _57842_ (_06170_, _06169_, _06168_);
  not _57843_ (_06171_, _06170_);
  nand _57844_ (_06172_, _06171_, _06042_);
  not _57845_ (_06173_, _06155_);
  nor _57846_ (_06174_, _06042_, _06173_);
  nand _57847_ (_06175_, _06174_, _06065_);
  nand _57848_ (_06176_, _06175_, _06172_);
  and _57849_ (_06177_, _06176_, _06041_);
  or _57850_ (_06178_, _06177_, _06162_);
  nand _57851_ (_06179_, _06178_, _06027_);
  and _57852_ (_06180_, _06179_, _06151_);
  or _57853_ (_06181_, _06180_, _06147_);
  or _57854_ (_06182_, _06181_, _06108_);
  or _57855_ (_06183_, _06182_, _00349_);
  and _57856_ (_06184_, _06079_, _06076_);
  nand _57857_ (_06185_, _06106_, _06096_);
  or _57858_ (_06186_, _06185_, _06184_);
  and _57859_ (_06187_, _06146_, _06112_);
  or _57860_ (_06188_, _06180_, _06187_);
  or _57861_ (_06189_, _06188_, _06186_);
  or _57862_ (_06190_, _06189_, _00031_);
  and _57863_ (_06191_, _06190_, _06183_);
  nand _57864_ (_06192_, _06179_, _06151_);
  or _57865_ (_06193_, _06192_, _06187_);
  or _57866_ (_06194_, _06193_, _06186_);
  or _57867_ (_06195_, _06194_, _00390_);
  or _57868_ (_06196_, _06188_, _06108_);
  or _57869_ (_06197_, _06196_, _00175_);
  and _57870_ (_06198_, _06197_, _06195_);
  and _57871_ (_06199_, _06198_, _06191_);
  or _57872_ (_06200_, _06193_, _06108_);
  or _57873_ (_06201_, _06200_, _00513_);
  or _57874_ (_06202_, _06185_, _06080_);
  or _57875_ (_06203_, _06202_, _06188_);
  or _57876_ (_06204_, _06203_, _00072_);
  and _57877_ (_06205_, _06204_, _06201_);
  or _57878_ (_06206_, _06192_, _06147_);
  or _57879_ (_06207_, _06206_, _06202_);
  or _57880_ (_06208_, _06207_, _00614_);
  or _57881_ (_06209_, _06206_, _06186_);
  or _57882_ (_06210_, _06209_, _00557_);
  and _57883_ (_06211_, _06210_, _06208_);
  and _57884_ (_06212_, _06211_, _06205_);
  and _57885_ (_06213_, _06212_, _06199_);
  or _57886_ (_06214_, _06107_, _06184_);
  or _57887_ (_06215_, _06214_, _06206_);
  or _57888_ (_06216_, _06215_, _00655_);
  or _57889_ (_06217_, _06214_, _06188_);
  or _57890_ (_06218_, _06217_, _00113_);
  and _57891_ (_06219_, _06218_, _06216_);
  or _57892_ (_06220_, _06202_, _06193_);
  or _57893_ (_06221_, _06220_, _00431_);
  or _57894_ (_06222_, _06214_, _06181_);
  or _57895_ (_06223_, _06222_, _00308_);
  and _57896_ (_06224_, _06223_, _06221_);
  and _57897_ (_06225_, _06224_, _06219_);
  or _57898_ (_06226_, _06214_, _06193_);
  or _57899_ (_06227_, _06226_, _00472_);
  or _57900_ (_06228_, _06186_, _06181_);
  or _57901_ (_06229_, _06228_, _00226_);
  and _57902_ (_06230_, _06229_, _06227_);
  or _57903_ (_06231_, _06206_, _06108_);
  or _57904_ (_06232_, _06231_, _00696_);
  or _57905_ (_06233_, _06202_, _06181_);
  or _57906_ (_06234_, _06233_, _00267_);
  and _57907_ (_06235_, _06234_, _06232_);
  and _57908_ (_06236_, _06235_, _06230_);
  and _57909_ (_06237_, _06236_, _06225_);
  nand _57910_ (_06238_, _06237_, _06213_);
  or _57911_ (_06239_, _06215_, _00675_);
  or _57912_ (_06240_, _06207_, _00634_);
  and _57913_ (_06241_, _06240_, _06239_);
  or _57914_ (_06242_, _06189_, _00051_);
  or _57915_ (_06243_, _06217_, _00133_);
  and _57916_ (_06244_, _06243_, _06242_);
  and _57917_ (_06245_, _06244_, _06241_);
  or _57918_ (_06246_, _06200_, _00533_);
  or _57919_ (_06247_, _06220_, _00451_);
  and _57920_ (_06248_, _06247_, _06246_);
  or _57921_ (_06249_, _06233_, _00287_);
  or _57922_ (_06250_, _06203_, _00092_);
  and _57923_ (_06251_, _06250_, _06249_);
  and _57924_ (_06252_, _06251_, _06248_);
  and _57925_ (_06253_, _06252_, _06245_);
  or _57926_ (_06254_, _06222_, _00328_);
  or _57927_ (_06255_, _06228_, _00246_);
  and _57928_ (_06256_, _06255_, _06254_);
  or _57929_ (_06257_, _06231_, _00716_);
  or _57930_ (_06258_, _06209_, _00589_);
  and _57931_ (_06259_, _06258_, _06257_);
  and _57932_ (_06260_, _06259_, _06256_);
  or _57933_ (_06261_, _06182_, _00369_);
  or _57934_ (_06262_, _06194_, _00410_);
  and _57935_ (_06263_, _06262_, _06261_);
  or _57936_ (_06264_, _06226_, _00492_);
  or _57937_ (_06265_, _06196_, _00205_);
  and _57938_ (_06266_, _06265_, _06264_);
  and _57939_ (_06267_, _06266_, _06263_);
  and _57940_ (_06268_, _06267_, _06260_);
  and _57941_ (_06269_, _06268_, _06253_);
  or _57942_ (_06270_, _06269_, _06238_);
  nor _57943_ (_06271_, _06270_, _05990_);
  nor _57944_ (_06272_, _06238_, _05990_);
  not _57945_ (_06273_, _06272_);
  nor _57946_ (_06274_, _06016_, \oc8051_golden_model_1.SP [0]);
  not _57947_ (_06275_, _06009_);
  not _57948_ (_06276_, _06008_);
  and _57949_ (_06277_, _06036_, _06276_);
  not _57950_ (_06278_, _06277_);
  nor _57951_ (_06279_, _06278_, _06238_);
  or _57952_ (_06280_, _06196_, _00186_);
  or _57953_ (_06281_, _06189_, _00036_);
  and _57954_ (_06282_, _06281_, _06280_);
  or _57955_ (_06283_, _06220_, _00436_);
  or _57956_ (_06284_, _06217_, _00118_);
  and _57957_ (_06285_, _06284_, _06283_);
  and _57958_ (_06286_, _06285_, _06282_);
  or _57959_ (_06287_, _06182_, _00354_);
  or _57960_ (_06288_, _06222_, _00313_);
  and _57961_ (_06289_, _06288_, _06287_);
  or _57962_ (_06290_, _06231_, _00701_);
  or _57963_ (_06291_, _06209_, _00565_);
  and _57964_ (_06292_, _06291_, _06290_);
  and _57965_ (_06293_, _06292_, _06289_);
  and _57966_ (_06294_, _06293_, _06286_);
  or _57967_ (_06295_, _06228_, _00231_);
  or _57968_ (_06296_, _06203_, _00077_);
  and _57969_ (_06297_, _06296_, _06295_);
  or _57970_ (_06298_, _06200_, _00518_);
  or _57971_ (_06299_, _06226_, _00477_);
  and _57972_ (_06300_, _06299_, _06298_);
  and _57973_ (_06301_, _06300_, _06297_);
  or _57974_ (_06302_, _06215_, _00660_);
  or _57975_ (_06303_, _06207_, _00619_);
  and _57976_ (_06304_, _06303_, _06302_);
  or _57977_ (_06305_, _06194_, _00395_);
  or _57978_ (_06306_, _06233_, _00272_);
  and _57979_ (_06307_, _06306_, _06305_);
  and _57980_ (_06308_, _06307_, _06304_);
  and _57981_ (_06309_, _06308_, _06301_);
  and _57982_ (_06310_, _06309_, _06294_);
  not _57983_ (_06311_, _06310_);
  and _57984_ (_06312_, _06311_, _06279_);
  not _57985_ (_06313_, _06037_);
  nor _57986_ (_06314_, _06034_, _05954_);
  and _57987_ (_06315_, _06314_, _05922_);
  and _57988_ (_06316_, _06315_, _06002_);
  not _57989_ (_06317_, _06316_);
  and _57990_ (_06318_, _05985_, _05954_);
  not _57991_ (_06319_, _06318_);
  or _57992_ (_06320_, _06319_, _05923_);
  nor _57993_ (_06321_, _06320_, _06003_);
  and _57994_ (_06322_, _06318_, _05923_);
  and _57995_ (_06323_, _06314_, _05921_);
  nor _57996_ (_06324_, _06323_, _06322_);
  nor _57997_ (_06325_, _06324_, _06003_);
  nor _57998_ (_06326_, _06325_, _06321_);
  and _57999_ (_06327_, _06326_, _06317_);
  and _58000_ (_06328_, _05921_, _05884_);
  and _58001_ (_06329_, _06328_, _06035_);
  and _58002_ (_06330_, _06329_, _06002_);
  and _58003_ (_06331_, _06035_, _06029_);
  and _58004_ (_06332_, _06331_, _06002_);
  nor _58005_ (_06333_, _06332_, _06330_);
  and _58006_ (_06334_, _06333_, _06327_);
  and _58007_ (_06335_, _06334_, _06313_);
  or _58008_ (_06336_, _06335_, _06238_);
  nor _58009_ (_06337_, _06336_, _06311_);
  and _58010_ (_06338_, _06328_, _05987_);
  and _58011_ (_06339_, _06338_, _06038_);
  not _58012_ (_06340_, _06339_);
  nor _58013_ (_06341_, _06340_, _06270_);
  not _58014_ (_06342_, \oc8051_golden_model_1.SP [0]);
  nor _58015_ (_06343_, _06049_, _06342_);
  not _58016_ (_06344_, _06048_);
  and _58017_ (_06345_, _06338_, _06344_);
  not _58018_ (_06346_, _06345_);
  nor _58019_ (_06347_, _06346_, _06270_);
  nor _58020_ (_06348_, _06346_, _06238_);
  not _58021_ (_06349_, _06348_);
  not _58022_ (_06350_, _06056_);
  and _58023_ (_06351_, _06350_, _05988_);
  and _58024_ (_06352_, _06338_, _06350_);
  not _58025_ (_06353_, _06352_);
  nor _58026_ (_06354_, _06353_, _06270_);
  not _58027_ (_06355_, _06051_);
  and _58028_ (_06356_, _06338_, _06355_);
  not _58029_ (_06357_, _06356_);
  or _58030_ (_06358_, _06357_, _06270_);
  not _58031_ (_06359_, _06060_);
  not _58032_ (_06360_, _06020_);
  and _58033_ (_06361_, _06338_, _06360_);
  not _58034_ (_06362_, _06361_);
  and _58035_ (_06363_, _06036_, _06360_);
  not _58036_ (_06364_, _06363_);
  and _58037_ (_06365_, _06269_, _06238_);
  not _58038_ (_06366_, _06238_);
  nor _58039_ (_06367_, _06209_, _00608_);
  nor _58040_ (_06368_, _06200_, _00548_);
  nor _58041_ (_06369_, _06368_, _06367_);
  nor _58042_ (_06370_, _06222_, _00343_);
  nor _58043_ (_06371_, _06233_, _00302_);
  nor _58044_ (_06372_, _06371_, _06370_);
  and _58045_ (_06373_, _06372_, _06369_);
  nor _58046_ (_06374_, _06226_, _00507_);
  nor _58047_ (_06375_, _06220_, _00466_);
  nor _58048_ (_06376_, _06375_, _06374_);
  nor _58049_ (_06377_, _06231_, _00731_);
  nor _58050_ (_06378_, _06207_, _00649_);
  nor _58051_ (_06379_, _06378_, _06377_);
  and _58052_ (_06380_, _06379_, _06376_);
  and _58053_ (_06381_, _06380_, _06373_);
  nor _58054_ (_06382_, _06189_, _00066_);
  nor _58055_ (_06383_, _06217_, _00162_);
  nor _58056_ (_06384_, _06383_, _06382_);
  nor _58057_ (_06385_, _06182_, _00384_);
  nor _58058_ (_06386_, _06228_, _00261_);
  nor _58059_ (_06387_, _06386_, _06385_);
  and _58060_ (_06388_, _06387_, _06384_);
  nor _58061_ (_06389_, _06215_, _00690_);
  nor _58062_ (_06390_, _06194_, _00425_);
  nor _58063_ (_06391_, _06390_, _06389_);
  nor _58064_ (_06392_, _06196_, _00220_);
  nor _58065_ (_06393_, _06203_, _00107_);
  nor _58066_ (_06394_, _06393_, _06392_);
  and _58067_ (_06395_, _06394_, _06391_);
  and _58068_ (_06396_, _06395_, _06388_);
  and _58069_ (_06397_, _06396_, _06381_);
  and _58070_ (_06398_, _06397_, _06366_);
  nor _58071_ (_06399_, _06398_, _06365_);
  and _58072_ (_06400_, _06338_, _06276_);
  and _58073_ (_06401_, _06338_, _06002_);
  nor _58074_ (_06402_, _06401_, _06400_);
  nor _58075_ (_06403_, _06402_, _06399_);
  and _58076_ (_06404_, _06344_, _05988_);
  nor _58077_ (_06405_, _06404_, _06345_);
  not _58078_ (_06406_, _06405_);
  and _58079_ (_06407_, _06406_, _06399_);
  nor _58080_ (_06408_, _06357_, _06399_);
  not _58081_ (_06409_, \oc8051_golden_model_1.SP [3]);
  and _58082_ (_06410_, _06355_, _05988_);
  and _58083_ (_06411_, _06410_, _06409_);
  not _58084_ (_06412_, _06036_);
  and _58085_ (_06413_, _06061_, _06051_);
  nor _58086_ (_06414_, _06413_, _06412_);
  not _58087_ (_06415_, _06414_);
  or _58088_ (_06416_, _06415_, _06269_);
  and _58089_ (_06417_, _06350_, _06036_);
  nor _58090_ (_06418_, _06410_, _06356_);
  not _58091_ (_06419_, \oc8051_golden_model_1.PSW [3]);
  or _58092_ (_06420_, _06414_, _06419_);
  and _58093_ (_06421_, _06420_, _06418_);
  or _58094_ (_06422_, _06421_, _06417_);
  and _58095_ (_06423_, _06422_, _06416_);
  or _58096_ (_06424_, _06423_, _06411_);
  nor _58097_ (_06425_, _06424_, _06408_);
  not _58098_ (_06426_, _06417_);
  nor _58099_ (_06427_, _06426_, _06269_);
  nor _58100_ (_06428_, _06427_, _06425_);
  nor _58101_ (_06429_, _06428_, _06352_);
  and _58102_ (_06430_, _06399_, _06352_);
  and _58103_ (_06431_, _06344_, _06036_);
  nor _58104_ (_06432_, _06431_, _06351_);
  not _58105_ (_06433_, _06432_);
  nor _58106_ (_06434_, _06433_, _06430_);
  not _58107_ (_06435_, _06434_);
  nor _58108_ (_06436_, _06435_, _06429_);
  and _58109_ (_06437_, _06433_, _06269_);
  or _58110_ (_06438_, _06437_, _06406_);
  nor _58111_ (_06439_, _06438_, _06436_);
  nor _58112_ (_06440_, _06439_, _06407_);
  nor _58113_ (_06441_, _06054_, _06034_);
  nor _58114_ (_06442_, _06441_, _06440_);
  not _58115_ (_06443_, _06054_);
  and _58116_ (_06444_, _06443_, _05988_);
  and _58117_ (_06445_, _06338_, _06443_);
  nor _58118_ (_06446_, _06445_, _06444_);
  not _58119_ (_06447_, _06446_);
  not _58120_ (_06448_, _06441_);
  nor _58121_ (_06449_, _06448_, _06269_);
  nor _58122_ (_06450_, _06449_, _06447_);
  not _58123_ (_06451_, _06450_);
  nor _58124_ (_06452_, _06451_, _06442_);
  and _58125_ (_06453_, _06038_, _06036_);
  nor _58126_ (_06454_, _06446_, _06399_);
  nor _58127_ (_06455_, _06454_, _06453_);
  not _58128_ (_06456_, _06455_);
  nor _58129_ (_06457_, _06456_, _06452_);
  not _58130_ (_06458_, _06453_);
  nor _58131_ (_06459_, _06458_, _06269_);
  nor _58132_ (_06460_, _06459_, _06457_);
  or _58133_ (_06461_, _06460_, _06339_);
  nand _58134_ (_06462_, _06399_, _06339_);
  and _58135_ (_06463_, _06462_, _06461_);
  or _58136_ (_06464_, _06463_, _06037_);
  not _58137_ (_06465_, _06402_);
  and _58138_ (_06466_, _06318_, _06033_);
  and _58139_ (_06467_, _06466_, _06344_);
  and _58140_ (_06468_, _06314_, _05923_);
  and _58141_ (_06469_, _06468_, _06344_);
  nor _58142_ (_06470_, _06469_, _06467_);
  and _58143_ (_06471_, _06035_, _05921_);
  and _58144_ (_06472_, _06471_, _06344_);
  not _58145_ (_06473_, _06472_);
  and _58146_ (_06474_, _06355_, _06036_);
  and _58147_ (_06475_, _06318_, _06029_);
  and _58148_ (_06476_, _06475_, _06344_);
  nor _58149_ (_06477_, _06476_, _06474_);
  and _58150_ (_06478_, _06477_, _06473_);
  and _58151_ (_06479_, _06478_, _06470_);
  and _58152_ (_06480_, _06314_, _06033_);
  and _58153_ (_06481_, _06480_, _06344_);
  nor _58154_ (_06482_, _06324_, _06048_);
  or _58155_ (_06483_, _06482_, _06481_);
  not _58156_ (_06484_, _06483_);
  and _58157_ (_06485_, _06484_, _06479_);
  and _58158_ (_06486_, _06038_, _05988_);
  not _58159_ (_06487_, _06486_);
  and _58160_ (_06488_, _06338_, _05996_);
  and _58161_ (_06489_, _06035_, _05923_);
  and _58162_ (_06490_, _06489_, _06344_);
  nor _58163_ (_06491_, _06490_, _06488_);
  and _58164_ (_06492_, _06491_, _06487_);
  and _58165_ (_06493_, _06318_, _06328_);
  and _58166_ (_06494_, _06493_, _06344_);
  not _58167_ (_06495_, _06494_);
  and _58168_ (_06496_, _06360_, _05988_);
  nor _58169_ (_06497_, _06496_, _06277_);
  and _58170_ (_06498_, _06497_, _06495_);
  and _58171_ (_06499_, _06498_, _06492_);
  not _58172_ (_06500_, _06431_);
  not _58173_ (_06501_, _06011_);
  and _58174_ (_06502_, _06030_, _06501_);
  and _58175_ (_06503_, _06338_, _05848_);
  nor _58176_ (_06504_, _06503_, _06502_);
  and _58177_ (_06505_, _06504_, _06500_);
  not _58178_ (_06506_, _06017_);
  and _58179_ (_06507_, _06030_, _06506_);
  not _58180_ (_06508_, _06022_);
  and _58181_ (_06509_, _06030_, _06508_);
  nor _58182_ (_06510_, _06509_, _06507_);
  not _58183_ (_06511_, _06015_);
  and _58184_ (_06512_, _06511_, _05988_);
  nor _58185_ (_06513_, _06512_, _05989_);
  and _58186_ (_06514_, _06513_, _06510_);
  and _58187_ (_06515_, _06514_, _06505_);
  and _58188_ (_06516_, _06515_, _06499_);
  and _58189_ (_06517_, _06516_, _06485_);
  nor _58190_ (_06518_, _06517_, _06113_);
  and _58191_ (_06519_, _06517_, _06127_);
  nor _58192_ (_06520_, _06519_, _06518_);
  not _58193_ (_06521_, _06150_);
  nor _58194_ (_06522_, _06517_, _06521_);
  and _58195_ (_06523_, _06517_, _06173_);
  nor _58196_ (_06524_, _06523_, _06522_);
  nor _58197_ (_06525_, _06524_, _06520_);
  nor _58198_ (_06526_, _06431_, _06512_);
  nor _58199_ (_06527_, _06502_, _05989_);
  and _58200_ (_06528_, _06527_, _06526_);
  nor _58201_ (_06529_, _06503_, \oc8051_golden_model_1.PC [0]);
  and _58202_ (_06530_, _06529_, _06510_);
  and _58203_ (_06531_, _06530_, _06528_);
  and _58204_ (_06532_, _06531_, _06499_);
  and _58205_ (_06533_, _06532_, _06485_);
  nor _58206_ (_06534_, _06533_, _05667_);
  and _58207_ (_06535_, _06533_, _05667_);
  nor _58208_ (_06536_, _06535_, _06534_);
  nor _58209_ (_06537_, _06517_, \oc8051_golden_model_1.PC [0]);
  and _58210_ (_06538_, _06517_, \oc8051_golden_model_1.PC [0]);
  nor _58211_ (_06539_, _06538_, _06537_);
  and _58212_ (_06540_, _06539_, _06536_);
  and _58213_ (_06541_, _06540_, _06525_);
  and _58214_ (_06542_, _06541_, _04760_);
  nor _58215_ (_06543_, _06539_, _06536_);
  not _58216_ (_06544_, _06520_);
  and _58217_ (_06545_, _06524_, _06544_);
  and _58218_ (_06546_, _06545_, _06543_);
  and _58219_ (_06547_, _06546_, _04739_);
  nor _58220_ (_06548_, _06547_, _06542_);
  not _58221_ (_06549_, _06536_);
  nor _58222_ (_06550_, _06539_, _06549_);
  and _58223_ (_06551_, _06550_, _06525_);
  and _58224_ (_06552_, _06551_, _04762_);
  nor _58225_ (_06553_, _06524_, _06544_);
  and _58226_ (_06554_, _06543_, _06553_);
  and _58227_ (_06555_, _06554_, _04768_);
  nor _58228_ (_06556_, _06555_, _06552_);
  and _58229_ (_06557_, _06556_, _06548_);
  and _58230_ (_06558_, _06539_, _06549_);
  and _58231_ (_06559_, _06524_, _06520_);
  and _58232_ (_06560_, _06559_, _06558_);
  and _58233_ (_06561_, _06560_, _04743_);
  and _58234_ (_06562_, _06559_, _06550_);
  and _58235_ (_06563_, _06562_, _04777_);
  nor _58236_ (_06564_, _06563_, _06561_);
  and _58237_ (_06565_, _06553_, _06540_);
  and _58238_ (_06566_, _06565_, _04749_);
  and _58239_ (_06567_, _06559_, _06540_);
  and _58240_ (_06568_, _06567_, _04741_);
  nor _58241_ (_06569_, _06568_, _06566_);
  and _58242_ (_06570_, _06569_, _06564_);
  and _58243_ (_06571_, _06570_, _06557_);
  and _58244_ (_06572_, _06558_, _06525_);
  and _58245_ (_06573_, _06572_, _04752_);
  and _58246_ (_06574_, _06543_, _06525_);
  and _58247_ (_06575_, _06574_, _04747_);
  nor _58248_ (_06576_, _06575_, _06573_);
  and _58249_ (_06577_, _06553_, _06558_);
  and _58250_ (_06578_, _06577_, _04766_);
  and _58251_ (_06579_, _06545_, _06550_);
  and _58252_ (_06580_, _06579_, _04773_);
  nor _58253_ (_06581_, _06580_, _06578_);
  and _58254_ (_06582_, _06581_, _06576_);
  and _58255_ (_06583_, _06553_, _06550_);
  and _58256_ (_06584_, _06583_, _04775_);
  and _58257_ (_06585_, _06545_, _06540_);
  and _58258_ (_06586_, _06585_, _04758_);
  nor _58259_ (_06587_, _06586_, _06584_);
  and _58260_ (_06588_, _06545_, _06558_);
  and _58261_ (_06589_, _06588_, _04754_);
  and _58262_ (_06590_, _06559_, _06543_);
  and _58263_ (_06591_, _06590_, _04771_);
  nor _58264_ (_06592_, _06591_, _06589_);
  and _58265_ (_06593_, _06592_, _06587_);
  and _58266_ (_06594_, _06593_, _06582_);
  and _58267_ (_06595_, _06594_, _06571_);
  nor _58268_ (_06596_, _06595_, _06313_);
  nor _58269_ (_06597_, _06596_, _06465_);
  and _58270_ (_06598_, _06597_, _06464_);
  or _58271_ (_06599_, _06598_, _06403_);
  and _58272_ (_06600_, _06036_, _06511_);
  not _58273_ (_06601_, _06600_);
  and _58274_ (_06602_, _06338_, _06508_);
  nor _58275_ (_06603_, _06602_, _06509_);
  and _58276_ (_06604_, _06036_, _06508_);
  not _58277_ (_06605_, _06604_);
  and _58278_ (_06606_, _06605_, _06603_);
  and _58279_ (_06607_, _06606_, _06601_);
  and _58280_ (_06608_, _06036_, _06506_);
  not _58281_ (_06609_, _06608_);
  and _58282_ (_06610_, _06338_, _06506_);
  nor _58283_ (_06611_, _06610_, _06507_);
  and _58284_ (_06612_, _06611_, _06609_);
  and _58285_ (_06613_, _06036_, _06501_);
  not _58286_ (_06614_, _06613_);
  and _58287_ (_06615_, _06338_, _06501_);
  nor _58288_ (_06616_, _06615_, _06502_);
  and _58289_ (_06617_, _06616_, _06614_);
  and _58290_ (_06618_, _06617_, _06612_);
  and _58291_ (_06619_, _06618_, _06607_);
  nand _58292_ (_06620_, _06619_, _06599_);
  and _58293_ (_06621_, _06338_, _06511_);
  not _58294_ (_06622_, _06269_);
  nor _58295_ (_06623_, _06619_, _06622_);
  nor _58296_ (_06624_, _06623_, _06621_);
  and _58297_ (_06625_, _06624_, _06620_);
  and _58298_ (_06626_, _06621_, \oc8051_golden_model_1.SP [3]);
  or _58299_ (_06627_, _06626_, _06512_);
  nor _58300_ (_06628_, _06627_, _06625_);
  not _58301_ (_06629_, _06512_);
  nor _58302_ (_06630_, _06629_, _06399_);
  or _58303_ (_06631_, _06630_, _06628_);
  and _58304_ (_06632_, _06631_, _06364_);
  and _58305_ (_06633_, _06363_, _06269_);
  or _58306_ (_06634_, _06633_, _06632_);
  nand _58307_ (_06635_, _06634_, _06362_);
  and _58308_ (_06636_, _06361_, _06409_);
  nor _58309_ (_06637_, _06636_, _06496_);
  and _58310_ (_06638_, _06637_, _06635_);
  and _58311_ (_06639_, _06036_, _05848_);
  and _58312_ (_06640_, _06399_, _06496_);
  or _58313_ (_06641_, _06640_, _06639_);
  nor _58314_ (_06642_, _06641_, _06638_);
  and _58315_ (_06643_, _06639_, _06269_);
  or _58316_ (_06644_, _06643_, _06642_);
  nand _58317_ (_06645_, _06644_, _05990_);
  and _58318_ (_06646_, _06036_, _05996_);
  nor _58319_ (_06647_, _06399_, _05990_);
  nor _58320_ (_06649_, _06647_, _06646_);
  nand _58321_ (_06650_, _06649_, _06645_);
  not _58322_ (_06651_, _06646_);
  nor _58323_ (_06652_, _06651_, _06269_);
  not _58324_ (_06653_, _06652_);
  and _58325_ (_06654_, _06653_, _06650_);
  nor _58326_ (_06655_, _06189_, _00061_);
  nor _58327_ (_06656_, _06217_, _00151_);
  nor _58328_ (_06657_, _06656_, _06655_);
  nor _58329_ (_06658_, _06207_, _00644_);
  nor _58330_ (_06659_, _06209_, _00603_);
  nor _58331_ (_06660_, _06659_, _06658_);
  and _58332_ (_06661_, _06660_, _06657_);
  nor _58333_ (_06662_, _06200_, _00543_);
  nor _58334_ (_06663_, _06220_, _00461_);
  nor _58335_ (_06664_, _06663_, _06662_);
  nor _58336_ (_06665_, _06233_, _00297_);
  nor _58337_ (_06666_, _06203_, _00102_);
  nor _58338_ (_06667_, _06666_, _06665_);
  and _58339_ (_06668_, _06667_, _06664_);
  and _58340_ (_06669_, _06668_, _06661_);
  nor _58341_ (_06670_, _06231_, _00726_);
  nor _58342_ (_06671_, _06215_, _00685_);
  nor _58343_ (_06672_, _06671_, _06670_);
  nor _58344_ (_06673_, _06222_, _00338_);
  nor _58345_ (_06674_, _06228_, _00256_);
  nor _58346_ (_06675_, _06674_, _06673_);
  and _58347_ (_06676_, _06675_, _06672_);
  nor _58348_ (_06677_, _06182_, _00379_);
  nor _58349_ (_06678_, _06194_, _00420_);
  nor _58350_ (_06679_, _06678_, _06677_);
  nor _58351_ (_06680_, _06226_, _00502_);
  nor _58352_ (_06681_, _06196_, _00215_);
  nor _58353_ (_06682_, _06681_, _06680_);
  and _58354_ (_06683_, _06682_, _06679_);
  and _58355_ (_06684_, _06683_, _06676_);
  and _58356_ (_06685_, _06684_, _06669_);
  nor _58357_ (_06686_, _06685_, _06238_);
  nor _58358_ (_06687_, _06352_, _06339_);
  nor _58359_ (_06688_, _06356_, _06496_);
  and _58360_ (_06689_, _06688_, _06687_);
  and _58361_ (_06690_, _06405_, _06402_);
  and _58362_ (_06691_, _06513_, _06446_);
  and _58363_ (_06692_, _06691_, _06690_);
  and _58364_ (_06693_, _06692_, _06689_);
  not _58365_ (_06694_, _06693_);
  and _58366_ (_06695_, _06694_, _06686_);
  not _58367_ (_06696_, _06695_);
  nor _58368_ (_06697_, _06189_, _00046_);
  nor _58369_ (_06698_, _06217_, _00128_);
  nor _58370_ (_06699_, _06698_, _06697_);
  nor _58371_ (_06700_, _06215_, _00670_);
  nor _58372_ (_06701_, _06222_, _00323_);
  nor _58373_ (_06702_, _06701_, _06700_);
  and _58374_ (_06703_, _06702_, _06699_);
  nor _58375_ (_06704_, _06200_, _00528_);
  nor _58376_ (_06705_, _06194_, _00405_);
  nor _58377_ (_06706_, _06705_, _06704_);
  nor _58378_ (_06707_, _06228_, _00241_);
  nor _58379_ (_06708_, _06203_, _00087_);
  nor _58380_ (_06709_, _06708_, _06707_);
  and _58381_ (_06710_, _06709_, _06706_);
  and _58382_ (_06711_, _06710_, _06703_);
  nor _58383_ (_06712_, _06209_, _00581_);
  nor _58384_ (_06713_, _06220_, _00446_);
  nor _58385_ (_06714_, _06713_, _06712_);
  nor _58386_ (_06715_, _06231_, _00711_);
  nor _58387_ (_06716_, _06207_, _00629_);
  nor _58388_ (_06717_, _06716_, _06715_);
  and _58389_ (_06718_, _06717_, _06714_);
  nor _58390_ (_06719_, _06226_, _00487_);
  nor _58391_ (_06720_, _06196_, _00200_);
  nor _58392_ (_06721_, _06720_, _06719_);
  nor _58393_ (_06722_, _06182_, _00364_);
  nor _58394_ (_06723_, _06233_, _00282_);
  nor _58395_ (_06724_, _06723_, _06722_);
  and _58396_ (_06725_, _06724_, _06721_);
  and _58397_ (_06726_, _06725_, _06718_);
  and _58398_ (_06727_, _06726_, _06711_);
  nor _58399_ (_06728_, _06417_, _06639_);
  nor _58400_ (_06729_, _06453_, _06441_);
  and _58401_ (_06730_, _06729_, _06728_);
  and _58402_ (_06731_, _06432_, _06415_);
  and _58403_ (_06732_, _06731_, _06730_);
  and _58404_ (_06733_, _06732_, _06618_);
  and _58405_ (_06734_, _06651_, _06607_);
  and _58406_ (_06735_, _06734_, _06364_);
  and _58407_ (_06736_, _06735_, _06733_);
  nor _58408_ (_06737_, _06736_, _06727_);
  not _58409_ (_06738_, _06737_);
  and _58410_ (_06739_, _06572_, _04706_);
  and _58411_ (_06740_, _06585_, _04712_);
  nor _58412_ (_06741_, _06740_, _06739_);
  and _58413_ (_06742_, _06588_, _04708_);
  and _58414_ (_06743_, _06590_, _04733_);
  nor _58415_ (_06744_, _06743_, _06742_);
  and _58416_ (_06745_, _06744_, _06741_);
  and _58417_ (_06746_, _06565_, _04703_);
  and _58418_ (_06747_, _06567_, _04695_);
  nor _58419_ (_06748_, _06747_, _06746_);
  and _58420_ (_06749_, _06583_, _04724_);
  and _58421_ (_06750_, _06554_, _04720_);
  nor _58422_ (_06751_, _06750_, _06749_);
  and _58423_ (_06752_, _06751_, _06748_);
  and _58424_ (_06753_, _06752_, _06745_);
  and _58425_ (_06754_, _06579_, _04722_);
  and _58426_ (_06755_, _06546_, _04693_);
  nor _58427_ (_06756_, _06755_, _06754_);
  and _58428_ (_06757_, _06541_, _04714_);
  and _58429_ (_06758_, _06560_, _04697_);
  nor _58430_ (_06759_, _06758_, _06757_);
  and _58431_ (_06760_, _06759_, _06756_);
  and _58432_ (_06761_, _06551_, _04716_);
  and _58433_ (_06762_, _06562_, _04726_);
  nor _58434_ (_06763_, _06762_, _06761_);
  and _58435_ (_06764_, _06574_, _04701_);
  and _58436_ (_06765_, _06577_, _04731_);
  nor _58437_ (_06766_, _06765_, _06764_);
  and _58438_ (_06767_, _06766_, _06763_);
  and _58439_ (_06768_, _06767_, _06760_);
  and _58440_ (_06769_, _06768_, _06753_);
  nor _58441_ (_06770_, _06769_, _06313_);
  not _58442_ (_06771_, \oc8051_golden_model_1.SP [2]);
  not _58443_ (_06772_, _06410_);
  nor _58444_ (_06773_, _06621_, _06361_);
  and _58445_ (_06774_, _06773_, _06772_);
  nor _58446_ (_06775_, _06774_, _06771_);
  not _58447_ (_06776_, _06775_);
  not _58448_ (_06777_, _06322_);
  not _58449_ (_06778_, _06038_);
  and _58450_ (_06779_, _06061_, _06778_);
  and _58451_ (_06780_, _06048_, _06015_);
  and _58452_ (_06781_, _06780_, _06020_);
  and _58453_ (_06782_, _06781_, _06779_);
  nor _58454_ (_06783_, _06782_, _06777_);
  not _58455_ (_06784_, _06783_);
  and _58456_ (_06785_, _06318_, _05921_);
  nor _58457_ (_06786_, _05808_, _05768_);
  and _58458_ (_06787_, _06786_, _06785_);
  not _58459_ (_06788_, _06787_);
  and _58460_ (_06789_, _06785_, _06508_);
  and _58461_ (_06790_, _06785_, _06002_);
  nor _58462_ (_06791_, _06790_, _06789_);
  and _58463_ (_06792_, _06318_, _05922_);
  not _58464_ (_06793_, _06792_);
  not _58465_ (_06794_, _05996_);
  and _58466_ (_06795_, _06056_, _06794_);
  nor _58467_ (_06796_, _06795_, _06793_);
  not _58468_ (_06797_, _06796_);
  and _58469_ (_06798_, _06797_, _06791_);
  and _58470_ (_06799_, _06798_, _06788_);
  and _58471_ (_06800_, _06799_, _06784_);
  and _58472_ (_06801_, _06800_, _06776_);
  and _58473_ (_06802_, _06322_, _06501_);
  and _58474_ (_06803_, _06466_, _06501_);
  nor _58475_ (_06804_, _06803_, _06802_);
  not _58476_ (_06805_, _06785_);
  and _58477_ (_06806_, _06048_, _06778_);
  and _58478_ (_06807_, _06806_, _06413_);
  nor _58479_ (_06808_, _06807_, _06805_);
  and _58480_ (_06809_, _06017_, _06015_);
  and _58481_ (_06810_, _06056_, _06011_);
  and _58482_ (_06811_, _06810_, _06809_);
  nor _58483_ (_06812_, _06811_, _06805_);
  nor _58484_ (_06813_, _06812_, _06808_);
  and _58485_ (_06814_, _06813_, _06804_);
  not _58486_ (_06815_, _06061_);
  and _58487_ (_06816_, _06466_, _06815_);
  nor _58488_ (_06817_, _06816_, _06467_);
  and _58489_ (_06818_, _06322_, _06002_);
  and _58490_ (_06819_, _06785_, _05848_);
  nor _58491_ (_06820_, _06819_, _06818_);
  and _58492_ (_06821_, _06820_, _06817_);
  or _58493_ (_06822_, _06038_, _06002_);
  nand _58494_ (_06823_, _06015_, _06020_);
  or _58495_ (_06824_, _06823_, _06822_);
  and _58496_ (_06825_, _06824_, _06466_);
  not _58497_ (_06826_, _06825_);
  and _58498_ (_06827_, _06792_, _06508_);
  and _58499_ (_06828_, _06792_, _06506_);
  nor _58500_ (_06829_, _06828_, _06827_);
  and _58501_ (_06830_, _06792_, _06355_);
  and _58502_ (_06831_, _06792_, _05848_);
  nor _58503_ (_06832_, _06831_, _06830_);
  and _58504_ (_06833_, _06832_, _06829_);
  and _58505_ (_06834_, _06833_, _06826_);
  and _58506_ (_06835_, _06834_, _06821_);
  and _58507_ (_06836_, _06835_, _06814_);
  and _58508_ (_06837_, _06836_, _06801_);
  not _58509_ (_06838_, _06837_);
  nor _58510_ (_06839_, _06838_, _06770_);
  and _58511_ (_06840_, _06839_, _06738_);
  and _58512_ (_06841_, _06840_, _06696_);
  nor _58513_ (_06842_, _06651_, _06310_);
  not _58514_ (_06843_, _06842_);
  nor _58515_ (_06844_, _06458_, _06310_);
  nor _58516_ (_06845_, _06446_, _06270_);
  nor _58517_ (_06846_, _06500_, _06310_);
  or _58518_ (_06847_, _06426_, _06310_);
  nor _58519_ (_06848_, _06415_, _06310_);
  nor _58520_ (_06849_, _06322_, _06036_);
  and _58521_ (_06850_, _06314_, _05884_);
  nor _58522_ (_06851_, _06850_, _06329_);
  and _58523_ (_06852_, _06851_, _06849_);
  nor _58524_ (_06853_, _06852_, _06061_);
  not _58525_ (_06854_, _06853_);
  and _58526_ (_06855_, _06493_, _06815_);
  not _58527_ (_06856_, _06059_);
  and _58528_ (_06857_, _06329_, _06856_);
  nor _58529_ (_06858_, _06857_, _06855_);
  not _58530_ (_06859_, _06329_);
  and _58531_ (_06860_, _06849_, _06859_);
  nor _58532_ (_06861_, _06860_, _06051_);
  not _58533_ (_06862_, _06861_);
  and _58534_ (_06863_, _06850_, _06355_);
  and _58535_ (_06864_, _06318_, _05884_);
  and _58536_ (_06865_, _06864_, _06355_);
  and _58537_ (_06866_, _06865_, _05921_);
  nor _58538_ (_06867_, _06866_, _06863_);
  and _58539_ (_06868_, _06867_, _06862_);
  and _58540_ (_06869_, _06868_, _06858_);
  and _58541_ (_06870_, _06869_, _06854_);
  or _58542_ (_06871_, _06870_, _06848_);
  nand _58543_ (_06872_, _06871_, _06357_);
  nand _58544_ (_06873_, _06358_, _06872_);
  and _58545_ (_06874_, _06410_, _06342_);
  nor _58546_ (_06875_, _06874_, _06417_);
  and _58547_ (_06876_, _05985_, _05884_);
  nor _58548_ (_06877_, _06329_, _06876_);
  nor _58549_ (_06878_, _06877_, _06056_);
  not _58550_ (_06879_, _06878_);
  and _58551_ (_06880_, _06879_, _06875_);
  nand _58552_ (_06881_, _06880_, _06873_);
  nand _58553_ (_06882_, _06881_, _06847_);
  and _58554_ (_06883_, _06882_, _06353_);
  or _58555_ (_06884_, _06354_, _06883_);
  and _58556_ (_06885_, _06351_, _06310_);
  nor _58557_ (_06886_, _06864_, _06036_);
  and _58558_ (_06887_, _06886_, _06851_);
  nor _58559_ (_06888_, _06887_, _06048_);
  nor _58560_ (_06889_, _06888_, _06885_);
  and _58561_ (_06890_, _06889_, _06884_);
  or _58562_ (_06891_, _06890_, _06846_);
  nand _58563_ (_06892_, _06891_, _06405_);
  nor _58564_ (_06893_, _06405_, _06270_);
  nor _58565_ (_06894_, _06893_, _06441_);
  nand _58566_ (_06895_, _06894_, _06892_);
  and _58567_ (_06896_, _06441_, _06310_);
  and _58568_ (_06897_, _06329_, _06443_);
  nor _58569_ (_06898_, _06897_, _06447_);
  not _58570_ (_06899_, _06898_);
  nor _58571_ (_06900_, _06899_, _06896_);
  and _58572_ (_06901_, _06900_, _06895_);
  or _58573_ (_06902_, _06901_, _06845_);
  and _58574_ (_06903_, _06314_, _06328_);
  or _58575_ (_06904_, _06493_, _06903_);
  and _58576_ (_06905_, _06904_, _06038_);
  not _58577_ (_06906_, _06905_);
  and _58578_ (_06907_, _06322_, _06038_);
  nor _58579_ (_06908_, _06907_, _06453_);
  and _58580_ (_06909_, _06329_, _06038_);
  and _58581_ (_06910_, _06468_, _06038_);
  nor _58582_ (_06911_, _06910_, _06909_);
  and _58583_ (_06912_, _06911_, _06908_);
  and _58584_ (_06913_, _06912_, _06906_);
  and _58585_ (_06914_, _06913_, _06902_);
  or _58586_ (_06915_, _06914_, _06844_);
  and _58587_ (_06916_, _06915_, _06340_);
  nor _58588_ (_06917_, _06916_, _06341_);
  nor _58589_ (_06918_, _06887_, _06003_);
  nor _58590_ (_06919_, _06918_, _06917_);
  and _58591_ (_06920_, _06541_, _04621_);
  and _58592_ (_06921_, _06590_, _04641_);
  nor _58593_ (_06922_, _06921_, _06920_);
  and _58594_ (_06923_, _06565_, _04610_);
  and _58595_ (_06924_, _06567_, _04602_);
  nor _58596_ (_06925_, _06924_, _06923_);
  and _58597_ (_06926_, _06925_, _06922_);
  and _58598_ (_06927_, _06577_, _04639_);
  and _58599_ (_06928_, _06562_, _04633_);
  nor _58600_ (_06929_, _06928_, _06927_);
  and _58601_ (_06930_, _06579_, _04629_);
  and _58602_ (_06931_, _06546_, _04600_);
  nor _58603_ (_06932_, _06931_, _06930_);
  and _58604_ (_06933_, _06932_, _06929_);
  and _58605_ (_06934_, _06933_, _06926_);
  and _58606_ (_06935_, _06588_, _04615_);
  and _58607_ (_06936_, _06560_, _04604_);
  nor _58608_ (_06937_, _06936_, _06935_);
  and _58609_ (_06938_, _06551_, _04623_);
  and _58610_ (_06939_, _06583_, _04631_);
  nor _58611_ (_06940_, _06939_, _06938_);
  and _58612_ (_06941_, _06940_, _06937_);
  and _58613_ (_06942_, _06574_, _04608_);
  and _58614_ (_06943_, _06554_, _04627_);
  nor _58615_ (_06944_, _06943_, _06942_);
  and _58616_ (_06945_, _06572_, _04613_);
  and _58617_ (_06946_, _06585_, _04619_);
  nor _58618_ (_06947_, _06946_, _06945_);
  and _58619_ (_06948_, _06947_, _06944_);
  and _58620_ (_06949_, _06948_, _06941_);
  and _58621_ (_06950_, _06949_, _06934_);
  nor _58622_ (_06951_, _06950_, _06313_);
  or _58623_ (_06952_, _06951_, _06919_);
  and _58624_ (_06953_, _06401_, _06270_);
  and _58625_ (_06954_, _06329_, _06276_);
  or _58626_ (_06955_, _06954_, _06400_);
  nor _58627_ (_06956_, _06955_, _06953_);
  and _58628_ (_06957_, _06956_, _06952_);
  not _58629_ (_06958_, _06400_);
  nor _58630_ (_06959_, _06958_, _06270_);
  or _58631_ (_06960_, _06959_, _06957_);
  nor _58632_ (_06961_, _06329_, _06903_);
  nor _58633_ (_06962_, _06961_, _06011_);
  not _58634_ (_06963_, _06962_);
  and _58635_ (_06964_, _06493_, _06501_);
  not _58636_ (_06965_, _06964_);
  and _58637_ (_06966_, _06468_, _06501_);
  nor _58638_ (_06967_, _06966_, _06802_);
  and _58639_ (_06968_, _06967_, _06965_);
  and _58640_ (_06969_, _06968_, _06963_);
  and _58641_ (_06970_, _06969_, _06960_);
  nor _58642_ (_06971_, _06617_, _06311_);
  and _58643_ (_06972_, _06468_, _06506_);
  not _58644_ (_06973_, _06972_);
  nor _58645_ (_06974_, _06864_, _06903_);
  nor _58646_ (_06975_, _06974_, _06017_);
  and _58647_ (_06976_, _06471_, _06506_);
  and _58648_ (_06977_, _06976_, _05884_);
  nor _58649_ (_06978_, _06977_, _06975_);
  and _58650_ (_06979_, _06978_, _06973_);
  not _58651_ (_06980_, _06979_);
  nor _58652_ (_06981_, _06980_, _06971_);
  and _58653_ (_06982_, _06981_, _06970_);
  nor _58654_ (_06983_, _06612_, _06311_);
  and _58655_ (_06984_, _06468_, _06508_);
  not _58656_ (_06985_, _06984_);
  nor _58657_ (_06986_, _06974_, _06022_);
  and _58658_ (_06987_, _06471_, _06508_);
  and _58659_ (_06988_, _06987_, _05884_);
  nor _58660_ (_06989_, _06988_, _06986_);
  and _58661_ (_06990_, _06989_, _06985_);
  not _58662_ (_06991_, _06990_);
  nor _58663_ (_06992_, _06991_, _06983_);
  and _58664_ (_06993_, _06992_, _06982_);
  nor _58665_ (_06994_, _06606_, _06311_);
  and _58666_ (_06995_, _06322_, _06511_);
  not _58667_ (_06996_, _06995_);
  and _58668_ (_06997_, _06903_, _06511_);
  nor _58669_ (_06998_, _06997_, _06600_);
  and _58670_ (_06999_, _06998_, _06996_);
  and _58671_ (_07000_, _06493_, _06511_);
  not _58672_ (_07001_, _07000_);
  and _58673_ (_07002_, _06329_, _06511_);
  and _58674_ (_07003_, _06468_, _06511_);
  nor _58675_ (_07004_, _07003_, _07002_);
  and _58676_ (_07005_, _07004_, _07001_);
  and _58677_ (_07006_, _07005_, _06999_);
  not _58678_ (_07007_, _07006_);
  nor _58679_ (_07008_, _07007_, _06994_);
  and _58680_ (_07009_, _07008_, _06993_);
  nor _58681_ (_07010_, _06601_, _06310_);
  or _58682_ (_07011_, _07010_, _07009_);
  and _58683_ (_07012_, _06621_, _06342_);
  nor _58684_ (_07013_, _07012_, _06512_);
  and _58685_ (_07014_, _07013_, _07011_);
  nor _58686_ (_07015_, _06629_, _06270_);
  or _58687_ (_07016_, _07015_, _07014_);
  and _58688_ (_07017_, _06468_, _06360_);
  not _58689_ (_07018_, _07017_);
  and _58690_ (_07019_, _06329_, _06360_);
  not _58691_ (_07020_, _07019_);
  and _58692_ (_07021_, _06322_, _06360_);
  nor _58693_ (_07022_, _07021_, _06363_);
  and _58694_ (_07023_, _06493_, _06360_);
  and _58695_ (_07024_, _06903_, _06360_);
  nor _58696_ (_07025_, _07024_, _07023_);
  and _58697_ (_07026_, _07025_, _07022_);
  and _58698_ (_07027_, _07026_, _07020_);
  and _58699_ (_07028_, _07027_, _07018_);
  and _58700_ (_07029_, _07028_, _07016_);
  nor _58701_ (_07030_, _06364_, _06310_);
  or _58702_ (_07031_, _07030_, _07029_);
  and _58703_ (_07032_, _06361_, _06342_);
  nor _58704_ (_07033_, _07032_, _06496_);
  and _58705_ (_07034_, _07033_, _07031_);
  not _58706_ (_07035_, _06496_);
  nor _58707_ (_07036_, _07035_, _06270_);
  or _58708_ (_07037_, _07036_, _07034_);
  not _58709_ (_07038_, _05848_);
  nor _58710_ (_07039_, _06851_, _07038_);
  not _58711_ (_07040_, _07039_);
  and _58712_ (_07041_, _06493_, _05848_);
  not _58713_ (_07042_, _07041_);
  and _58714_ (_07043_, _06322_, _05848_);
  nor _58715_ (_07044_, _07043_, _06639_);
  and _58716_ (_07045_, _07044_, _07042_);
  and _58717_ (_07046_, _07045_, _07040_);
  and _58718_ (_07047_, _07046_, _07037_);
  not _58719_ (_07048_, _06639_);
  nor _58720_ (_07049_, _07048_, _06310_);
  or _58721_ (_07050_, _07049_, _07047_);
  and _58722_ (_07051_, _07050_, _05990_);
  or _58723_ (_07052_, _07051_, _06271_);
  nor _58724_ (_07053_, _06886_, _06794_);
  not _58725_ (_07054_, _07053_);
  and _58726_ (_07055_, _06471_, _05996_);
  and _58727_ (_07056_, _07055_, _05884_);
  and _58728_ (_07057_, _06850_, _05996_);
  nor _58729_ (_07058_, _07057_, _07056_);
  and _58730_ (_07059_, _07058_, _07054_);
  nand _58731_ (_07060_, _07059_, _07052_);
  and _58732_ (_07061_, _07060_, _06843_);
  nand _58733_ (_07062_, _07061_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _58734_ (_07063_, _06200_, _00538_);
  nor _58735_ (_07064_, _06182_, _00374_);
  nor _58736_ (_07065_, _07064_, _07063_);
  nor _58737_ (_07066_, _06222_, _00333_);
  nor _58738_ (_07067_, _06203_, _00097_);
  nor _58739_ (_07068_, _07067_, _07066_);
  and _58740_ (_07069_, _07068_, _07065_);
  nor _58741_ (_07070_, _06231_, _00721_);
  nor _58742_ (_07071_, _06196_, _00210_);
  nor _58743_ (_07072_, _07071_, _07070_);
  nor _58744_ (_07073_, _06215_, _00680_);
  nor _58745_ (_07074_, _06220_, _00456_);
  nor _58746_ (_07075_, _07074_, _07073_);
  and _58747_ (_07076_, _07075_, _07072_);
  and _58748_ (_07077_, _07076_, _07069_);
  nor _58749_ (_07078_, _06233_, _00292_);
  nor _58750_ (_07079_, _06228_, _00251_);
  nor _58751_ (_07080_, _07079_, _07078_);
  nor _58752_ (_07081_, _06226_, _00497_);
  nor _58753_ (_07082_, _06189_, _00056_);
  nor _58754_ (_07083_, _07082_, _07081_);
  and _58755_ (_07084_, _07083_, _07080_);
  nor _58756_ (_07085_, _06207_, _00639_);
  nor _58757_ (_07086_, _06217_, _00140_);
  nor _58758_ (_07087_, _07086_, _07085_);
  nor _58759_ (_07088_, _06209_, _00597_);
  nor _58760_ (_07089_, _06194_, _00415_);
  nor _58761_ (_07090_, _07089_, _07088_);
  and _58762_ (_07091_, _07090_, _07087_);
  and _58763_ (_07092_, _07091_, _07084_);
  and _58764_ (_07093_, _07092_, _07077_);
  nor _58765_ (_07094_, _07093_, _06238_);
  and _58766_ (_07095_, _07094_, _06694_);
  not _58767_ (_07096_, _07095_);
  nor _58768_ (_07097_, _06200_, _00523_);
  nor _58769_ (_07098_, _06203_, _00082_);
  nor _58770_ (_07099_, _07098_, _07097_);
  nor _58771_ (_07100_, _06231_, _00706_);
  nor _58772_ (_07101_, _06222_, _00318_);
  nor _58773_ (_07102_, _07101_, _07100_);
  and _58774_ (_07103_, _07102_, _07099_);
  nor _58775_ (_07104_, _06226_, _00482_);
  nor _58776_ (_07105_, _06220_, _00441_);
  nor _58777_ (_07106_, _07105_, _07104_);
  nor _58778_ (_07107_, _06215_, _00665_);
  nor _58779_ (_07108_, _06196_, _00195_);
  nor _58780_ (_07109_, _07108_, _07107_);
  and _58781_ (_07110_, _07109_, _07106_);
  and _58782_ (_07111_, _07110_, _07103_);
  nor _58783_ (_07112_, _06228_, _00236_);
  nor _58784_ (_07113_, _06189_, _00041_);
  nor _58785_ (_07114_, _07113_, _07112_);
  nor _58786_ (_07115_, _06182_, _00359_);
  nor _58787_ (_07116_, _06233_, _00277_);
  nor _58788_ (_07117_, _07116_, _07115_);
  and _58789_ (_07118_, _07117_, _07114_);
  nor _58790_ (_07119_, _06194_, _00400_);
  nor _58791_ (_07120_, _06217_, _00123_);
  nor _58792_ (_07121_, _07120_, _07119_);
  nor _58793_ (_07122_, _06207_, _00624_);
  nor _58794_ (_07123_, _06209_, _00573_);
  nor _58795_ (_07124_, _07123_, _07122_);
  and _58796_ (_07125_, _07124_, _07121_);
  and _58797_ (_07126_, _07125_, _07118_);
  and _58798_ (_07127_, _07126_, _07111_);
  nor _58799_ (_07128_, _07127_, _06736_);
  not _58800_ (_07129_, _07128_);
  and _58801_ (_07130_, _06574_, _04657_);
  and _58802_ (_07131_, _06565_, _04660_);
  nor _58803_ (_07132_, _07131_, _07130_);
  and _58804_ (_07133_, _06541_, _04674_);
  and _58805_ (_07134_, _06551_, _04685_);
  nor _58806_ (_07135_, _07134_, _07133_);
  and _58807_ (_07136_, _07135_, _07132_);
  and _58808_ (_07137_, _06585_, _04668_);
  and _58809_ (_07138_, _06579_, _04676_);
  nor _58810_ (_07139_, _07138_, _07137_);
  and _58811_ (_07140_, _06546_, _04647_);
  and _58812_ (_07141_, _06562_, _04680_);
  nor _58813_ (_07142_, _07141_, _07140_);
  and _58814_ (_07143_, _07142_, _07139_);
  and _58815_ (_07144_, _07143_, _07136_);
  and _58816_ (_07145_, _06577_, _04671_);
  and _58817_ (_07146_, _06560_, _04651_);
  nor _58818_ (_07147_, _07146_, _07145_);
  and _58819_ (_07148_, _06554_, _04666_);
  and _58820_ (_07149_, _06567_, _04649_);
  nor _58821_ (_07150_, _07149_, _07148_);
  and _58822_ (_07151_, _07150_, _07147_);
  and _58823_ (_07152_, _06572_, _04655_);
  and _58824_ (_07153_, _06590_, _04687_);
  nor _58825_ (_07154_, _07153_, _07152_);
  and _58826_ (_07155_, _06583_, _04678_);
  and _58827_ (_07156_, _06588_, _04662_);
  nor _58828_ (_07157_, _07156_, _07155_);
  and _58829_ (_07158_, _07157_, _07154_);
  and _58830_ (_07159_, _07158_, _07151_);
  and _58831_ (_07160_, _07159_, _07144_);
  nor _58832_ (_07161_, _07160_, _06313_);
  not _58833_ (_07162_, _06903_);
  and _58834_ (_07163_, _06061_, _06048_);
  and _58835_ (_07164_, _07163_, _06011_);
  nor _58836_ (_07165_, _07164_, _07162_);
  not _58837_ (_07166_, _07165_);
  and _58838_ (_07167_, _06314_, _06029_);
  not _58839_ (_07168_, _07167_);
  and _58840_ (_07169_, _07163_, _06015_);
  nor _58841_ (_07170_, _07169_, _07168_);
  nor _58842_ (_07171_, _07170_, _06808_);
  and _58843_ (_07172_, _07171_, _07166_);
  not _58844_ (_07173_, _06819_);
  and _58845_ (_07174_, _07173_, _06791_);
  and _58846_ (_07175_, _07174_, _06788_);
  not _58847_ (_07176_, _06812_);
  and _58848_ (_07177_, _06323_, _05848_);
  nor _58849_ (_07178_, _07177_, _07024_);
  nor _58850_ (_07179_, _06010_, _05767_);
  and _58851_ (_07180_, _07179_, _07167_);
  nor _58852_ (_07181_, _07180_, _06997_);
  and _58853_ (_07182_, _07181_, _07178_);
  and _58854_ (_07183_, _07182_, _07176_);
  and _58855_ (_07184_, _07183_, _07175_);
  not _58856_ (_07185_, \oc8051_golden_model_1.SP [1]);
  nor _58857_ (_07186_, _06774_, _07185_);
  nand _58858_ (_07187_, _06051_, _06017_);
  or _58859_ (_07188_, _06822_, _06508_);
  nor _58860_ (_07189_, _07188_, _07187_);
  nand _58861_ (_07190_, _07189_, _06795_);
  and _58862_ (_07191_, _07190_, _06323_);
  nor _58863_ (_07192_, _07191_, _07186_);
  and _58864_ (_07193_, _07192_, _07184_);
  and _58865_ (_07194_, _07193_, _07172_);
  not _58866_ (_07195_, _07194_);
  nor _58867_ (_07196_, _07195_, _07161_);
  and _58868_ (_07197_, _07196_, _07129_);
  and _58869_ (_07198_, _07197_, _07096_);
  nand _58870_ (_07199_, _07060_, _06843_);
  nand _58871_ (_07200_, _07199_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _58872_ (_07201_, _07200_, _07198_);
  nand _58873_ (_07202_, _07201_, _07062_);
  nand _58874_ (_07203_, _07199_, \oc8051_golden_model_1.IRAM[3] [0]);
  not _58875_ (_07204_, _07198_);
  nand _58876_ (_07205_, _07061_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _58877_ (_07206_, _07205_, _07204_);
  nand _58878_ (_07207_, _07206_, _07203_);
  nand _58879_ (_07208_, _07207_, _07202_);
  nand _58880_ (_07209_, _07208_, _06841_);
  not _58881_ (_07210_, _06841_);
  not _58882_ (_07211_, \oc8051_golden_model_1.IRAM[7] [0]);
  or _58883_ (_07212_, _07061_, _07211_);
  nand _58884_ (_07213_, _07061_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _58885_ (_07214_, _07213_, _07204_);
  nand _58886_ (_07215_, _07214_, _07212_);
  nand _58887_ (_07216_, _07061_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand _58888_ (_07217_, _07199_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _58889_ (_07218_, _07217_, _07198_);
  nand _58890_ (_07219_, _07218_, _07216_);
  nand _58891_ (_07220_, _07219_, _07215_);
  nand _58892_ (_07221_, _07220_, _07210_);
  nand _58893_ (_07222_, _07221_, _07209_);
  nand _58894_ (_07223_, _07222_, _06654_);
  not _58895_ (_07224_, _06654_);
  nand _58896_ (_07225_, _07199_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _58897_ (_07226_, _07061_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _58898_ (_07227_, _07226_, _07204_);
  nand _58899_ (_07228_, _07227_, _07225_);
  nand _58900_ (_07229_, _07061_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand _58901_ (_07230_, _07199_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _58902_ (_07231_, _07230_, _07198_);
  nand _58903_ (_07232_, _07231_, _07229_);
  nand _58904_ (_07233_, _07232_, _07228_);
  nand _58905_ (_07234_, _07233_, _06841_);
  not _58906_ (_07235_, \oc8051_golden_model_1.IRAM[15] [0]);
  or _58907_ (_07236_, _07061_, _07235_);
  not _58908_ (_07237_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _58909_ (_07238_, _07199_, _07237_);
  and _58910_ (_07239_, _07238_, _07204_);
  nand _58911_ (_07240_, _07239_, _07236_);
  nand _58912_ (_07241_, _07061_, \oc8051_golden_model_1.IRAM[12] [0]);
  not _58913_ (_07242_, \oc8051_golden_model_1.IRAM[13] [0]);
  or _58914_ (_07243_, _07061_, _07242_);
  and _58915_ (_07244_, _07243_, _07198_);
  nand _58916_ (_07245_, _07244_, _07241_);
  nand _58917_ (_07246_, _07245_, _07240_);
  nand _58918_ (_07247_, _07246_, _07210_);
  nand _58919_ (_07248_, _07247_, _07234_);
  nand _58920_ (_07249_, _07248_, _07224_);
  and _58921_ (_07250_, _07249_, _07223_);
  and _58922_ (_07251_, _07250_, _06359_);
  nor _58923_ (_07252_, _06471_, _06315_);
  nor _58924_ (_07253_, _07252_, _06028_);
  or _58925_ (_07254_, _06489_, _05993_);
  or _58926_ (_07255_, _07254_, _07253_);
  and _58927_ (_07256_, _07255_, _06856_);
  not _58928_ (_07257_, _07256_);
  nor _58929_ (_07258_, _07257_, _07251_);
  and _58930_ (_07259_, _06475_, _06815_);
  not _58931_ (_07260_, _07259_);
  nor _58932_ (_07261_, _07260_, _06238_);
  and _58933_ (_07262_, _07261_, _06310_);
  nor _58934_ (_07263_, _07262_, _07258_);
  and _58935_ (_07264_, _06816_, \oc8051_golden_model_1.SP [0]);
  not _58936_ (_07265_, _07264_);
  nor _58937_ (_07266_, _06865_, _06863_);
  and _58938_ (_07267_, _07266_, _07265_);
  and _58939_ (_07268_, _07267_, _07263_);
  and _58940_ (_07269_, _06471_, _06355_);
  not _58941_ (_07270_, _07269_);
  nor _58942_ (_07271_, _07270_, _07250_);
  not _58943_ (_07272_, _07271_);
  and _58944_ (_07273_, _07272_, _07268_);
  nor _58945_ (_07274_, _06357_, _06238_);
  not _58946_ (_07275_, _06474_);
  nor _58947_ (_07276_, _07275_, _06238_);
  and _58948_ (_07277_, _07276_, _06310_);
  nor _58949_ (_07278_, _07277_, _07274_);
  and _58950_ (_07279_, _07278_, _07273_);
  not _58951_ (_07280_, _07279_);
  and _58952_ (_07281_, _07280_, _06358_);
  nor _58953_ (_07282_, _06052_, _06342_);
  nor _58954_ (_07283_, _07282_, _07281_);
  nor _58955_ (_07284_, _06772_, _06238_);
  and _58956_ (_07285_, _07284_, _06310_);
  and _58957_ (_07286_, _06876_, _06350_);
  nor _58958_ (_07287_, _07286_, _07285_);
  and _58959_ (_07288_, _07287_, _07283_);
  and _58960_ (_07289_, _06471_, _06350_);
  not _58961_ (_07290_, _07289_);
  nor _58962_ (_07291_, _07290_, _07250_);
  not _58963_ (_07292_, _07291_);
  and _58964_ (_07293_, _07292_, _07288_);
  nor _58965_ (_07294_, _06353_, _06238_);
  nor _58966_ (_07295_, _06426_, _06238_);
  and _58967_ (_07296_, _07295_, _06310_);
  nor _58968_ (_07297_, _07296_, _07294_);
  and _58969_ (_07298_, _07297_, _07293_);
  nor _58970_ (_07299_, _07298_, _06354_);
  or _58971_ (_07300_, _07299_, _06351_);
  nand _58972_ (_07301_, _06351_, _06342_);
  nand _58973_ (_07302_, _07301_, _07300_);
  and _58974_ (_07303_, _07302_, _06349_);
  nor _58975_ (_07304_, _07303_, _06347_);
  and _58976_ (_07305_, _06441_, _05884_);
  or _58977_ (_07306_, _07305_, _07304_);
  nor _58978_ (_07307_, _07306_, _06343_);
  nor _58979_ (_07308_, _06340_, _06238_);
  and _58980_ (_07309_, _06471_, _06443_);
  not _58981_ (_07310_, _07309_);
  nor _58982_ (_07311_, _07310_, _07250_);
  nor _58983_ (_07312_, _07311_, _07308_);
  and _58984_ (_07313_, _07312_, _07307_);
  nor _58985_ (_07314_, _07313_, _06341_);
  nor _58986_ (_07315_, _07314_, _06039_);
  and _58987_ (_07316_, _06039_, _06342_);
  nor _58988_ (_07317_, _07316_, _07315_);
  and _58989_ (_07318_, _06876_, _06276_);
  or _58990_ (_07319_, _07318_, _07317_);
  nor _58991_ (_07320_, _07319_, _06337_);
  not _58992_ (_07321_, _07250_);
  and _58993_ (_07322_, _06471_, _06276_);
  and _58994_ (_07323_, _07322_, _07321_);
  nor _58995_ (_07324_, _07323_, _06279_);
  and _58996_ (_07325_, _07324_, _07320_);
  nor _58997_ (_07326_, _07325_, _06312_);
  nor _58998_ (_07327_, _07326_, _06275_);
  nor _58999_ (_07328_, _06009_, \oc8051_golden_model_1.SP [0]);
  nor _59000_ (_07329_, _07328_, _07327_);
  not _59001_ (_07330_, _06018_);
  not _59002_ (_07331_, _06610_);
  nor _59003_ (_07332_, _07331_, _06238_);
  not _59004_ (_07333_, _07332_);
  not _59005_ (_07334_, _06502_);
  nor _59006_ (_07335_, _07334_, _06238_);
  not _59007_ (_07336_, _07335_);
  not _59008_ (_07337_, _06615_);
  nor _59009_ (_07338_, _07337_, _06238_);
  not _59010_ (_07339_, _06507_);
  nor _59011_ (_07340_, _07339_, _06238_);
  nor _59012_ (_07341_, _07340_, _07338_);
  and _59013_ (_07342_, _07341_, _07336_);
  and _59014_ (_07343_, _07342_, _07333_);
  nor _59015_ (_07344_, _07343_, _06311_);
  nor _59016_ (_07345_, _07344_, _07330_);
  not _59017_ (_07346_, _07345_);
  nor _59018_ (_07347_, _07346_, _07329_);
  nor _59019_ (_07348_, _06018_, \oc8051_golden_model_1.SP [0]);
  nor _59020_ (_07349_, _07348_, _07347_);
  not _59021_ (_07350_, _06016_);
  nor _59022_ (_07351_, _06603_, _06238_);
  and _59023_ (_07352_, _07351_, _06310_);
  nor _59024_ (_07353_, _07352_, _07350_);
  not _59025_ (_07354_, _07353_);
  nor _59026_ (_07355_, _07354_, _07349_);
  nor _59027_ (_07356_, _07355_, _06274_);
  and _59028_ (_07357_, _06876_, _05848_);
  nor _59029_ (_07358_, _07357_, _07356_);
  nor _59030_ (_07359_, _07048_, _06238_);
  and _59031_ (_07360_, _06471_, _05848_);
  not _59032_ (_07361_, _07360_);
  nor _59033_ (_07362_, _07361_, _07250_);
  nor _59034_ (_07363_, _07362_, _07359_);
  and _59035_ (_07364_, _07363_, _07358_);
  and _59036_ (_07365_, _07359_, _06311_);
  nor _59037_ (_07366_, _07365_, _07364_);
  nor _59038_ (_07367_, _06503_, _05998_);
  nor _59039_ (_07368_, _07367_, _06342_);
  nor _59040_ (_07369_, _07368_, _07366_);
  and _59041_ (_07370_, _07369_, _06273_);
  nor _59042_ (_07371_, _07370_, _06271_);
  and _59043_ (_07372_, _06864_, _05996_);
  or _59044_ (_07373_, _07372_, _07057_);
  nor _59045_ (_07374_, _07373_, _07371_);
  not _59046_ (_07375_, _07055_);
  nor _59047_ (_07376_, _07250_, _07375_);
  not _59048_ (_07377_, _07376_);
  and _59049_ (_07378_, _07377_, _07374_);
  nor _59050_ (_07379_, _06651_, _06238_);
  and _59051_ (_07380_, _07379_, _06310_);
  not _59052_ (_07381_, _07380_);
  and _59053_ (_07382_, _07381_, _07378_);
  not _59054_ (_07383_, _07127_);
  and _59055_ (_07384_, _07379_, _07383_);
  and _59056_ (_07385_, _07094_, _05989_);
  and _59057_ (_07386_, _07185_, \oc8051_golden_model_1.SP [0]);
  and _59058_ (_07387_, \oc8051_golden_model_1.SP [1], _06342_);
  nor _59059_ (_07388_, _07387_, _07386_);
  nor _59060_ (_07389_, _07388_, _06016_);
  and _59061_ (_07390_, _07383_, _06279_);
  and _59062_ (_07391_, _07094_, _06339_);
  not _59063_ (_07392_, _07388_);
  and _59064_ (_07393_, _07392_, _06351_);
  not _59065_ (_07394_, _06351_);
  and _59066_ (_07395_, _06471_, _06856_);
  nand _59067_ (_07396_, _07061_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand _59068_ (_07397_, _07199_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _59069_ (_07398_, _07397_, _07198_);
  nand _59070_ (_07399_, _07398_, _07396_);
  not _59071_ (_07400_, \oc8051_golden_model_1.IRAM[3] [1]);
  or _59072_ (_07401_, _07061_, _07400_);
  not _59073_ (_07402_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _59074_ (_07403_, _07199_, _07402_);
  and _59075_ (_07404_, _07403_, _07204_);
  nand _59076_ (_07405_, _07404_, _07401_);
  nand _59077_ (_07406_, _07405_, _07399_);
  nand _59078_ (_07407_, _07406_, _06841_);
  not _59079_ (_07408_, \oc8051_golden_model_1.IRAM[7] [1]);
  or _59080_ (_07409_, _07061_, _07408_);
  not _59081_ (_07410_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _59082_ (_07411_, _07199_, _07410_);
  and _59083_ (_07412_, _07411_, _07204_);
  nand _59084_ (_07413_, _07412_, _07409_);
  nand _59085_ (_07414_, _07061_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand _59086_ (_07415_, _07199_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _59087_ (_07416_, _07415_, _07198_);
  nand _59088_ (_07417_, _07416_, _07414_);
  nand _59089_ (_07418_, _07417_, _07413_);
  nand _59090_ (_07419_, _07418_, _07210_);
  nand _59091_ (_07420_, _07419_, _07407_);
  nand _59092_ (_07421_, _07420_, _06654_);
  not _59093_ (_07422_, \oc8051_golden_model_1.IRAM[11] [1]);
  or _59094_ (_07423_, _07061_, _07422_);
  not _59095_ (_07424_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _59096_ (_07425_, _07199_, _07424_);
  and _59097_ (_07426_, _07425_, _07204_);
  nand _59098_ (_07427_, _07426_, _07423_);
  nand _59099_ (_07428_, _07061_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand _59100_ (_07429_, _07199_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _59101_ (_07430_, _07429_, _07198_);
  nand _59102_ (_07431_, _07430_, _07428_);
  nand _59103_ (_07432_, _07431_, _07427_);
  nand _59104_ (_07433_, _07432_, _06841_);
  not _59105_ (_07434_, \oc8051_golden_model_1.IRAM[15] [1]);
  or _59106_ (_07435_, _07061_, _07434_);
  not _59107_ (_07436_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _59108_ (_07437_, _07199_, _07436_);
  and _59109_ (_07438_, _07437_, _07204_);
  nand _59110_ (_07439_, _07438_, _07435_);
  nand _59111_ (_07440_, _07061_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand _59112_ (_07441_, _07199_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _59113_ (_07442_, _07441_, _07198_);
  nand _59114_ (_07443_, _07442_, _07440_);
  nand _59115_ (_07444_, _07443_, _07439_);
  nand _59116_ (_07445_, _07444_, _07210_);
  nand _59117_ (_07446_, _07445_, _07433_);
  nand _59118_ (_07447_, _07446_, _07224_);
  nand _59119_ (_07448_, _07447_, _07421_);
  and _59120_ (_07449_, _07448_, _06359_);
  or _59121_ (_07450_, _07449_, _07395_);
  and _59122_ (_07451_, _07261_, _07127_);
  or _59123_ (_07452_, _07451_, _07450_);
  and _59124_ (_07453_, _07388_, _06816_);
  not _59125_ (_07454_, _07453_);
  and _59126_ (_07455_, _06315_, _06355_);
  nor _59127_ (_07456_, _07455_, _06830_);
  and _59128_ (_07457_, _07456_, _07454_);
  not _59129_ (_07458_, _07457_);
  nor _59130_ (_07459_, _07458_, _07452_);
  and _59131_ (_07460_, _07448_, _07269_);
  nor _59132_ (_07461_, _07460_, _07276_);
  and _59133_ (_07462_, _07461_, _07459_);
  and _59134_ (_07463_, _07276_, _07383_);
  nor _59135_ (_07464_, _07463_, _07462_);
  and _59136_ (_07465_, _07093_, _07274_);
  nor _59137_ (_07466_, _07465_, _07464_);
  nor _59138_ (_07467_, _07392_, _06052_);
  nor _59139_ (_07468_, _07467_, _07284_);
  and _59140_ (_07469_, _07468_, _07466_);
  and _59141_ (_07470_, _07284_, _07383_);
  nor _59142_ (_07471_, _07470_, _07469_);
  and _59143_ (_07472_, _05985_, _05922_);
  and _59144_ (_07473_, _07472_, _06350_);
  nor _59145_ (_07474_, _07473_, _07471_);
  and _59146_ (_07475_, _07448_, _07289_);
  nor _59147_ (_07476_, _07475_, _07295_);
  and _59148_ (_07477_, _07476_, _07474_);
  and _59149_ (_07478_, _07295_, _07383_);
  nor _59150_ (_07479_, _07478_, _07477_);
  and _59151_ (_07480_, _07093_, _07294_);
  nor _59152_ (_07481_, _07480_, _07479_);
  and _59153_ (_07482_, _07481_, _07394_);
  nor _59154_ (_07483_, _07482_, _07393_);
  and _59155_ (_07484_, _06348_, _07093_);
  or _59156_ (_07485_, _07484_, _07483_);
  nor _59157_ (_07486_, _07392_, _06049_);
  and _59158_ (_07487_, _07472_, _06443_);
  nor _59159_ (_07488_, _07487_, _07486_);
  not _59160_ (_07489_, _07488_);
  nor _59161_ (_07490_, _07489_, _07485_);
  and _59162_ (_07491_, _07448_, _07309_);
  nor _59163_ (_07492_, _07491_, _07308_);
  and _59164_ (_07493_, _07492_, _07490_);
  nor _59165_ (_07494_, _07493_, _07391_);
  nor _59166_ (_07495_, _07494_, _06039_);
  and _59167_ (_07496_, _07392_, _06039_);
  nor _59168_ (_07497_, _07496_, _07495_);
  nor _59169_ (_07498_, _06336_, _07383_);
  and _59170_ (_07499_, _07472_, _06276_);
  nor _59171_ (_07500_, _07499_, _07498_);
  not _59172_ (_07501_, _07500_);
  nor _59173_ (_07502_, _07501_, _07497_);
  and _59174_ (_07503_, _07448_, _07322_);
  nor _59175_ (_07504_, _07503_, _06279_);
  and _59176_ (_07505_, _07504_, _07502_);
  nor _59177_ (_07506_, _07505_, _07390_);
  nor _59178_ (_07507_, _07506_, _06275_);
  nor _59179_ (_07508_, _07388_, _06009_);
  nor _59180_ (_07509_, _07508_, _07507_);
  nor _59181_ (_07510_, _07343_, _07383_);
  nor _59182_ (_07511_, _07510_, _07330_);
  not _59183_ (_07512_, _07511_);
  nor _59184_ (_07513_, _07512_, _07509_);
  nor _59185_ (_07514_, _07388_, _06018_);
  nor _59186_ (_07515_, _07514_, _07513_);
  and _59187_ (_07516_, _07351_, _07127_);
  nor _59188_ (_07517_, _07516_, _07350_);
  not _59189_ (_07518_, _07517_);
  nor _59190_ (_07519_, _07518_, _07515_);
  nor _59191_ (_07520_, _07519_, _07389_);
  and _59192_ (_07521_, _06315_, _05848_);
  or _59193_ (_07522_, _07521_, _06831_);
  nor _59194_ (_07523_, _07522_, _07520_);
  and _59195_ (_07524_, _07448_, _07360_);
  nor _59196_ (_07525_, _07524_, _07359_);
  and _59197_ (_07526_, _07525_, _07523_);
  and _59198_ (_07527_, _07359_, _07383_);
  nor _59199_ (_07528_, _07527_, _07526_);
  nor _59200_ (_07529_, _07392_, _07367_);
  nor _59201_ (_07530_, _07529_, _06272_);
  not _59202_ (_07531_, _07530_);
  nor _59203_ (_07532_, _07531_, _07528_);
  nor _59204_ (_07533_, _07532_, _07385_);
  and _59205_ (_07534_, _06792_, _05996_);
  and _59206_ (_07535_, _06315_, _05996_);
  nor _59207_ (_07536_, _07535_, _07534_);
  not _59208_ (_07537_, _07536_);
  nor _59209_ (_07538_, _07537_, _07533_);
  and _59210_ (_07539_, _07448_, _07055_);
  nor _59211_ (_07540_, _07539_, _07379_);
  and _59212_ (_07541_, _07540_, _07538_);
  nor _59213_ (_07542_, _07541_, _07384_);
  not _59214_ (_07543_, _00000_);
  or _59215_ (_07544_, _06238_, _06003_);
  nor _59216_ (_07545_, _06322_, _07167_);
  nor _59217_ (_07546_, _06471_, _06903_);
  and _59218_ (_07547_, _07546_, _07545_);
  nor _59219_ (_07548_, _07547_, _07544_);
  not _59220_ (_07549_, _07548_);
  and _59221_ (_07550_, _06056_, _06008_);
  not _59222_ (_07551_, _07550_);
  and _59223_ (_07552_, _07551_, _06468_);
  not _59224_ (_07553_, _07552_);
  and _59225_ (_07554_, _06480_, _06276_);
  nor _59226_ (_07555_, _07554_, _07056_);
  and _59227_ (_07556_, _07555_, _07553_);
  nor _59228_ (_07557_, _06320_, _06008_);
  and _59229_ (_07558_, _07055_, _06028_);
  nor _59230_ (_07559_, _07558_, _07557_);
  nor _59231_ (_07560_, _07252_, _06059_);
  or _59232_ (_07561_, _07521_, _07360_);
  nor _59233_ (_07562_, _07561_, _07560_);
  and _59234_ (_07563_, _07562_, _07559_);
  not _59235_ (_07564_, _06816_);
  nor _59236_ (_07565_, _07322_, _07269_);
  and _59237_ (_07566_, _07565_, _07564_);
  and _59238_ (_07567_, _07367_, _06019_);
  and _59239_ (_07568_, _07567_, _07566_);
  and _59240_ (_07569_, _07568_, _07563_);
  and _59241_ (_07570_, _07569_, _07556_);
  nor _59242_ (_07571_, _06324_, _06008_);
  not _59243_ (_07572_, _07571_);
  and _59244_ (_07573_, _06489_, _06856_);
  and _59245_ (_07574_, _06856_, _06036_);
  nor _59246_ (_07575_, _07574_, _07573_);
  nand _59247_ (_07576_, _07575_, _06060_);
  or _59248_ (_07577_, _06323_, _06318_);
  and _59249_ (_07578_, _07577_, _06443_);
  nor _59250_ (_07579_, _07578_, _07576_);
  and _59251_ (_07580_, _07579_, _07572_);
  and _59252_ (_07581_, _06318_, _05996_);
  nor _59253_ (_07582_, _07289_, _07581_);
  not _59254_ (_07583_, _05923_);
  and _59255_ (_07584_, _06314_, _07583_);
  and _59256_ (_07585_, _07584_, _06350_);
  nor _59257_ (_07586_, _07585_, _07455_);
  and _59258_ (_07587_, _07586_, _07582_);
  and _59259_ (_07588_, _06318_, _05848_);
  nor _59260_ (_07589_, _07588_, _06351_);
  and _59261_ (_07590_, _06323_, _06355_);
  and _59262_ (_07591_, _06314_, _05996_);
  nor _59263_ (_07592_, _07591_, _07590_);
  and _59264_ (_07593_, _07592_, _07589_);
  and _59265_ (_07594_, _07593_, _07587_);
  and _59266_ (_07595_, _06052_, _06009_);
  not _59267_ (_07596_, _06049_);
  nor _59268_ (_07597_, _07596_, _06039_);
  and _59269_ (_07598_, _07597_, _07595_);
  and _59270_ (_07599_, _06056_, _06051_);
  nor _59271_ (_07600_, _07599_, _06319_);
  and _59272_ (_07601_, _06315_, _06443_);
  nor _59273_ (_07602_, _07601_, _07600_);
  nor _59274_ (_07603_, _07309_, _07177_);
  and _59275_ (_07604_, _07603_, _07602_);
  and _59276_ (_07605_, _07604_, _07598_);
  and _59277_ (_07606_, _07605_, _07594_);
  and _59278_ (_07607_, _07606_, _07580_);
  and _59279_ (_07608_, _07607_, _07570_);
  not _59280_ (_07609_, _07608_);
  not _59281_ (_07610_, _06321_);
  nor _59282_ (_07611_, _06316_, _06037_);
  and _59283_ (_07612_, _07611_, _07610_);
  nor _59284_ (_07613_, _07612_, _06238_);
  nor _59285_ (_07614_, _07613_, _07609_);
  nor _59286_ (_07615_, _07261_, _06272_);
  and _59287_ (_07616_, _07615_, _07614_);
  and _59288_ (_07617_, _07616_, _07549_);
  nor _59289_ (_07618_, _07379_, _06279_);
  nor _59290_ (_07619_, _07295_, _07284_);
  and _59291_ (_07620_, _07619_, _07618_);
  nor _59292_ (_07621_, _07359_, _06348_);
  nor _59293_ (_07622_, _07332_, _07276_);
  and _59294_ (_07623_, _07622_, _07621_);
  and _59295_ (_07624_, _07623_, _07620_);
  nor _59296_ (_07625_, _07351_, _07294_);
  nor _59297_ (_07626_, _07308_, _07274_);
  and _59298_ (_07627_, _07626_, _07625_);
  and _59299_ (_07628_, _07627_, _07342_);
  and _59300_ (_07629_, _07628_, _07624_);
  and _59301_ (_07630_, _07629_, _07617_);
  nor _59302_ (_07631_, _07630_, _07543_);
  not _59303_ (_07632_, _07631_);
  nor _59304_ (_07633_, _07632_, _07542_);
  and _59305_ (_07634_, _07633_, _07382_);
  not _59306_ (_07635_, _07634_);
  nand _59307_ (_07636_, _07061_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand _59308_ (_07637_, _07199_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _59309_ (_07638_, _07637_, _07198_);
  nand _59310_ (_07639_, _07638_, _07636_);
  nand _59311_ (_07640_, _07199_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand _59312_ (_07641_, _07061_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _59313_ (_07642_, _07641_, _07204_);
  nand _59314_ (_07643_, _07642_, _07640_);
  nand _59315_ (_07644_, _07643_, _07639_);
  nand _59316_ (_07645_, _07644_, _06841_);
  nand _59317_ (_07646_, _07199_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand _59318_ (_07647_, _07061_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _59319_ (_07648_, _07647_, _07204_);
  nand _59320_ (_07649_, _07648_, _07646_);
  nand _59321_ (_07650_, _07061_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand _59322_ (_07651_, _07199_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _59323_ (_07652_, _07651_, _07198_);
  nand _59324_ (_07653_, _07652_, _07650_);
  nand _59325_ (_07654_, _07653_, _07649_);
  nand _59326_ (_07655_, _07654_, _07210_);
  nand _59327_ (_07656_, _07655_, _07645_);
  nand _59328_ (_07657_, _07656_, _06654_);
  nand _59329_ (_07658_, _07199_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _59330_ (_07659_, _07061_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _59331_ (_07660_, _07659_, _07204_);
  nand _59332_ (_07661_, _07660_, _07658_);
  nand _59333_ (_07662_, _07061_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _59334_ (_07663_, _07199_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _59335_ (_07664_, _07663_, _07198_);
  nand _59336_ (_07665_, _07664_, _07662_);
  nand _59337_ (_07666_, _07665_, _07661_);
  nand _59338_ (_07667_, _07666_, _06841_);
  nand _59339_ (_07668_, _07199_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _59340_ (_07669_, _07061_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _59341_ (_07670_, _07669_, _07204_);
  nand _59342_ (_07671_, _07670_, _07668_);
  nand _59343_ (_07672_, _07061_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _59344_ (_07673_, _07199_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _59345_ (_07674_, _07673_, _07198_);
  nand _59346_ (_07675_, _07674_, _07672_);
  nand _59347_ (_07676_, _07675_, _07671_);
  nand _59348_ (_07677_, _07676_, _07210_);
  nand _59349_ (_07678_, _07677_, _07667_);
  nand _59350_ (_07679_, _07678_, _07224_);
  nand _59351_ (_07680_, _07679_, _07657_);
  and _59352_ (_07681_, _07680_, _07055_);
  and _59353_ (_07682_, _07680_, _07360_);
  and _59354_ (_07683_, _07680_, _07309_);
  and _59355_ (_07684_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _59356_ (_07685_, _07684_, \oc8051_golden_model_1.SP [2]);
  nor _59357_ (_07686_, _07685_, \oc8051_golden_model_1.SP [3]);
  and _59358_ (_07687_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _59359_ (_07688_, _07687_, \oc8051_golden_model_1.SP [3]);
  and _59360_ (_07689_, _07688_, \oc8051_golden_model_1.SP [0]);
  nor _59361_ (_07690_, _07689_, _07686_);
  and _59362_ (_07691_, _07690_, _07596_);
  not _59363_ (_07692_, _06052_);
  and _59364_ (_07693_, _07274_, _06397_);
  and _59365_ (_07694_, _07680_, _07269_);
  and _59366_ (_07695_, _07690_, _06816_);
  and _59367_ (_07696_, _07680_, _06359_);
  and _59368_ (_07697_, _06060_, _06419_);
  nor _59369_ (_07698_, _07697_, _07696_);
  nor _59370_ (_07699_, _07698_, _07261_);
  and _59371_ (_07700_, _07261_, _06269_);
  nor _59372_ (_07701_, _07700_, _06816_);
  not _59373_ (_07702_, _07701_);
  nor _59374_ (_07703_, _07702_, _07699_);
  or _59375_ (_07704_, _07703_, _07269_);
  nor _59376_ (_07705_, _07704_, _07695_);
  or _59377_ (_07706_, _07705_, _07276_);
  nor _59378_ (_07707_, _07706_, _07694_);
  and _59379_ (_07708_, _07276_, _06622_);
  or _59380_ (_07709_, _07708_, _07274_);
  nor _59381_ (_07710_, _07709_, _07707_);
  nor _59382_ (_07711_, _07710_, _07693_);
  nor _59383_ (_07712_, _07711_, _07692_);
  nor _59384_ (_07713_, _07690_, _06052_);
  nor _59385_ (_07714_, _07713_, _07284_);
  not _59386_ (_07715_, _07714_);
  nor _59387_ (_07716_, _07715_, _07712_);
  and _59388_ (_07717_, _07284_, _06622_);
  nor _59389_ (_07718_, _07717_, _07289_);
  not _59390_ (_07719_, _07718_);
  nor _59391_ (_07720_, _07719_, _07716_);
  and _59392_ (_07721_, _07680_, _07289_);
  nor _59393_ (_07722_, _07721_, _07295_);
  not _59394_ (_07723_, _07722_);
  nor _59395_ (_07724_, _07723_, _07720_);
  and _59396_ (_07725_, _07295_, _06622_);
  or _59397_ (_07726_, _07725_, _07294_);
  nor _59398_ (_07727_, _07726_, _07724_);
  and _59399_ (_07728_, _06397_, _07294_);
  nor _59400_ (_07729_, _07728_, _07727_);
  and _59401_ (_07730_, _07729_, _07394_);
  and _59402_ (_07731_, _07690_, _06351_);
  nor _59403_ (_07732_, _07731_, _07730_);
  nor _59404_ (_07733_, _07732_, _06348_);
  and _59405_ (_07734_, _06348_, _06399_);
  or _59406_ (_07735_, _07734_, _07733_);
  and _59407_ (_07736_, _07735_, _06049_);
  or _59408_ (_07737_, _07736_, _07309_);
  nor _59409_ (_07738_, _07737_, _07691_);
  or _59410_ (_07739_, _07738_, _07308_);
  nor _59411_ (_07740_, _07739_, _07683_);
  not _59412_ (_07741_, _06397_);
  and _59413_ (_07742_, _07308_, _07741_);
  or _59414_ (_07743_, _07742_, _06039_);
  or _59415_ (_07744_, _07743_, _07740_);
  not _59416_ (_07745_, _06039_);
  or _59417_ (_07746_, _07690_, _07745_);
  and _59418_ (_07747_, _07746_, _06336_);
  and _59419_ (_07748_, _07747_, _07744_);
  nor _59420_ (_07749_, _06336_, _06269_);
  nor _59421_ (_07750_, _07749_, _07322_);
  not _59422_ (_07751_, _07750_);
  nor _59423_ (_07752_, _07751_, _07748_);
  and _59424_ (_07753_, _07680_, _07322_);
  nor _59425_ (_07754_, _07753_, _06279_);
  not _59426_ (_07755_, _07754_);
  nor _59427_ (_07756_, _07755_, _07752_);
  nor _59428_ (_07757_, _06278_, _06270_);
  nor _59429_ (_07758_, _07757_, _07756_);
  nor _59430_ (_07759_, _07758_, _06275_);
  and _59431_ (_07760_, _07690_, _06275_);
  not _59432_ (_07761_, _07760_);
  and _59433_ (_07762_, _07761_, _07343_);
  not _59434_ (_07763_, _07762_);
  nor _59435_ (_07764_, _07763_, _07759_);
  nor _59436_ (_07765_, _07343_, _06622_);
  nor _59437_ (_07766_, _07765_, _07330_);
  not _59438_ (_07767_, _07766_);
  nor _59439_ (_07768_, _07767_, _07764_);
  and _59440_ (_07769_, _07690_, _07330_);
  nor _59441_ (_07770_, _07769_, _07351_);
  not _59442_ (_07771_, _07770_);
  nor _59443_ (_07772_, _07771_, _07768_);
  and _59444_ (_07773_, _07351_, _06269_);
  nor _59445_ (_07774_, _07773_, _07350_);
  not _59446_ (_07775_, _07774_);
  nor _59447_ (_07776_, _07775_, _07772_);
  and _59448_ (_07777_, _07690_, _07350_);
  nor _59449_ (_07778_, _07777_, _07360_);
  not _59450_ (_07779_, _07778_);
  nor _59451_ (_07780_, _07779_, _07776_);
  or _59452_ (_07781_, _07780_, _07359_);
  nor _59453_ (_07782_, _07781_, _07682_);
  not _59454_ (_07783_, _07367_);
  and _59455_ (_07784_, _07359_, _06622_);
  nor _59456_ (_07785_, _07784_, _07783_);
  not _59457_ (_07786_, _07785_);
  nor _59458_ (_07787_, _07786_, _07782_);
  nor _59459_ (_07788_, _07690_, _07367_);
  nor _59460_ (_07789_, _07788_, _06272_);
  not _59461_ (_07790_, _07789_);
  nor _59462_ (_07791_, _07790_, _07787_);
  and _59463_ (_07792_, _06272_, _07741_);
  or _59464_ (_07793_, _07792_, _07055_);
  nor _59465_ (_07794_, _07793_, _07791_);
  or _59466_ (_07795_, _07794_, _07379_);
  nor _59467_ (_07796_, _07795_, _07681_);
  and _59468_ (_07797_, _07379_, _06622_);
  nor _59469_ (_07798_, _07797_, _07796_);
  not _59470_ (_07799_, _06727_);
  and _59471_ (_07800_, _07379_, _07799_);
  and _59472_ (_07801_, _06686_, _05989_);
  nor _59473_ (_07802_, _07684_, \oc8051_golden_model_1.SP [2]);
  nor _59474_ (_07803_, _07802_, _07685_);
  not _59475_ (_07804_, _07803_);
  nor _59476_ (_07805_, _07804_, _06016_);
  and _59477_ (_07806_, _07799_, _06279_);
  and _59478_ (_07807_, _06686_, _06339_);
  and _59479_ (_07808_, _07803_, _06351_);
  and _59480_ (_07809_, _07276_, _07799_);
  nand _59481_ (_07810_, _07061_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand _59482_ (_07811_, _07199_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _59483_ (_07812_, _07811_, _07198_);
  nand _59484_ (_07813_, _07812_, _07810_);
  nand _59485_ (_07814_, _07199_, \oc8051_golden_model_1.IRAM[3] [2]);
  nand _59486_ (_07815_, _07061_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _59487_ (_07816_, _07815_, _07204_);
  nand _59488_ (_07817_, _07816_, _07814_);
  nand _59489_ (_07818_, _07817_, _07813_);
  nand _59490_ (_07819_, _07818_, _06841_);
  nand _59491_ (_07820_, _07199_, \oc8051_golden_model_1.IRAM[7] [2]);
  nand _59492_ (_07821_, _07061_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _59493_ (_07822_, _07821_, _07204_);
  nand _59494_ (_07823_, _07822_, _07820_);
  nand _59495_ (_07824_, _07061_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand _59496_ (_07825_, _07199_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _59497_ (_07826_, _07825_, _07198_);
  nand _59498_ (_07827_, _07826_, _07824_);
  nand _59499_ (_07828_, _07827_, _07823_);
  nand _59500_ (_07829_, _07828_, _07210_);
  nand _59501_ (_07830_, _07829_, _07819_);
  nand _59502_ (_07831_, _07830_, _06654_);
  nand _59503_ (_07832_, _07199_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _59504_ (_07833_, _07061_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _59505_ (_07834_, _07833_, _07204_);
  nand _59506_ (_07835_, _07834_, _07832_);
  nand _59507_ (_07836_, _07061_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _59508_ (_07837_, _07199_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _59509_ (_07838_, _07837_, _07198_);
  nand _59510_ (_07839_, _07838_, _07836_);
  nand _59511_ (_07840_, _07839_, _07835_);
  nand _59512_ (_07841_, _07840_, _06841_);
  nand _59513_ (_07842_, _07199_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _59514_ (_07843_, _07061_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _59515_ (_07844_, _07843_, _07204_);
  nand _59516_ (_07845_, _07844_, _07842_);
  nand _59517_ (_07846_, _07061_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _59518_ (_07847_, _07199_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _59519_ (_07848_, _07847_, _07198_);
  nand _59520_ (_07849_, _07848_, _07846_);
  nand _59521_ (_07850_, _07849_, _07845_);
  nand _59522_ (_07851_, _07850_, _07210_);
  nand _59523_ (_07852_, _07851_, _07841_);
  nand _59524_ (_07853_, _07852_, _07224_);
  nand _59525_ (_07854_, _07853_, _07831_);
  or _59526_ (_07855_, _07854_, _05992_);
  and _59527_ (_07856_, _07855_, _07576_);
  and _59528_ (_07857_, _07261_, _06727_);
  nor _59529_ (_07858_, _07857_, _07856_);
  and _59530_ (_07859_, _07804_, _06816_);
  and _59531_ (_07860_, _06314_, _06355_);
  nor _59532_ (_07861_, _07860_, _07859_);
  and _59533_ (_07862_, _07861_, _07858_);
  and _59534_ (_07863_, _07854_, _07269_);
  nor _59535_ (_07864_, _07863_, _07276_);
  and _59536_ (_07865_, _07864_, _07862_);
  nor _59537_ (_07866_, _07865_, _07809_);
  and _59538_ (_07867_, _07274_, _06685_);
  or _59539_ (_07868_, _07867_, _07866_);
  nor _59540_ (_07869_, _07803_, _06052_);
  nor _59541_ (_07870_, _07869_, _07284_);
  not _59542_ (_07871_, _07870_);
  nor _59543_ (_07872_, _07871_, _07868_);
  and _59544_ (_07873_, _07284_, _07799_);
  nor _59545_ (_07874_, _07873_, _07872_);
  and _59546_ (_07875_, _06314_, _06350_);
  nor _59547_ (_07876_, _07875_, _07874_);
  and _59548_ (_07877_, _07854_, _07289_);
  nor _59549_ (_07878_, _07877_, _07295_);
  and _59550_ (_07879_, _07878_, _07876_);
  and _59551_ (_07880_, _07295_, _07799_);
  nor _59552_ (_07881_, _07880_, _07879_);
  and _59553_ (_07882_, _06685_, _07294_);
  nor _59554_ (_07883_, _07882_, _07881_);
  and _59555_ (_07884_, _07883_, _07394_);
  nor _59556_ (_07885_, _07884_, _07808_);
  and _59557_ (_07886_, _06348_, _06685_);
  or _59558_ (_07887_, _07886_, _07885_);
  nor _59559_ (_07888_, _07803_, _06049_);
  and _59560_ (_07889_, _06323_, _06443_);
  or _59561_ (_07890_, _07889_, _07601_);
  nor _59562_ (_07891_, _07890_, _07888_);
  not _59563_ (_07892_, _07891_);
  nor _59564_ (_07893_, _07892_, _07887_);
  and _59565_ (_07894_, _07854_, _07309_);
  nor _59566_ (_07895_, _07894_, _07308_);
  and _59567_ (_07896_, _07895_, _07893_);
  nor _59568_ (_07897_, _07896_, _07807_);
  nor _59569_ (_07898_, _07897_, _06039_);
  and _59570_ (_07899_, _07803_, _06039_);
  nor _59571_ (_07900_, _07899_, _07898_);
  nor _59572_ (_07901_, _06336_, _07799_);
  and _59573_ (_07902_, _06314_, _06276_);
  nor _59574_ (_07903_, _07902_, _07901_);
  not _59575_ (_07904_, _07903_);
  nor _59576_ (_07905_, _07904_, _07900_);
  and _59577_ (_07906_, _07854_, _07322_);
  nor _59578_ (_07907_, _07906_, _06279_);
  and _59579_ (_07908_, _07907_, _07905_);
  nor _59580_ (_07909_, _07908_, _07806_);
  nor _59581_ (_07910_, _07909_, _06275_);
  nor _59582_ (_07911_, _07804_, _06009_);
  nor _59583_ (_07912_, _07911_, _07910_);
  nor _59584_ (_07913_, _07343_, _07799_);
  nor _59585_ (_07914_, _07913_, _07330_);
  not _59586_ (_07915_, _07914_);
  nor _59587_ (_07916_, _07915_, _07912_);
  nor _59588_ (_07917_, _07804_, _06018_);
  nor _59589_ (_07918_, _07917_, _07916_);
  and _59590_ (_07919_, _07351_, _06727_);
  nor _59591_ (_07920_, _07919_, _07350_);
  not _59592_ (_07921_, _07920_);
  nor _59593_ (_07922_, _07921_, _07918_);
  nor _59594_ (_07923_, _07922_, _07805_);
  and _59595_ (_07924_, _06314_, _05848_);
  nor _59596_ (_07925_, _07924_, _07923_);
  and _59597_ (_07926_, _07854_, _07360_);
  nor _59598_ (_07927_, _07926_, _07359_);
  and _59599_ (_07928_, _07927_, _07925_);
  and _59600_ (_07929_, _07359_, _07799_);
  nor _59601_ (_07930_, _07929_, _07928_);
  nor _59602_ (_07931_, _07803_, _07367_);
  nor _59603_ (_07932_, _07931_, _06272_);
  not _59604_ (_07933_, _07932_);
  nor _59605_ (_07934_, _07933_, _07930_);
  nor _59606_ (_07935_, _07934_, _07801_);
  nor _59607_ (_07936_, _07935_, _07591_);
  and _59608_ (_07937_, _07854_, _07055_);
  nor _59609_ (_07938_, _07937_, _07379_);
  and _59610_ (_07939_, _07938_, _07936_);
  nor _59611_ (_07940_, _07939_, _07800_);
  nor _59612_ (_07941_, _07940_, _07632_);
  not _59613_ (_07942_, _07941_);
  or _59614_ (_07943_, _07942_, _07798_);
  nor _59615_ (_07944_, _07943_, _07635_);
  nor _59616_ (_07945_, _07944_, _05659_);
  and _59617_ (_07946_, _06397_, _06238_);
  and _59618_ (_07947_, _07946_, _06685_);
  and _59619_ (_07948_, _07947_, _07093_);
  not _59620_ (_07949_, _07948_);
  and _59621_ (_07950_, _07127_, _06310_);
  not _59622_ (_07951_, _07950_);
  or _59623_ (_07952_, _06727_, _06269_);
  or _59624_ (_07953_, _07952_, _07951_);
  nor _59625_ (_07954_, _07953_, _07949_);
  and _59626_ (_07955_, _07954_, \oc8051_golden_model_1.TH0 [7]);
  and _59627_ (_07956_, _07127_, _06311_);
  and _59628_ (_07957_, _07956_, _06727_);
  and _59629_ (_07958_, _07957_, _06622_);
  not _59630_ (_07959_, _07093_);
  and _59631_ (_07960_, _07959_, _06685_);
  and _59632_ (_07961_, _07960_, _07946_);
  and _59633_ (_07962_, _07961_, _07958_);
  and _59634_ (_07963_, _07962_, \oc8051_golden_model_1.SBUF [7]);
  nor _59635_ (_07964_, _07963_, _07955_);
  and _59636_ (_07965_, _07958_, _07948_);
  and _59637_ (_07966_, _07965_, \oc8051_golden_model_1.TMOD [7]);
  and _59638_ (_07967_, _07950_, _06727_);
  and _59639_ (_07968_, _07967_, _06622_);
  and _59640_ (_07969_, _07968_, _07961_);
  and _59641_ (_07970_, _07969_, \oc8051_golden_model_1.SCON [7]);
  nor _59642_ (_07971_, _07970_, _07966_);
  and _59643_ (_07972_, _07971_, _07964_);
  nor _59644_ (_07973_, _07127_, _06311_);
  nand _59645_ (_07974_, _06727_, _06622_);
  nor _59646_ (_07975_, _07974_, _07949_);
  and _59647_ (_07976_, _07975_, _07973_);
  and _59648_ (_07977_, _07976_, \oc8051_golden_model_1.TL0 [7]);
  not _59649_ (_07978_, _07977_);
  not _59650_ (_07979_, _07956_);
  or _59651_ (_07980_, _07979_, _07952_);
  nor _59652_ (_07981_, _07980_, _07949_);
  and _59653_ (_07982_, _07981_, \oc8051_golden_model_1.TH1 [7]);
  not _59654_ (_07983_, _06685_);
  and _59655_ (_07984_, _07093_, _07983_);
  and _59656_ (_07985_, _07984_, _07946_);
  and _59657_ (_07986_, _07985_, _07968_);
  and _59658_ (_07987_, _07986_, \oc8051_golden_model_1.IE [7]);
  nor _59659_ (_07988_, _07987_, _07982_);
  and _59660_ (_07989_, _07988_, _07978_);
  nor _59661_ (_07990_, _07127_, _06310_);
  and _59662_ (_07991_, _07990_, _07975_);
  and _59663_ (_07992_, _07991_, \oc8051_golden_model_1.TL1 [7]);
  and _59664_ (_07993_, _07948_, _06269_);
  and _59665_ (_07994_, _07990_, _06727_);
  and _59666_ (_07995_, _07994_, _07993_);
  and _59667_ (_07996_, _07995_, \oc8051_golden_model_1.DPH [7]);
  nor _59668_ (_07997_, _07996_, _07992_);
  and _59669_ (_07998_, _07997_, _07989_);
  and _59670_ (_07999_, _07998_, _07972_);
  and _59671_ (_08000_, _07973_, _06727_);
  and _59672_ (_08001_, _08000_, _07993_);
  and _59673_ (_08002_, _08001_, \oc8051_golden_model_1.DPL [7]);
  not _59674_ (_08003_, _08002_);
  and _59675_ (_08004_, _07993_, _07957_);
  and _59676_ (_08005_, _08004_, \oc8051_golden_model_1.SP [7]);
  and _59677_ (_08006_, _07968_, _07948_);
  and _59678_ (_08007_, _08006_, \oc8051_golden_model_1.TCON [7]);
  nor _59679_ (_08008_, _08007_, _08005_);
  and _59680_ (_08009_, _08008_, _08003_);
  nand _59681_ (_08010_, _06727_, _06269_);
  nor _59682_ (_08011_, _08010_, _07951_);
  nor _59683_ (_08012_, _06397_, _06366_);
  and _59684_ (_08013_, _08012_, _07960_);
  and _59685_ (_08014_, _08013_, _08011_);
  and _59686_ (_08015_, _08014_, \oc8051_golden_model_1.PSW [7]);
  and _59687_ (_08016_, _08012_, _07984_);
  and _59688_ (_08017_, _08016_, _08011_);
  and _59689_ (_08018_, _08017_, \oc8051_golden_model_1.ACC [7]);
  nor _59690_ (_08019_, _08018_, _08015_);
  nor _59691_ (_08020_, _07093_, _06685_);
  and _59692_ (_08021_, _08020_, _07946_);
  and _59693_ (_08022_, _08021_, _07968_);
  and _59694_ (_08023_, _08022_, \oc8051_golden_model_1.IP [7]);
  and _59695_ (_08024_, _08020_, _08012_);
  and _59696_ (_08025_, _08024_, _08011_);
  and _59697_ (_08026_, _08025_, \oc8051_golden_model_1.B [7]);
  nor _59698_ (_08027_, _08026_, _08023_);
  and _59699_ (_08028_, _08027_, _08019_);
  and _59700_ (_08029_, _08011_, _07961_);
  and _59701_ (_08030_, _08029_, \oc8051_golden_model_1.P1INREG [7]);
  not _59702_ (_08031_, _08030_);
  and _59703_ (_08032_, _08011_, _07985_);
  and _59704_ (_08033_, _08032_, \oc8051_golden_model_1.P2INREG [7]);
  and _59705_ (_08034_, _08021_, _08011_);
  and _59706_ (_08035_, _08034_, \oc8051_golden_model_1.P3INREG [7]);
  nor _59707_ (_08036_, _08035_, _08033_);
  and _59708_ (_08037_, _08036_, _08031_);
  and _59709_ (_08038_, _08037_, _08028_);
  and _59710_ (_08039_, _08011_, _07948_);
  and _59711_ (_08040_, _08039_, \oc8051_golden_model_1.P0INREG [7]);
  and _59712_ (_08041_, _07990_, _07799_);
  and _59713_ (_08042_, _08041_, _07993_);
  and _59714_ (_08043_, _08042_, \oc8051_golden_model_1.PCON [7]);
  nor _59715_ (_08044_, _08043_, _08040_);
  and _59716_ (_08045_, _08044_, _08038_);
  and _59717_ (_08046_, _08045_, _08009_);
  and _59718_ (_08047_, _08046_, _07999_);
  not _59719_ (_08048_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _59720_ (_08049_, _07199_, _08048_);
  not _59721_ (_08050_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _59722_ (_08051_, _07061_, _08050_);
  and _59723_ (_08052_, _08051_, _07198_);
  nand _59724_ (_08053_, _08052_, _08049_);
  not _59725_ (_08054_, \oc8051_golden_model_1.IRAM[3] [7]);
  or _59726_ (_08055_, _07061_, _08054_);
  not _59727_ (_08056_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _59728_ (_08057_, _07199_, _08056_);
  and _59729_ (_08058_, _08057_, _07204_);
  nand _59730_ (_08059_, _08058_, _08055_);
  nand _59731_ (_08060_, _08059_, _08053_);
  nand _59732_ (_08061_, _08060_, _06841_);
  not _59733_ (_08062_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _59734_ (_08063_, _07061_, _08062_);
  not _59735_ (_08064_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _59736_ (_08065_, _07199_, _08064_);
  and _59737_ (_08066_, _08065_, _07204_);
  nand _59738_ (_08067_, _08066_, _08063_);
  not _59739_ (_08068_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _59740_ (_08069_, _07199_, _08068_);
  not _59741_ (_08070_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _59742_ (_08071_, _07061_, _08070_);
  and _59743_ (_08072_, _08071_, _07198_);
  nand _59744_ (_08073_, _08072_, _08069_);
  nand _59745_ (_08074_, _08073_, _08067_);
  nand _59746_ (_08075_, _08074_, _07210_);
  nand _59747_ (_08076_, _08075_, _08061_);
  nand _59748_ (_08077_, _08076_, _06654_);
  not _59749_ (_08078_, \oc8051_golden_model_1.IRAM[11] [7]);
  or _59750_ (_08079_, _07061_, _08078_);
  not _59751_ (_08080_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _59752_ (_08081_, _07199_, _08080_);
  and _59753_ (_08082_, _08081_, _07204_);
  nand _59754_ (_08083_, _08082_, _08079_);
  not _59755_ (_08084_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _59756_ (_08085_, _07199_, _08084_);
  not _59757_ (_08086_, \oc8051_golden_model_1.IRAM[9] [7]);
  or _59758_ (_08087_, _07061_, _08086_);
  and _59759_ (_08088_, _08087_, _07198_);
  nand _59760_ (_08089_, _08088_, _08085_);
  nand _59761_ (_08090_, _08089_, _08083_);
  nand _59762_ (_08091_, _08090_, _06841_);
  or _59763_ (_08092_, _07061_, _05659_);
  not _59764_ (_08093_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _59765_ (_08094_, _07199_, _08093_);
  and _59766_ (_08095_, _08094_, _07204_);
  nand _59767_ (_08096_, _08095_, _08092_);
  not _59768_ (_08097_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _59769_ (_08098_, _07199_, _08097_);
  not _59770_ (_08099_, \oc8051_golden_model_1.IRAM[13] [7]);
  or _59771_ (_08100_, _07061_, _08099_);
  and _59772_ (_08101_, _08100_, _07198_);
  nand _59773_ (_08102_, _08101_, _08098_);
  nand _59774_ (_08103_, _08102_, _08096_);
  nand _59775_ (_08104_, _08103_, _07210_);
  nand _59776_ (_08105_, _08104_, _08091_);
  nand _59777_ (_08106_, _08105_, _07224_);
  nand _59778_ (_08107_, _08106_, _08077_);
  or _59779_ (_08108_, _08107_, _06238_);
  and _59780_ (_08109_, _08108_, _08047_);
  not _59781_ (_08110_, _08109_);
  and _59782_ (_08111_, _08022_, \oc8051_golden_model_1.IP [6]);
  not _59783_ (_08112_, _08111_);
  and _59784_ (_08113_, _08014_, \oc8051_golden_model_1.PSW [6]);
  not _59785_ (_08114_, _08113_);
  and _59786_ (_08115_, _08017_, \oc8051_golden_model_1.ACC [6]);
  and _59787_ (_08116_, _08025_, \oc8051_golden_model_1.B [6]);
  nor _59788_ (_08117_, _08116_, _08115_);
  and _59789_ (_08118_, _08117_, _08114_);
  and _59790_ (_08119_, _08118_, _08112_);
  and _59791_ (_08120_, _08006_, \oc8051_golden_model_1.TCON [6]);
  and _59792_ (_08121_, _07954_, \oc8051_golden_model_1.TH0 [6]);
  nor _59793_ (_08122_, _08121_, _08120_);
  and _59794_ (_08123_, _07991_, \oc8051_golden_model_1.TL1 [6]);
  and _59795_ (_08124_, _08029_, \oc8051_golden_model_1.P1INREG [6]);
  nor _59796_ (_08125_, _08124_, _08123_);
  and _59797_ (_08126_, _08125_, _08122_);
  and _59798_ (_08127_, _07969_, \oc8051_golden_model_1.SCON [6]);
  and _59799_ (_08128_, _07981_, \oc8051_golden_model_1.TH1 [6]);
  nor _59800_ (_08129_, _08128_, _08127_);
  and _59801_ (_08130_, _07965_, \oc8051_golden_model_1.TMOD [6]);
  not _59802_ (_08131_, _07973_);
  or _59803_ (_08132_, _08131_, _07974_);
  nor _59804_ (_08133_, _08132_, _07949_);
  and _59805_ (_08134_, _08133_, \oc8051_golden_model_1.TL0 [6]);
  nor _59806_ (_08135_, _08134_, _08130_);
  and _59807_ (_08136_, _08135_, _08129_);
  and _59808_ (_08137_, _08136_, _08126_);
  and _59809_ (_08138_, _08137_, _08119_);
  and _59810_ (_08139_, _08042_, \oc8051_golden_model_1.PCON [6]);
  not _59811_ (_08140_, _08139_);
  and _59812_ (_08141_, _07962_, \oc8051_golden_model_1.SBUF [6]);
  and _59813_ (_08142_, _07986_, \oc8051_golden_model_1.IE [6]);
  nor _59814_ (_08143_, _08142_, _08141_);
  and _59815_ (_08144_, _08143_, _08140_);
  and _59816_ (_08145_, _08032_, \oc8051_golden_model_1.P2INREG [6]);
  and _59817_ (_08146_, _08034_, \oc8051_golden_model_1.P3INREG [6]);
  nor _59818_ (_08147_, _08146_, _08145_);
  and _59819_ (_08148_, _08147_, _08144_);
  and _59820_ (_08149_, _08039_, \oc8051_golden_model_1.P0INREG [6]);
  not _59821_ (_08150_, _08149_);
  not _59822_ (_08151_, _07990_);
  nor _59823_ (_08152_, _08010_, _08151_);
  and _59824_ (_08153_, _08152_, _07948_);
  and _59825_ (_08154_, _08153_, \oc8051_golden_model_1.DPH [6]);
  not _59826_ (_08155_, _08154_);
  and _59827_ (_08156_, _08004_, \oc8051_golden_model_1.SP [6]);
  or _59828_ (_08157_, _08010_, _08131_);
  nor _59829_ (_08158_, _08157_, _07949_);
  and _59830_ (_08159_, _08158_, \oc8051_golden_model_1.DPL [6]);
  nor _59831_ (_08160_, _08159_, _08156_);
  and _59832_ (_08161_, _08160_, _08155_);
  and _59833_ (_08162_, _08161_, _08150_);
  and _59834_ (_08163_, _08162_, _08148_);
  and _59835_ (_08164_, _08163_, _08138_);
  nand _59836_ (_08165_, _07061_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand _59837_ (_08166_, _07199_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _59838_ (_08167_, _08166_, _07198_);
  nand _59839_ (_08168_, _08167_, _08165_);
  nand _59840_ (_08169_, _07199_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand _59841_ (_08170_, _07061_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _59842_ (_08171_, _08170_, _07204_);
  nand _59843_ (_08172_, _08171_, _08169_);
  nand _59844_ (_08173_, _08172_, _08168_);
  nand _59845_ (_08174_, _08173_, _06841_);
  nand _59846_ (_08175_, _07199_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand _59847_ (_08176_, _07061_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _59848_ (_08177_, _08176_, _07204_);
  nand _59849_ (_08178_, _08177_, _08175_);
  nand _59850_ (_08179_, _07061_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand _59851_ (_08180_, _07199_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _59852_ (_08181_, _08180_, _07198_);
  nand _59853_ (_08182_, _08181_, _08179_);
  nand _59854_ (_08183_, _08182_, _08178_);
  nand _59855_ (_08184_, _08183_, _07210_);
  nand _59856_ (_08185_, _08184_, _08174_);
  nand _59857_ (_08186_, _08185_, _06654_);
  nand _59858_ (_08187_, _07199_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _59859_ (_08188_, _07061_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _59860_ (_08189_, _08188_, _07204_);
  nand _59861_ (_08190_, _08189_, _08187_);
  nand _59862_ (_08191_, _07061_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _59863_ (_08192_, _07199_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _59864_ (_08193_, _08192_, _07198_);
  nand _59865_ (_08194_, _08193_, _08191_);
  nand _59866_ (_08195_, _08194_, _08190_);
  nand _59867_ (_08196_, _08195_, _06841_);
  nand _59868_ (_08197_, _07199_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _59869_ (_08198_, _07061_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _59870_ (_08199_, _08198_, _07204_);
  nand _59871_ (_08200_, _08199_, _08197_);
  nand _59872_ (_08201_, _07061_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _59873_ (_08202_, _07199_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _59874_ (_08203_, _08202_, _07198_);
  nand _59875_ (_08204_, _08203_, _08201_);
  nand _59876_ (_08205_, _08204_, _08200_);
  nand _59877_ (_08206_, _08205_, _07210_);
  nand _59878_ (_08207_, _08206_, _08196_);
  nand _59879_ (_08208_, _08207_, _07224_);
  nand _59880_ (_08209_, _08208_, _08186_);
  or _59881_ (_08210_, _08209_, _06238_);
  and _59882_ (_08211_, _08210_, _08164_);
  not _59883_ (_08212_, _08211_);
  and _59884_ (_08213_, _07965_, \oc8051_golden_model_1.TMOD [5]);
  and _59885_ (_08214_, _07981_, \oc8051_golden_model_1.TH1 [5]);
  nor _59886_ (_08215_, _08214_, _08213_);
  and _59887_ (_08216_, _07954_, \oc8051_golden_model_1.TH0 [5]);
  and _59888_ (_08217_, _07969_, \oc8051_golden_model_1.SCON [5]);
  nor _59889_ (_08218_, _08217_, _08216_);
  and _59890_ (_08219_, _08218_, _08215_);
  and _59891_ (_08220_, _07995_, \oc8051_golden_model_1.DPH [5]);
  not _59892_ (_08221_, _08220_);
  and _59893_ (_08222_, _07991_, \oc8051_golden_model_1.TL1 [5]);
  and _59894_ (_08223_, _07976_, \oc8051_golden_model_1.TL0 [5]);
  nor _59895_ (_08224_, _08223_, _08222_);
  and _59896_ (_08225_, _08224_, _08221_);
  and _59897_ (_08226_, _08225_, _08219_);
  and _59898_ (_08227_, _08042_, \oc8051_golden_model_1.PCON [5]);
  not _59899_ (_08228_, _08227_);
  and _59900_ (_08229_, _08022_, \oc8051_golden_model_1.IP [5]);
  not _59901_ (_08230_, _08229_);
  and _59902_ (_08231_, _08014_, \oc8051_golden_model_1.PSW [5]);
  and _59903_ (_08232_, _08017_, \oc8051_golden_model_1.ACC [5]);
  nor _59904_ (_08233_, _08232_, _08231_);
  and _59905_ (_08234_, _08233_, _08230_);
  and _59906_ (_08235_, _07962_, \oc8051_golden_model_1.SBUF [5]);
  not _59907_ (_08236_, _08235_);
  and _59908_ (_08237_, _07986_, \oc8051_golden_model_1.IE [5]);
  and _59909_ (_08238_, _08025_, \oc8051_golden_model_1.B [5]);
  nor _59910_ (_08239_, _08238_, _08237_);
  and _59911_ (_08240_, _08239_, _08236_);
  and _59912_ (_08241_, _08240_, _08234_);
  and _59913_ (_08242_, _08241_, _08228_);
  and _59914_ (_08243_, _08001_, \oc8051_golden_model_1.DPL [5]);
  not _59915_ (_08244_, _08243_);
  and _59916_ (_08245_, _08004_, \oc8051_golden_model_1.SP [5]);
  and _59917_ (_08246_, _08006_, \oc8051_golden_model_1.TCON [5]);
  nor _59918_ (_08247_, _08246_, _08245_);
  and _59919_ (_08248_, _08247_, _08244_);
  and _59920_ (_08249_, _08039_, \oc8051_golden_model_1.P0INREG [5]);
  not _59921_ (_08250_, _08249_);
  and _59922_ (_08251_, _08029_, \oc8051_golden_model_1.P1INREG [5]);
  not _59923_ (_08252_, _08251_);
  and _59924_ (_08253_, _08032_, \oc8051_golden_model_1.P2INREG [5]);
  and _59925_ (_08254_, _08034_, \oc8051_golden_model_1.P3INREG [5]);
  nor _59926_ (_08255_, _08254_, _08253_);
  and _59927_ (_08256_, _08255_, _08252_);
  and _59928_ (_08257_, _08256_, _08250_);
  and _59929_ (_08258_, _08257_, _08248_);
  and _59930_ (_08259_, _08258_, _08242_);
  and _59931_ (_08260_, _08259_, _08226_);
  nand _59932_ (_08261_, _07061_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand _59933_ (_08262_, _07199_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _59934_ (_08263_, _08262_, _07198_);
  nand _59935_ (_08264_, _08263_, _08261_);
  nand _59936_ (_08265_, _07199_, \oc8051_golden_model_1.IRAM[3] [5]);
  nand _59937_ (_08266_, _07061_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _59938_ (_08267_, _08266_, _07204_);
  nand _59939_ (_08268_, _08267_, _08265_);
  nand _59940_ (_08269_, _08268_, _08264_);
  nand _59941_ (_08270_, _08269_, _06841_);
  nand _59942_ (_08271_, _07199_, \oc8051_golden_model_1.IRAM[7] [5]);
  nand _59943_ (_08272_, _07061_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _59944_ (_08273_, _08272_, _07204_);
  nand _59945_ (_08274_, _08273_, _08271_);
  nand _59946_ (_08275_, _07061_, \oc8051_golden_model_1.IRAM[4] [5]);
  nand _59947_ (_08276_, _07199_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _59948_ (_08277_, _08276_, _07198_);
  nand _59949_ (_08278_, _08277_, _08275_);
  nand _59950_ (_08279_, _08278_, _08274_);
  nand _59951_ (_08280_, _08279_, _07210_);
  nand _59952_ (_08281_, _08280_, _08270_);
  nand _59953_ (_08282_, _08281_, _06654_);
  nand _59954_ (_08283_, _07199_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _59955_ (_08284_, _07061_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _59956_ (_08285_, _08284_, _07204_);
  nand _59957_ (_08286_, _08285_, _08283_);
  nand _59958_ (_08287_, _07061_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand _59959_ (_08288_, _07199_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _59960_ (_08289_, _08288_, _07198_);
  nand _59961_ (_08290_, _08289_, _08287_);
  nand _59962_ (_08291_, _08290_, _08286_);
  nand _59963_ (_08292_, _08291_, _06841_);
  nand _59964_ (_08293_, _07199_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _59965_ (_08294_, _07061_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _59966_ (_08295_, _08294_, _07204_);
  nand _59967_ (_08296_, _08295_, _08293_);
  nand _59968_ (_08297_, _07061_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand _59969_ (_08298_, _07199_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _59970_ (_08299_, _08298_, _07198_);
  nand _59971_ (_08300_, _08299_, _08297_);
  nand _59972_ (_08301_, _08300_, _08296_);
  nand _59973_ (_08302_, _08301_, _07210_);
  nand _59974_ (_08303_, _08302_, _08292_);
  nand _59975_ (_08304_, _08303_, _07224_);
  nand _59976_ (_08305_, _08304_, _08282_);
  or _59977_ (_08306_, _08305_, _06238_);
  and _59978_ (_08307_, _08306_, _08260_);
  not _59979_ (_08308_, _08307_);
  and _59980_ (_08309_, _07965_, \oc8051_golden_model_1.TMOD [3]);
  and _59981_ (_08310_, _07981_, \oc8051_golden_model_1.TH1 [3]);
  nor _59982_ (_08311_, _08310_, _08309_);
  and _59983_ (_08312_, _07954_, \oc8051_golden_model_1.TH0 [3]);
  and _59984_ (_08313_, _07969_, \oc8051_golden_model_1.SCON [3]);
  nor _59985_ (_08314_, _08313_, _08312_);
  and _59986_ (_08315_, _08314_, _08311_);
  and _59987_ (_08316_, _07995_, \oc8051_golden_model_1.DPH [3]);
  not _59988_ (_08317_, _08316_);
  and _59989_ (_08318_, _07991_, \oc8051_golden_model_1.TL1 [3]);
  and _59990_ (_08319_, _07976_, \oc8051_golden_model_1.TL0 [3]);
  nor _59991_ (_08320_, _08319_, _08318_);
  and _59992_ (_08321_, _08320_, _08317_);
  and _59993_ (_08322_, _08321_, _08315_);
  and _59994_ (_08323_, _08042_, \oc8051_golden_model_1.PCON [3]);
  not _59995_ (_08324_, _08323_);
  and _59996_ (_08325_, _08022_, \oc8051_golden_model_1.IP [3]);
  not _59997_ (_08326_, _08325_);
  and _59998_ (_08327_, _08014_, \oc8051_golden_model_1.PSW [3]);
  and _59999_ (_08328_, _08017_, \oc8051_golden_model_1.ACC [3]);
  nor _60000_ (_08329_, _08328_, _08327_);
  and _60001_ (_08330_, _08329_, _08326_);
  and _60002_ (_08331_, _07962_, \oc8051_golden_model_1.SBUF [3]);
  not _60003_ (_08332_, _08331_);
  and _60004_ (_08333_, _07986_, \oc8051_golden_model_1.IE [3]);
  and _60005_ (_08334_, _08025_, \oc8051_golden_model_1.B [3]);
  nor _60006_ (_08335_, _08334_, _08333_);
  and _60007_ (_08336_, _08335_, _08332_);
  and _60008_ (_08337_, _08336_, _08330_);
  and _60009_ (_08338_, _08337_, _08324_);
  and _60010_ (_08339_, _08001_, \oc8051_golden_model_1.DPL [3]);
  not _60011_ (_08340_, _08339_);
  and _60012_ (_08341_, _08004_, \oc8051_golden_model_1.SP [3]);
  and _60013_ (_08342_, _08006_, \oc8051_golden_model_1.TCON [3]);
  nor _60014_ (_08343_, _08342_, _08341_);
  and _60015_ (_08344_, _08343_, _08340_);
  and _60016_ (_08345_, _08039_, \oc8051_golden_model_1.P0INREG [3]);
  not _60017_ (_08346_, _08345_);
  and _60018_ (_08347_, _08029_, \oc8051_golden_model_1.P1INREG [3]);
  not _60019_ (_08348_, _08347_);
  and _60020_ (_08349_, _08032_, \oc8051_golden_model_1.P2INREG [3]);
  and _60021_ (_08350_, _08034_, \oc8051_golden_model_1.P3INREG [3]);
  nor _60022_ (_08351_, _08350_, _08349_);
  and _60023_ (_08352_, _08351_, _08348_);
  and _60024_ (_08353_, _08352_, _08346_);
  and _60025_ (_08354_, _08353_, _08344_);
  and _60026_ (_08355_, _08354_, _08338_);
  and _60027_ (_08356_, _08355_, _08322_);
  or _60028_ (_08357_, _07680_, _06238_);
  and _60029_ (_08358_, _08357_, _08356_);
  not _60030_ (_08359_, _08358_);
  and _60031_ (_08360_, _08014_, \oc8051_golden_model_1.PSW [1]);
  and _60032_ (_08361_, _08025_, \oc8051_golden_model_1.B [1]);
  nor _60033_ (_08362_, _08361_, _08360_);
  and _60034_ (_08363_, _08022_, \oc8051_golden_model_1.IP [1]);
  and _60035_ (_08364_, _08017_, \oc8051_golden_model_1.ACC [1]);
  nor _60036_ (_08365_, _08364_, _08363_);
  and _60037_ (_08366_, _08365_, _08362_);
  and _60038_ (_08367_, _08039_, \oc8051_golden_model_1.P0INREG [1]);
  and _60039_ (_08368_, _08153_, \oc8051_golden_model_1.DPH [1]);
  nor _60040_ (_08369_, _08368_, _08367_);
  and _60041_ (_08370_, _08369_, _08366_);
  and _60042_ (_08371_, _08042_, \oc8051_golden_model_1.PCON [1]);
  not _60043_ (_08372_, _08371_);
  and _60044_ (_08373_, _07962_, \oc8051_golden_model_1.SBUF [1]);
  and _60045_ (_08374_, _07986_, \oc8051_golden_model_1.IE [1]);
  nor _60046_ (_08375_, _08374_, _08373_);
  and _60047_ (_08376_, _08375_, _08372_);
  and _60048_ (_08377_, _08032_, \oc8051_golden_model_1.P2INREG [1]);
  and _60049_ (_08378_, _08034_, \oc8051_golden_model_1.P3INREG [1]);
  nor _60050_ (_08379_, _08378_, _08377_);
  and _60051_ (_08380_, _08379_, _08376_);
  and _60052_ (_08381_, _07954_, \oc8051_golden_model_1.TH0 [1]);
  and _60053_ (_08382_, _08006_, \oc8051_golden_model_1.TCON [1]);
  nor _60054_ (_08383_, _08382_, _08381_);
  and _60055_ (_08384_, _07991_, \oc8051_golden_model_1.TL1 [1]);
  and _60056_ (_08385_, _08029_, \oc8051_golden_model_1.P1INREG [1]);
  nor _60057_ (_08386_, _08385_, _08384_);
  and _60058_ (_08387_, _08386_, _08383_);
  and _60059_ (_08388_, _07969_, \oc8051_golden_model_1.SCON [1]);
  and _60060_ (_08389_, _07981_, \oc8051_golden_model_1.TH1 [1]);
  nor _60061_ (_08390_, _08389_, _08388_);
  and _60062_ (_08391_, _07965_, \oc8051_golden_model_1.TMOD [1]);
  and _60063_ (_08392_, _08133_, \oc8051_golden_model_1.TL0 [1]);
  nor _60064_ (_08393_, _08392_, _08391_);
  and _60065_ (_08394_, _08393_, _08390_);
  and _60066_ (_08395_, _08394_, _08387_);
  and _60067_ (_08396_, _08004_, \oc8051_golden_model_1.SP [1]);
  and _60068_ (_08397_, _08158_, \oc8051_golden_model_1.DPL [1]);
  nor _60069_ (_08398_, _08397_, _08396_);
  and _60070_ (_08399_, _08398_, _08395_);
  and _60071_ (_08400_, _08399_, _08380_);
  and _60072_ (_08401_, _08400_, _08370_);
  or _60073_ (_08402_, _07448_, _06238_);
  and _60074_ (_08403_, _08402_, _08401_);
  not _60075_ (_08404_, _08403_);
  and _60076_ (_08405_, _07954_, \oc8051_golden_model_1.TH0 [0]);
  and _60077_ (_08406_, _07981_, \oc8051_golden_model_1.TH1 [0]);
  nor _60078_ (_08407_, _08406_, _08405_);
  and _60079_ (_08408_, _07965_, \oc8051_golden_model_1.TMOD [0]);
  and _60080_ (_08409_, _07969_, \oc8051_golden_model_1.SCON [0]);
  nor _60081_ (_08410_, _08409_, _08408_);
  and _60082_ (_08411_, _08410_, _08407_);
  and _60083_ (_08412_, _08022_, \oc8051_golden_model_1.IP [0]);
  and _60084_ (_08413_, _08017_, \oc8051_golden_model_1.ACC [0]);
  nor _60085_ (_08414_, _08413_, _08412_);
  and _60086_ (_08415_, _08014_, \oc8051_golden_model_1.PSW [0]);
  and _60087_ (_08416_, _08025_, \oc8051_golden_model_1.B [0]);
  nor _60088_ (_08417_, _08416_, _08415_);
  and _60089_ (_08418_, _08417_, _08414_);
  not _60090_ (_08419_, _08418_);
  and _60091_ (_08420_, _07976_, \oc8051_golden_model_1.TL0 [0]);
  nor _60092_ (_08421_, _08420_, _08419_);
  and _60093_ (_08422_, _07991_, \oc8051_golden_model_1.TL1 [0]);
  and _60094_ (_08423_, _07995_, \oc8051_golden_model_1.DPH [0]);
  nor _60095_ (_08424_, _08423_, _08422_);
  and _60096_ (_08425_, _08424_, _08421_);
  and _60097_ (_08426_, _08425_, _08411_);
  and _60098_ (_08427_, _08004_, \oc8051_golden_model_1.SP [0]);
  not _60099_ (_08428_, _08427_);
  and _60100_ (_08429_, _08006_, \oc8051_golden_model_1.TCON [0]);
  and _60101_ (_08430_, _08001_, \oc8051_golden_model_1.DPL [0]);
  nor _60102_ (_08431_, _08430_, _08429_);
  and _60103_ (_08432_, _08431_, _08428_);
  and _60104_ (_08433_, _08042_, \oc8051_golden_model_1.PCON [0]);
  not _60105_ (_08434_, _08433_);
  and _60106_ (_08435_, _07962_, \oc8051_golden_model_1.SBUF [0]);
  and _60107_ (_08436_, _07986_, \oc8051_golden_model_1.IE [0]);
  nor _60108_ (_08437_, _08436_, _08435_);
  and _60109_ (_08438_, _08437_, _08434_);
  and _60110_ (_08439_, _08039_, \oc8051_golden_model_1.P0INREG [0]);
  not _60111_ (_08440_, _08439_);
  and _60112_ (_08441_, _08029_, \oc8051_golden_model_1.P1INREG [0]);
  not _60113_ (_08442_, _08441_);
  and _60114_ (_08443_, _08032_, \oc8051_golden_model_1.P2INREG [0]);
  and _60115_ (_08444_, _08034_, \oc8051_golden_model_1.P3INREG [0]);
  nor _60116_ (_08445_, _08444_, _08443_);
  and _60117_ (_08446_, _08445_, _08442_);
  and _60118_ (_08447_, _08446_, _08440_);
  and _60119_ (_08448_, _08447_, _08438_);
  and _60120_ (_08449_, _08448_, _08432_);
  and _60121_ (_08450_, _08449_, _08426_);
  and _60122_ (_08451_, _07250_, _06366_);
  not _60123_ (_08452_, _08451_);
  nand _60124_ (_08453_, _08452_, _08450_);
  and _60125_ (_08454_, _08453_, _08404_);
  and _60126_ (_08455_, _07954_, \oc8051_golden_model_1.TH0 [2]);
  and _60127_ (_08456_, _07969_, \oc8051_golden_model_1.SCON [2]);
  nor _60128_ (_08457_, _08456_, _08455_);
  and _60129_ (_08458_, _07965_, \oc8051_golden_model_1.TMOD [2]);
  and _60130_ (_08459_, _07981_, \oc8051_golden_model_1.TH1 [2]);
  nor _60131_ (_08460_, _08459_, _08458_);
  and _60132_ (_08461_, _08460_, _08457_);
  and _60133_ (_08462_, _08014_, \oc8051_golden_model_1.PSW [2]);
  and _60134_ (_08463_, _08017_, \oc8051_golden_model_1.ACC [2]);
  nor _60135_ (_08464_, _08463_, _08462_);
  and _60136_ (_08465_, _08022_, \oc8051_golden_model_1.IP [2]);
  and _60137_ (_08466_, _08025_, \oc8051_golden_model_1.B [2]);
  nor _60138_ (_08467_, _08466_, _08465_);
  and _60139_ (_08468_, _08467_, _08464_);
  and _60140_ (_08469_, _07995_, \oc8051_golden_model_1.DPH [2]);
  not _60141_ (_08470_, _08469_);
  and _60142_ (_08471_, _08470_, _08468_);
  and _60143_ (_08472_, _07991_, \oc8051_golden_model_1.TL1 [2]);
  and _60144_ (_08473_, _07976_, \oc8051_golden_model_1.TL0 [2]);
  nor _60145_ (_08474_, _08473_, _08472_);
  and _60146_ (_08475_, _08474_, _08471_);
  and _60147_ (_08476_, _08475_, _08461_);
  and _60148_ (_08477_, _08001_, \oc8051_golden_model_1.DPL [2]);
  not _60149_ (_08478_, _08477_);
  and _60150_ (_08479_, _08004_, \oc8051_golden_model_1.SP [2]);
  and _60151_ (_08480_, _08006_, \oc8051_golden_model_1.TCON [2]);
  nor _60152_ (_08481_, _08480_, _08479_);
  and _60153_ (_08482_, _08481_, _08478_);
  and _60154_ (_08483_, _08042_, \oc8051_golden_model_1.PCON [2]);
  not _60155_ (_08484_, _08483_);
  and _60156_ (_08485_, _07962_, \oc8051_golden_model_1.SBUF [2]);
  and _60157_ (_08486_, _07986_, \oc8051_golden_model_1.IE [2]);
  nor _60158_ (_08487_, _08486_, _08485_);
  and _60159_ (_08488_, _08487_, _08484_);
  and _60160_ (_08489_, _08039_, \oc8051_golden_model_1.P0INREG [2]);
  not _60161_ (_08490_, _08489_);
  and _60162_ (_08491_, _08029_, \oc8051_golden_model_1.P1INREG [2]);
  not _60163_ (_08492_, _08491_);
  and _60164_ (_08493_, _08032_, \oc8051_golden_model_1.P2INREG [2]);
  and _60165_ (_08494_, _08034_, \oc8051_golden_model_1.P3INREG [2]);
  nor _60166_ (_08495_, _08494_, _08493_);
  and _60167_ (_08496_, _08495_, _08492_);
  and _60168_ (_08497_, _08496_, _08490_);
  and _60169_ (_08498_, _08497_, _08488_);
  and _60170_ (_08499_, _08498_, _08482_);
  and _60171_ (_08500_, _08499_, _08476_);
  or _60172_ (_08501_, _07854_, _06238_);
  and _60173_ (_08502_, _08501_, _08500_);
  not _60174_ (_08503_, _08502_);
  and _60175_ (_08504_, _08503_, _08454_);
  and _60176_ (_08505_, _08504_, _08359_);
  and _60177_ (_08506_, _07954_, \oc8051_golden_model_1.TH0 [4]);
  and _60178_ (_08507_, _07981_, \oc8051_golden_model_1.TH1 [4]);
  nor _60179_ (_08508_, _08507_, _08506_);
  and _60180_ (_08509_, _07965_, \oc8051_golden_model_1.TMOD [4]);
  and _60181_ (_08510_, _07969_, \oc8051_golden_model_1.SCON [4]);
  nor _60182_ (_08511_, _08510_, _08509_);
  and _60183_ (_08512_, _08511_, _08508_);
  and _60184_ (_08513_, _08014_, \oc8051_golden_model_1.PSW [4]);
  and _60185_ (_08514_, _08017_, \oc8051_golden_model_1.ACC [4]);
  nor _60186_ (_08515_, _08514_, _08513_);
  and _60187_ (_08516_, _08022_, \oc8051_golden_model_1.IP [4]);
  and _60188_ (_08517_, _08025_, \oc8051_golden_model_1.B [4]);
  nor _60189_ (_08518_, _08517_, _08516_);
  and _60190_ (_08519_, _08518_, _08515_);
  and _60191_ (_08520_, _07976_, \oc8051_golden_model_1.TL0 [4]);
  not _60192_ (_08521_, _08520_);
  and _60193_ (_08522_, _08521_, _08519_);
  and _60194_ (_08523_, _07991_, \oc8051_golden_model_1.TL1 [4]);
  and _60195_ (_08524_, _07995_, \oc8051_golden_model_1.DPH [4]);
  nor _60196_ (_08525_, _08524_, _08523_);
  and _60197_ (_08526_, _08525_, _08522_);
  and _60198_ (_08527_, _08526_, _08512_);
  and _60199_ (_08528_, _08004_, \oc8051_golden_model_1.SP [4]);
  not _60200_ (_08529_, _08528_);
  and _60201_ (_08530_, _08006_, \oc8051_golden_model_1.TCON [4]);
  and _60202_ (_08531_, _08001_, \oc8051_golden_model_1.DPL [4]);
  nor _60203_ (_08532_, _08531_, _08530_);
  and _60204_ (_08533_, _08532_, _08529_);
  and _60205_ (_08534_, _08042_, \oc8051_golden_model_1.PCON [4]);
  not _60206_ (_08535_, _08534_);
  and _60207_ (_08536_, _07962_, \oc8051_golden_model_1.SBUF [4]);
  and _60208_ (_08537_, _07986_, \oc8051_golden_model_1.IE [4]);
  nor _60209_ (_08538_, _08537_, _08536_);
  and _60210_ (_08539_, _08538_, _08535_);
  and _60211_ (_08540_, _08039_, \oc8051_golden_model_1.P0INREG [4]);
  not _60212_ (_08541_, _08540_);
  and _60213_ (_08542_, _08029_, \oc8051_golden_model_1.P1INREG [4]);
  not _60214_ (_08543_, _08542_);
  and _60215_ (_08544_, _08032_, \oc8051_golden_model_1.P2INREG [4]);
  and _60216_ (_08545_, _08034_, \oc8051_golden_model_1.P3INREG [4]);
  nor _60217_ (_08546_, _08545_, _08544_);
  and _60218_ (_08547_, _08546_, _08543_);
  and _60219_ (_08548_, _08547_, _08541_);
  and _60220_ (_08549_, _08548_, _08539_);
  and _60221_ (_08550_, _08549_, _08533_);
  and _60222_ (_08551_, _08550_, _08527_);
  nand _60223_ (_08552_, _07061_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand _60224_ (_08553_, _07199_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _60225_ (_08554_, _08553_, _07198_);
  nand _60226_ (_08555_, _08554_, _08552_);
  nand _60227_ (_08556_, _07199_, \oc8051_golden_model_1.IRAM[3] [4]);
  nand _60228_ (_08557_, _07061_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _60229_ (_08558_, _08557_, _07204_);
  nand _60230_ (_08559_, _08558_, _08556_);
  nand _60231_ (_08560_, _08559_, _08555_);
  nand _60232_ (_08561_, _08560_, _06841_);
  nand _60233_ (_08562_, _07199_, \oc8051_golden_model_1.IRAM[7] [4]);
  nand _60234_ (_08563_, _07061_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _60235_ (_08564_, _08563_, _07204_);
  nand _60236_ (_08565_, _08564_, _08562_);
  nand _60237_ (_08566_, _07061_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand _60238_ (_08567_, _07199_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _60239_ (_08568_, _08567_, _07198_);
  nand _60240_ (_08569_, _08568_, _08566_);
  nand _60241_ (_08570_, _08569_, _08565_);
  nand _60242_ (_08571_, _08570_, _07210_);
  nand _60243_ (_08572_, _08571_, _08561_);
  nand _60244_ (_08573_, _08572_, _06654_);
  nand _60245_ (_08574_, _07199_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _60246_ (_08575_, _07061_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _60247_ (_08576_, _08575_, _07204_);
  nand _60248_ (_08577_, _08576_, _08574_);
  nand _60249_ (_08578_, _07061_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand _60250_ (_08579_, _07199_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _60251_ (_08580_, _08579_, _07198_);
  nand _60252_ (_08581_, _08580_, _08578_);
  nand _60253_ (_08582_, _08581_, _08577_);
  nand _60254_ (_08583_, _08582_, _06841_);
  nand _60255_ (_08584_, _07199_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _60256_ (_08585_, _07061_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _60257_ (_08586_, _08585_, _07204_);
  nand _60258_ (_08587_, _08586_, _08584_);
  nand _60259_ (_08588_, _07061_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand _60260_ (_08589_, _07199_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _60261_ (_08590_, _08589_, _07198_);
  nand _60262_ (_08591_, _08590_, _08588_);
  nand _60263_ (_08592_, _08591_, _08587_);
  nand _60264_ (_08593_, _08592_, _07210_);
  nand _60265_ (_08594_, _08593_, _08583_);
  nand _60266_ (_08595_, _08594_, _07224_);
  nand _60267_ (_08596_, _08595_, _08573_);
  or _60268_ (_08597_, _08596_, _06238_);
  and _60269_ (_08598_, _08597_, _08551_);
  not _60270_ (_08599_, _08598_);
  and _60271_ (_08600_, _08599_, _08505_);
  and _60272_ (_08601_, _08600_, _08308_);
  and _60273_ (_08602_, _08601_, _08212_);
  or _60274_ (_08603_, _08602_, _08110_);
  nand _60275_ (_08604_, _08602_, _08110_);
  and _60276_ (_08605_, _08604_, _08603_);
  and _60277_ (_08606_, _08605_, _07379_);
  and _60278_ (_08607_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _60279_ (_08608_, _08607_, \oc8051_golden_model_1.PC [6]);
  and _60280_ (_08609_, _05705_, \oc8051_golden_model_1.PC [2]);
  and _60281_ (_08610_, _08609_, \oc8051_golden_model_1.PC [3]);
  and _60282_ (_08611_, _08610_, _08608_);
  and _60283_ (_08612_, _08611_, \oc8051_golden_model_1.PC [7]);
  nor _60284_ (_08613_, _08611_, \oc8051_golden_model_1.PC [7]);
  nor _60285_ (_08614_, _08613_, _08612_);
  not _60286_ (_08615_, _08614_);
  nand _60287_ (_08616_, _08615_, _06503_);
  and _60288_ (_08617_, _08608_, _06148_);
  and _60289_ (_08618_, _08617_, \oc8051_golden_model_1.PC [7]);
  nor _60290_ (_08619_, _08617_, \oc8051_golden_model_1.PC [7]);
  nor _60291_ (_08620_, _08619_, _08618_);
  or _60292_ (_08621_, _08620_, _06009_);
  not _60293_ (_08622_, _07557_);
  and _60294_ (_08623_, _06315_, _06276_);
  nor _60295_ (_08624_, _08623_, _07322_);
  and _60296_ (_08625_, _08624_, _07572_);
  and _60297_ (_08626_, _08625_, _08622_);
  and _60298_ (_08627_, _08626_, _06278_);
  or _60299_ (_08628_, _08627_, _06238_);
  not _60300_ (_08629_, _07294_);
  nor _60301_ (_08630_, _07094_, _06686_);
  and _60302_ (_08631_, _08630_, _06270_);
  and _60303_ (_08632_, _08631_, _06399_);
  and _60304_ (_08633_, _08632_, _07948_);
  and _60305_ (_08634_, _08633_, \oc8051_golden_model_1.TCON [7]);
  not _60306_ (_08635_, _06399_);
  and _60307_ (_08636_, _08631_, _08635_);
  and _60308_ (_08637_, _08024_, _08636_);
  and _60309_ (_08638_, _08637_, \oc8051_golden_model_1.B [7]);
  nor _60310_ (_08639_, _08638_, _08634_);
  and _60311_ (_08640_, _08013_, _08636_);
  and _60312_ (_08641_, _08640_, \oc8051_golden_model_1.PSW [7]);
  not _60313_ (_08642_, _08641_);
  and _60314_ (_08643_, _08632_, _08021_);
  and _60315_ (_08644_, _08643_, \oc8051_golden_model_1.IP [7]);
  and _60316_ (_08645_, _08016_, _08636_);
  and _60317_ (_08646_, _08645_, \oc8051_golden_model_1.ACC [7]);
  nor _60318_ (_08647_, _08646_, _08644_);
  and _60319_ (_08648_, _08647_, _08642_);
  and _60320_ (_08649_, _08648_, _08639_);
  and _60321_ (_08650_, _08632_, _07961_);
  and _60322_ (_08651_, _08650_, \oc8051_golden_model_1.SCON [7]);
  and _60323_ (_08652_, _08632_, _07985_);
  and _60324_ (_08653_, _08652_, \oc8051_golden_model_1.IE [7]);
  nor _60325_ (_08654_, _08653_, _08651_);
  and _60326_ (_08655_, _08636_, _07985_);
  and _60327_ (_08656_, _08655_, \oc8051_golden_model_1.P2INREG [7]);
  and _60328_ (_08657_, _08021_, _08636_);
  and _60329_ (_08658_, _08657_, \oc8051_golden_model_1.P3INREG [7]);
  nor _60330_ (_08659_, _08658_, _08656_);
  and _60331_ (_08660_, _07993_, \oc8051_golden_model_1.P0INREG [7]);
  and _60332_ (_08661_, _08636_, _07961_);
  and _60333_ (_08662_, _08661_, \oc8051_golden_model_1.P1INREG [7]);
  nor _60334_ (_08663_, _08662_, _08660_);
  and _60335_ (_08664_, _08663_, _08659_);
  and _60336_ (_08665_, _08664_, _08654_);
  and _60337_ (_08666_, _08665_, _08649_);
  and _60338_ (_08667_, _08666_, _08108_);
  nor _60339_ (_08668_, _08667_, _08041_);
  or _60340_ (_08669_, _08668_, _08629_);
  not _60341_ (_08670_, _07274_);
  not _60342_ (_08671_, _08041_);
  nand _60343_ (_08672_, _08667_, _08671_);
  or _60344_ (_08673_, _08672_, _08670_);
  not _60345_ (_08674_, _08107_);
  and _60346_ (_08675_, _08596_, _08305_);
  and _60347_ (_08676_, _07854_, _07680_);
  and _60348_ (_08677_, _07448_, _07321_);
  and _60349_ (_08678_, _08677_, _08676_);
  and _60350_ (_08679_, _08678_, _08675_);
  and _60351_ (_08680_, _08679_, _08209_);
  or _60352_ (_08681_, _08680_, _08674_);
  nand _60353_ (_08682_, _08680_, _08674_);
  and _60354_ (_08683_, _08682_, _08681_);
  nor _60355_ (_08684_, _06319_, _06051_);
  nor _60356_ (_08685_, _07860_, _08684_);
  or _60357_ (_08686_, _08685_, _08683_);
  not _60358_ (_08687_, _08685_);
  not _60359_ (_08688_, \oc8051_golden_model_1.ACC [7]);
  nor _60360_ (_08689_, _06816_, _08688_);
  and _60361_ (_08690_, _08620_, _06816_);
  or _60362_ (_08691_, _08690_, _08689_);
  or _60363_ (_08692_, _08691_, _08687_);
  and _60364_ (_08693_, _08692_, _08686_);
  or _60365_ (_08694_, _08693_, _07269_);
  nor _60366_ (_08695_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _60367_ (_08696_, _08695_, _06771_);
  nor _60368_ (_08697_, _08696_, _06409_);
  nor _60369_ (_08698_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _60370_ (_08699_, _08698_, _06409_);
  and _60371_ (_08700_, _08699_, _06342_);
  nor _60372_ (_08701_, _08700_, _08697_);
  nor _60373_ (_08702_, _08701_, _06773_);
  and _60374_ (_08703_, _07680_, _07310_);
  not _60375_ (_08704_, _06773_);
  and _60376_ (_08705_, _07309_, _06269_);
  or _60377_ (_08706_, _08705_, _08704_);
  nor _60378_ (_08707_, _08706_, _08703_);
  nor _60379_ (_08708_, _08707_, _08702_);
  not _60380_ (_08709_, _08708_);
  nor _60381_ (_08710_, _07854_, _07309_);
  nor _60382_ (_08711_, _07310_, _06727_);
  nor _60383_ (_08712_, _08711_, _08704_);
  not _60384_ (_08713_, _08712_);
  nor _60385_ (_08714_, _08713_, _08710_);
  nor _60386_ (_08715_, _08695_, _06771_);
  nor _60387_ (_08716_, _08715_, _08696_);
  and _60388_ (_08717_, _08716_, _08704_);
  nor _60389_ (_08718_, _08717_, _08714_);
  not _60390_ (_08719_, _08718_);
  or _60391_ (_08720_, _07309_, _07250_);
  and _60392_ (_08721_, _07309_, _06310_);
  nor _60393_ (_08722_, _08721_, _08704_);
  nand _60394_ (_08723_, _08722_, _08720_);
  nor _60395_ (_08724_, _06773_, \oc8051_golden_model_1.SP [0]);
  not _60396_ (_08725_, _08724_);
  and _60397_ (_08726_, _08725_, _08723_);
  or _60398_ (_08727_, _08726_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor _60399_ (_08728_, _07310_, _07127_);
  nor _60400_ (_08729_, _07448_, _07309_);
  or _60401_ (_08730_, _08729_, _08728_);
  nand _60402_ (_08731_, _08730_, _06773_);
  nor _60403_ (_08732_, _07392_, _06773_);
  not _60404_ (_08733_, _08732_);
  and _60405_ (_08734_, _08733_, _08731_);
  nand _60406_ (_08735_, _08726_, _08084_);
  and _60407_ (_08736_, _08735_, _08734_);
  nand _60408_ (_08737_, _08736_, _08727_);
  nand _60409_ (_08738_, _08726_, _08080_);
  nor _60410_ (_08739_, _08726_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor _60411_ (_08740_, _08739_, _08734_);
  nand _60412_ (_08741_, _08740_, _08738_);
  nand _60413_ (_08742_, _08741_, _08737_);
  and _60414_ (_08743_, _08742_, _08719_);
  or _60415_ (_08744_, _08726_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand _60416_ (_08745_, _08726_, _08097_);
  and _60417_ (_08746_, _08745_, _08734_);
  nand _60418_ (_08747_, _08746_, _08744_);
  nand _60419_ (_08748_, _08726_, _08093_);
  nor _60420_ (_08749_, _08726_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor _60421_ (_08750_, _08749_, _08734_);
  nand _60422_ (_08751_, _08750_, _08748_);
  nand _60423_ (_08752_, _08751_, _08747_);
  and _60424_ (_08753_, _08752_, _08718_);
  nor _60425_ (_08754_, _08753_, _08743_);
  nand _60426_ (_08755_, _08754_, _08709_);
  nand _60427_ (_08756_, _08726_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor _60428_ (_08757_, _08726_, _08062_);
  nor _60429_ (_08758_, _08757_, _08734_);
  nand _60430_ (_08759_, _08758_, _08756_);
  nand _60431_ (_08760_, _08726_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _60432_ (_08761_, _08726_, _08070_);
  and _60433_ (_08762_, _08761_, _08734_);
  nand _60434_ (_08763_, _08762_, _08760_);
  nand _60435_ (_08764_, _08763_, _08759_);
  nand _60436_ (_08765_, _08764_, _08718_);
  nand _60437_ (_08766_, _08726_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _60438_ (_08767_, _08726_, _08054_);
  nor _60439_ (_08768_, _08767_, _08734_);
  nand _60440_ (_08769_, _08768_, _08766_);
  nand _60441_ (_08770_, _08726_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _60442_ (_08771_, _08726_, _08050_);
  and _60443_ (_08772_, _08771_, _08734_);
  nand _60444_ (_08773_, _08772_, _08770_);
  nand _60445_ (_08774_, _08773_, _08769_);
  nand _60446_ (_08775_, _08774_, _08719_);
  nand _60447_ (_08776_, _08775_, _08765_);
  nand _60448_ (_08777_, _08776_, _08708_);
  and _60449_ (_08778_, _08777_, _08755_);
  or _60450_ (_08779_, _08778_, _07270_);
  and _60451_ (_08780_, _08779_, _08694_);
  or _60452_ (_08781_, _08780_, _07276_);
  not _60453_ (_08782_, _07276_);
  and _60454_ (_08783_, _08598_, _08307_);
  nor _60455_ (_08784_, _08453_, _08404_);
  and _60456_ (_08785_, _08502_, _08358_);
  and _60457_ (_08786_, _08785_, _08784_);
  and _60458_ (_08787_, _08786_, _08783_);
  and _60459_ (_08788_, _08787_, _08211_);
  or _60460_ (_08789_, _08788_, _08110_);
  nand _60461_ (_08790_, _08788_, _08110_);
  and _60462_ (_08791_, _08790_, _08789_);
  or _60463_ (_08792_, _08791_, _08782_);
  and _60464_ (_08793_, _08792_, _08781_);
  or _60465_ (_08794_, _08793_, _07274_);
  and _60466_ (_08795_, _08794_, _08673_);
  or _60467_ (_08796_, _08795_, _07692_);
  nor _60468_ (_08797_, _08620_, _06052_);
  nor _60469_ (_08798_, _08797_, _07284_);
  and _60470_ (_08799_, _08798_, _08796_);
  and _60471_ (_08800_, _08674_, _07284_);
  or _60472_ (_08801_, _08800_, _07294_);
  or _60473_ (_08802_, _08801_, _08799_);
  and _60474_ (_08803_, _08802_, _08669_);
  or _60475_ (_08804_, _08803_, _06351_);
  nand _60476_ (_08805_, _08109_, _06351_);
  and _60477_ (_08806_, _08805_, _06349_);
  and _60478_ (_08807_, _08806_, _08804_);
  nor _60479_ (_08808_, _08667_, _08671_);
  not _60480_ (_08809_, _08808_);
  and _60481_ (_08810_, _08809_, _08672_);
  and _60482_ (_08811_, _08810_, _06348_);
  or _60483_ (_08812_, _08811_, _08807_);
  and _60484_ (_08813_, _08812_, _06049_);
  not _60485_ (_08814_, _08620_);
  nor _60486_ (_08815_, _08814_, _06049_);
  or _60487_ (_08816_, _08815_, _06441_);
  or _60488_ (_08817_, _08816_, _08813_);
  nand _60489_ (_08818_, _08109_, _06441_);
  and _60490_ (_08819_, _08818_, _08817_);
  or _60491_ (_08820_, _08819_, _07309_);
  not _60492_ (_08821_, _07308_);
  nand _60493_ (_08822_, _08778_, _06366_);
  and _60494_ (_08823_, _08047_, _07309_);
  nand _60495_ (_08824_, _08823_, _08822_);
  and _60496_ (_08825_, _08824_, _08821_);
  and _60497_ (_08826_, _08825_, _08820_);
  and _60498_ (_08827_, _08041_, \oc8051_golden_model_1.PSW [7]);
  or _60499_ (_08828_, _08827_, _08668_);
  and _60500_ (_08829_, _08828_, _07308_);
  or _60501_ (_08830_, _08829_, _06039_);
  or _60502_ (_08831_, _08830_, _08826_);
  nor _60503_ (_08832_, _06327_, _06238_);
  and _60504_ (_08833_, _08814_, _06039_);
  nor _60505_ (_08834_, _08833_, _08832_);
  and _60506_ (_08835_, _08834_, _08831_);
  not _60507_ (_08836_, _08832_);
  nor _60508_ (_08837_, _08836_, _08107_);
  nor _60509_ (_08838_, _06333_, _06238_);
  or _60510_ (_08839_, _08838_, _08837_);
  or _60511_ (_08840_, _08839_, _08835_);
  nor _60512_ (_08841_, _06238_, _06313_);
  not _60513_ (_08842_, _08841_);
  not _60514_ (_08843_, _06471_);
  or _60515_ (_08844_, _07544_, _08843_);
  or _60516_ (_08845_, _08844_, _08778_);
  and _60517_ (_08846_, _08845_, _08842_);
  and _60518_ (_08847_, _08846_, _08840_);
  not _60519_ (_08848_, _08626_);
  and _60520_ (_08849_, _06541_, _04443_);
  and _60521_ (_08850_, _06565_, _04458_);
  nor _60522_ (_08851_, _08850_, _08849_);
  and _60523_ (_08852_, _06579_, _04481_);
  and _60524_ (_08853_, _06560_, _04453_);
  nor _60525_ (_08854_, _08853_, _08852_);
  and _60526_ (_08855_, _08854_, _08851_);
  and _60527_ (_08856_, _06551_, _04500_);
  and _60528_ (_08857_, _06574_, _04502_);
  nor _60529_ (_08858_, _08857_, _08856_);
  and _60530_ (_08859_, _06572_, _04479_);
  and _60531_ (_08860_, _06554_, _04492_);
  nor _60532_ (_08861_, _08860_, _08859_);
  and _60533_ (_08862_, _08861_, _08858_);
  and _60534_ (_08863_, _08862_, _08855_);
  and _60535_ (_08864_, _06546_, _04489_);
  and _60536_ (_08865_, _06567_, _04470_);
  nor _60537_ (_08866_, _08865_, _08864_);
  and _60538_ (_08867_, _06585_, _04486_);
  and _60539_ (_08868_, _06588_, _04475_);
  nor _60540_ (_08869_, _08868_, _08867_);
  and _60541_ (_08870_, _08869_, _08866_);
  and _60542_ (_08871_, _06583_, _04463_);
  and _60543_ (_08872_, _06577_, _04467_);
  nor _60544_ (_08873_, _08872_, _08871_);
  and _60545_ (_08874_, _06590_, _04495_);
  and _60546_ (_08875_, _06562_, _04414_);
  nor _60547_ (_08876_, _08875_, _08874_);
  and _60548_ (_08877_, _08876_, _08873_);
  and _60549_ (_08878_, _08877_, _08870_);
  and _60550_ (_08879_, _08878_, _08863_);
  not _60551_ (_08880_, _08879_);
  nor _60552_ (_08881_, _08880_, _08107_);
  and _60553_ (_08882_, _07160_, _06950_);
  and _60554_ (_08883_, _06769_, _06595_);
  and _60555_ (_08884_, _08883_, _08882_);
  and _60556_ (_08885_, _06541_, _04898_);
  and _60557_ (_08886_, _06560_, _04881_);
  nor _60558_ (_08887_, _08886_, _08885_);
  and _60559_ (_08888_, _06565_, _04887_);
  and _60560_ (_08890_, _06590_, _04909_);
  nor _60561_ (_08891_, _08890_, _08888_);
  and _60562_ (_08892_, _08891_, _08887_);
  and _60563_ (_08893_, _06577_, _04904_);
  and _60564_ (_08894_, _06562_, _04915_);
  nor _60565_ (_08895_, _08894_, _08893_);
  and _60566_ (_08896_, _06579_, _04911_);
  and _60567_ (_08897_, _06546_, _04877_);
  nor _60568_ (_08898_, _08897_, _08896_);
  and _60569_ (_08899_, _08898_, _08895_);
  and _60570_ (_08901_, _08899_, _08892_);
  and _60571_ (_08902_, _06588_, _04892_);
  and _60572_ (_08903_, _06567_, _04879_);
  nor _60573_ (_08904_, _08903_, _08902_);
  and _60574_ (_08905_, _06572_, _04890_);
  and _60575_ (_08906_, _06583_, _04913_);
  nor _60576_ (_08907_, _08906_, _08905_);
  and _60577_ (_08908_, _08907_, _08904_);
  and _60578_ (_08909_, _06551_, _04900_);
  and _60579_ (_08910_, _06554_, _04906_);
  nor _60580_ (_08912_, _08910_, _08909_);
  and _60581_ (_08913_, _06574_, _04885_);
  and _60582_ (_08914_, _06585_, _04896_);
  nor _60583_ (_08915_, _08914_, _08913_);
  and _60584_ (_08916_, _08915_, _08912_);
  and _60585_ (_08917_, _08916_, _08908_);
  and _60586_ (_08918_, _08917_, _08901_);
  and _60587_ (_08919_, _08918_, _08880_);
  and _60588_ (_08920_, _06588_, _04846_);
  and _60589_ (_08921_, _06567_, _04831_);
  nor _60590_ (_08923_, _08921_, _08920_);
  and _60591_ (_08924_, _06574_, _04841_);
  and _60592_ (_08925_, _06554_, _04852_);
  nor _60593_ (_08926_, _08925_, _08924_);
  and _60594_ (_08927_, _08926_, _08923_);
  and _60595_ (_08928_, _06562_, _04864_);
  and _60596_ (_08929_, _06560_, _04835_);
  nor _60597_ (_08930_, _08929_, _08928_);
  and _60598_ (_08931_, _06579_, _04860_);
  and _60599_ (_08932_, _06546_, _04833_);
  nor _60600_ (_08934_, _08932_, _08931_);
  and _60601_ (_08935_, _08934_, _08930_);
  and _60602_ (_08936_, _08935_, _08927_);
  and _60603_ (_08937_, _06541_, _04858_);
  and _60604_ (_08938_, _06551_, _04869_);
  nor _60605_ (_08939_, _08938_, _08937_);
  and _60606_ (_08940_, _06572_, _04839_);
  and _60607_ (_08941_, _06565_, _04844_);
  nor _60608_ (_08942_, _08941_, _08940_);
  and _60609_ (_08943_, _08942_, _08939_);
  and _60610_ (_08945_, _06583_, _04862_);
  and _60611_ (_08946_, _06577_, _04871_);
  nor _60612_ (_08947_, _08946_, _08945_);
  and _60613_ (_08948_, _06585_, _04850_);
  and _60614_ (_08949_, _06590_, _04855_);
  nor _60615_ (_08950_, _08949_, _08948_);
  and _60616_ (_08951_, _08950_, _08947_);
  and _60617_ (_08952_, _08951_, _08943_);
  and _60618_ (_08953_, _08952_, _08936_);
  not _60619_ (_08954_, _08953_);
  and _60620_ (_08956_, _06585_, _04804_);
  and _60621_ (_08957_, _06560_, _04789_);
  nor _60622_ (_08958_, _08957_, _08956_);
  and _60623_ (_08959_, _06551_, _04823_);
  and _60624_ (_08960_, _06567_, _04785_);
  nor _60625_ (_08961_, _08960_, _08959_);
  and _60626_ (_08962_, _08961_, _08958_);
  and _60627_ (_08963_, _06572_, _04793_);
  and _60628_ (_08964_, _06574_, _04795_);
  nor _60629_ (_08965_, _08964_, _08963_);
  and _60630_ (_08966_, _06588_, _04800_);
  and _60631_ (_08967_, _06546_, _04787_);
  nor _60632_ (_08968_, _08967_, _08966_);
  and _60633_ (_08969_, _08968_, _08965_);
  and _60634_ (_08970_, _08969_, _08962_);
  and _60635_ (_08971_, _06583_, _04816_);
  and _60636_ (_08972_, _06554_, _04806_);
  nor _60637_ (_08973_, _08972_, _08971_);
  and _60638_ (_08974_, _06590_, _04809_);
  and _60639_ (_08975_, _06562_, _04818_);
  nor _60640_ (_08976_, _08975_, _08974_);
  and _60641_ (_08977_, _08976_, _08973_);
  and _60642_ (_08978_, _06541_, _04812_);
  and _60643_ (_08979_, _06579_, _04814_);
  nor _60644_ (_08980_, _08979_, _08978_);
  and _60645_ (_08981_, _06565_, _04798_);
  and _60646_ (_08982_, _06577_, _04825_);
  nor _60647_ (_08983_, _08982_, _08981_);
  and _60648_ (_08984_, _08983_, _08980_);
  and _60649_ (_08985_, _08984_, _08977_);
  and _60650_ (_08986_, _08985_, _08970_);
  and _60651_ (_08987_, _08986_, _08954_);
  and _60652_ (_08988_, _08987_, _08919_);
  and _60653_ (_08989_, _08988_, _08884_);
  and _60654_ (_08990_, _08989_, \oc8051_golden_model_1.P2INREG [7]);
  and _60655_ (_08991_, _08986_, _08953_);
  and _60656_ (_08992_, _08991_, _08919_);
  and _60657_ (_08993_, _08992_, _08884_);
  and _60658_ (_08994_, _08993_, \oc8051_golden_model_1.P0INREG [7]);
  not _60659_ (_08995_, _08986_);
  and _60660_ (_08996_, _08995_, _08953_);
  and _60661_ (_08997_, _08996_, _08919_);
  and _60662_ (_08998_, _08997_, _08884_);
  and _60663_ (_08999_, _08998_, \oc8051_golden_model_1.P1INREG [7]);
  nor _60664_ (_09000_, _08986_, _08953_);
  and _60665_ (_09001_, _09000_, _08919_);
  and _60666_ (_09002_, _09001_, _08884_);
  and _60667_ (_09003_, _09002_, \oc8051_golden_model_1.P3INREG [7]);
  or _60668_ (_09004_, _09003_, _08999_);
  or _60669_ (_09005_, _09004_, _08994_);
  or _60670_ (_09006_, _09005_, _08990_);
  and _60671_ (_09007_, _08992_, _08883_);
  not _60672_ (_09008_, _06950_);
  and _60673_ (_09009_, _07160_, _09008_);
  and _60674_ (_09010_, _09009_, _09007_);
  and _60675_ (_09011_, _09010_, \oc8051_golden_model_1.SP [7]);
  not _60676_ (_09012_, _07160_);
  and _60677_ (_09013_, _09012_, _06950_);
  not _60678_ (_09014_, _06595_);
  and _60679_ (_09015_, _06769_, _09014_);
  and _60680_ (_09016_, _09015_, _08992_);
  and _60681_ (_09017_, _09016_, _09013_);
  and _60682_ (_09018_, _09017_, \oc8051_golden_model_1.TL0 [7]);
  or _60683_ (_09019_, _09018_, _09011_);
  or _60684_ (_09020_, _09019_, _09006_);
  nor _60685_ (_09021_, _08918_, _08879_);
  and _60686_ (_09022_, _09021_, _08884_);
  and _60687_ (_09023_, _09022_, _08996_);
  and _60688_ (_09024_, _09023_, \oc8051_golden_model_1.PSW [7]);
  and _60689_ (_09025_, _09015_, _08882_);
  and _60690_ (_09026_, _09025_, _09001_);
  and _60691_ (_09027_, _09026_, \oc8051_golden_model_1.IP [7]);
  and _60692_ (_09028_, _09022_, _08987_);
  and _60693_ (_09029_, _09028_, \oc8051_golden_model_1.ACC [7]);
  and _60694_ (_09030_, _09022_, _09000_);
  and _60695_ (_09031_, _09030_, \oc8051_golden_model_1.B [7]);
  or _60696_ (_09032_, _09031_, _09029_);
  or _60697_ (_09033_, _09032_, _09027_);
  or _60698_ (_09034_, _09033_, _09024_);
  and _60699_ (_09035_, _09025_, _08997_);
  and _60700_ (_09036_, _09035_, \oc8051_golden_model_1.SCON [7]);
  and _60701_ (_09037_, _09015_, _09009_);
  and _60702_ (_09038_, _09037_, _08997_);
  and _60703_ (_09039_, _09038_, \oc8051_golden_model_1.SBUF [7]);
  or _60704_ (_09040_, _09039_, _09036_);
  and _60705_ (_09041_, _09025_, _08988_);
  and _60706_ (_09042_, _09041_, \oc8051_golden_model_1.IE [7]);
  or _60707_ (_09043_, _09042_, _09040_);
  or _60708_ (_09044_, _09043_, _09034_);
  or _60709_ (_09045_, _09044_, _09020_);
  nor _60710_ (_09046_, _06769_, _06595_);
  and _60711_ (_09047_, _09046_, _08992_);
  and _60712_ (_09048_, _09047_, _08882_);
  and _60713_ (_09049_, _09048_, \oc8051_golden_model_1.TH0 [7]);
  nor _60714_ (_09050_, _07160_, _06950_);
  and _60715_ (_09051_, _09050_, _08992_);
  and _60716_ (_09052_, _09051_, _09015_);
  and _60717_ (_09053_, _09052_, \oc8051_golden_model_1.TL1 [7]);
  or _60718_ (_09054_, _09053_, _09049_);
  and _60719_ (_09055_, _09025_, _08992_);
  and _60720_ (_09056_, _09055_, \oc8051_golden_model_1.TCON [7]);
  not _60721_ (_09057_, _06769_);
  and _60722_ (_09058_, _09057_, _06595_);
  and _60723_ (_09059_, _09051_, _09058_);
  and _60724_ (_09060_, _09059_, \oc8051_golden_model_1.PCON [7]);
  or _60725_ (_09061_, _09060_, _09056_);
  or _60726_ (_09062_, _09061_, _09054_);
  and _60727_ (_09063_, _09037_, _08992_);
  and _60728_ (_09064_, _09063_, \oc8051_golden_model_1.TMOD [7]);
  and _60729_ (_09065_, _09051_, _08883_);
  and _60730_ (_09066_, _09065_, \oc8051_golden_model_1.DPH [7]);
  or _60731_ (_09067_, _09066_, _09064_);
  and _60732_ (_09068_, _09013_, _09007_);
  and _60733_ (_09069_, _09068_, \oc8051_golden_model_1.DPL [7]);
  and _60734_ (_09070_, _09047_, _09009_);
  and _60735_ (_09071_, _09070_, \oc8051_golden_model_1.TH1 [7]);
  or _60736_ (_09072_, _09071_, _09069_);
  or _60737_ (_09073_, _09072_, _09067_);
  or _60738_ (_09074_, _09073_, _09062_);
  or _60739_ (_09075_, _09074_, _09045_);
  or _60740_ (_09076_, _09075_, _08881_);
  and _60741_ (_09077_, _09076_, _08841_);
  or _60742_ (_09078_, _09077_, _08848_);
  or _60743_ (_09079_, _09078_, _08847_);
  and _60744_ (_09080_, _09079_, _08628_);
  and _60745_ (_09081_, _08880_, _06279_);
  or _60746_ (_09082_, _09081_, _06275_);
  or _60747_ (_09083_, _09082_, _09080_);
  and _60748_ (_09084_, _09083_, _08621_);
  or _60749_ (_09085_, _09084_, _07335_);
  not _60750_ (_09086_, _07338_);
  nand _60751_ (_09087_, _08879_, _08109_);
  nor _60752_ (_09088_, _08879_, _08109_);
  not _60753_ (_09089_, _09088_);
  and _60754_ (_09090_, _09089_, _09087_);
  or _60755_ (_09091_, _09090_, _07336_);
  and _60756_ (_09092_, _09091_, _09086_);
  and _60757_ (_09093_, _09092_, _09085_);
  nor _60758_ (_09094_, _08109_, _08688_);
  and _60759_ (_09095_, _08109_, _08688_);
  nor _60760_ (_09096_, _09095_, _09094_);
  nor _60761_ (_09097_, _09096_, _07340_);
  nor _60762_ (_09098_, _09097_, _07341_);
  or _60763_ (_09099_, _09098_, _09093_);
  not _60764_ (_09100_, _07340_);
  or _60765_ (_09101_, _09088_, _09100_);
  and _60766_ (_09102_, _09101_, _07333_);
  and _60767_ (_09103_, _09102_, _09099_);
  and _60768_ (_09104_, _09094_, _07332_);
  or _60769_ (_09105_, _09104_, _07330_);
  or _60770_ (_09106_, _09105_, _09103_);
  not _60771_ (_09107_, _06509_);
  nor _60772_ (_09108_, _09107_, _06238_);
  nor _60773_ (_09109_, _08620_, _06018_);
  nor _60774_ (_09110_, _09109_, _09108_);
  and _60775_ (_09111_, _09110_, _09106_);
  not _60776_ (_09112_, _06602_);
  nor _60777_ (_09113_, _09112_, _06238_);
  and _60778_ (_09114_, _09087_, _09108_);
  or _60779_ (_09115_, _09114_, _09113_);
  or _60780_ (_09116_, _09115_, _09111_);
  nand _60781_ (_09117_, _09095_, _09113_);
  and _60782_ (_09118_, _09117_, _06016_);
  and _60783_ (_09119_, _09118_, _09116_);
  or _60784_ (_09120_, _08814_, _06016_);
  not _60785_ (_09121_, _07561_);
  nor _60786_ (_09122_, _07177_, _07588_);
  and _60787_ (_09123_, _09122_, _09121_);
  nand _60788_ (_09124_, _09123_, _09120_);
  or _60789_ (_09125_, _09124_, _09119_);
  not _60790_ (_09126_, _08726_);
  or _60791_ (_09127_, _09126_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _60792_ (_09128_, _08726_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _60793_ (_09129_, _09128_, _09127_);
  nand _60794_ (_09130_, _09129_, _08734_);
  not _60795_ (_09131_, _08734_);
  or _60796_ (_09132_, _09126_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _60797_ (_09133_, _08726_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _60798_ (_09134_, _09133_, _09132_);
  nand _60799_ (_09135_, _09134_, _09131_);
  nand _60800_ (_09136_, _09135_, _09130_);
  nand _60801_ (_09137_, _09136_, _08718_);
  or _60802_ (_09138_, _09126_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _60803_ (_09139_, _08726_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _60804_ (_09140_, _09139_, _09138_);
  nand _60805_ (_09141_, _09140_, _08734_);
  or _60806_ (_09142_, _09126_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _60807_ (_09143_, _08726_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _60808_ (_09144_, _09143_, _09142_);
  nand _60809_ (_09145_, _09144_, _09131_);
  nand _60810_ (_09146_, _09145_, _09141_);
  nand _60811_ (_09147_, _09146_, _08719_);
  nand _60812_ (_09148_, _09147_, _09137_);
  nand _60813_ (_09149_, _09148_, _08709_);
  nand _60814_ (_09150_, _08719_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _60815_ (_09151_, _08718_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor _60816_ (_09152_, _09151_, _08734_);
  and _60817_ (_09153_, _09152_, _09150_);
  nand _60818_ (_09154_, _08719_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand _60819_ (_09155_, _08718_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _60820_ (_09156_, _09155_, _08734_);
  and _60821_ (_09157_, _09156_, _09154_);
  or _60822_ (_09158_, _09157_, _09153_);
  and _60823_ (_09159_, _09158_, _08726_);
  nand _60824_ (_09160_, _08719_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _60825_ (_09161_, _08718_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor _60826_ (_09162_, _09161_, _08734_);
  and _60827_ (_09163_, _09162_, _09160_);
  nand _60828_ (_09164_, _08719_, \oc8051_golden_model_1.IRAM[1] [6]);
  nand _60829_ (_09165_, _08718_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _60830_ (_09166_, _09165_, _08734_);
  and _60831_ (_09167_, _09166_, _09164_);
  or _60832_ (_09168_, _09167_, _09163_);
  and _60833_ (_09169_, _09168_, _09126_);
  or _60834_ (_09170_, _09169_, _09159_);
  nand _60835_ (_09171_, _09170_, _08708_);
  and _60836_ (_09172_, _09171_, _09149_);
  not _60837_ (_09173_, _09172_);
  or _60838_ (_09174_, _09126_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _60839_ (_09175_, _08726_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _60840_ (_09176_, _09175_, _09174_);
  nand _60841_ (_09177_, _09176_, _08734_);
  or _60842_ (_09178_, _09126_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _60843_ (_09179_, _08726_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _60844_ (_09180_, _09179_, _09178_);
  nand _60845_ (_09181_, _09180_, _09131_);
  nand _60846_ (_09182_, _09181_, _09177_);
  nand _60847_ (_09183_, _09182_, _08718_);
  or _60848_ (_09184_, _09126_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _60849_ (_09185_, _08726_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _60850_ (_09186_, _09185_, _09184_);
  nand _60851_ (_09187_, _09186_, _08734_);
  or _60852_ (_09188_, _09126_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _60853_ (_09189_, _08726_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _60854_ (_09190_, _09189_, _09188_);
  nand _60855_ (_09191_, _09190_, _09131_);
  nand _60856_ (_09192_, _09191_, _09187_);
  nand _60857_ (_09193_, _09192_, _08719_);
  nand _60858_ (_09194_, _09193_, _09183_);
  nand _60859_ (_09195_, _09194_, _08709_);
  nand _60860_ (_09196_, _08719_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _60861_ (_09197_, _08718_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor _60862_ (_09198_, _09197_, _08734_);
  and _60863_ (_09199_, _09198_, _09196_);
  nand _60864_ (_09200_, _08719_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand _60865_ (_09201_, _08718_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _60866_ (_09202_, _09201_, _08734_);
  and _60867_ (_09203_, _09202_, _09200_);
  or _60868_ (_09204_, _09203_, _09199_);
  and _60869_ (_09205_, _09204_, _08726_);
  nand _60870_ (_09206_, _08719_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _60871_ (_09207_, _08718_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor _60872_ (_09208_, _09207_, _08734_);
  and _60873_ (_09209_, _09208_, _09206_);
  nand _60874_ (_09210_, _08719_, \oc8051_golden_model_1.IRAM[1] [5]);
  nand _60875_ (_09211_, _08718_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _60876_ (_09212_, _09211_, _08734_);
  and _60877_ (_09213_, _09212_, _09210_);
  or _60878_ (_09214_, _09213_, _09209_);
  and _60879_ (_09215_, _09214_, _09126_);
  or _60880_ (_09216_, _09215_, _09205_);
  nand _60881_ (_09217_, _09216_, _08708_);
  and _60882_ (_09218_, _09217_, _09195_);
  not _60883_ (_09219_, _09218_);
  or _60884_ (_09220_, _09126_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _60885_ (_09221_, _08726_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _60886_ (_09222_, _09221_, _09220_);
  nand _60887_ (_09223_, _09222_, _08734_);
  or _60888_ (_09224_, _09126_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _60889_ (_09225_, _08726_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _60890_ (_09226_, _09225_, _09224_);
  nand _60891_ (_09227_, _09226_, _09131_);
  nand _60892_ (_09228_, _09227_, _09223_);
  nand _60893_ (_09229_, _09228_, _08718_);
  or _60894_ (_09230_, _09126_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _60895_ (_09231_, _08726_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _60896_ (_09232_, _09231_, _09230_);
  nand _60897_ (_09233_, _09232_, _08734_);
  or _60898_ (_09234_, _09126_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _60899_ (_09235_, _08726_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _60900_ (_09236_, _09235_, _09234_);
  nand _60901_ (_09237_, _09236_, _09131_);
  nand _60902_ (_09238_, _09237_, _09233_);
  nand _60903_ (_09239_, _09238_, _08719_);
  nand _60904_ (_09240_, _09239_, _09229_);
  nand _60905_ (_09241_, _09240_, _08709_);
  nand _60906_ (_09242_, _08719_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _60907_ (_09243_, _08718_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor _60908_ (_09244_, _09243_, _08734_);
  and _60909_ (_09245_, _09244_, _09242_);
  nand _60910_ (_09246_, _08719_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand _60911_ (_09247_, _08718_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _60912_ (_09248_, _09247_, _08734_);
  and _60913_ (_09249_, _09248_, _09246_);
  or _60914_ (_09250_, _09249_, _09245_);
  and _60915_ (_09251_, _09250_, _08726_);
  nand _60916_ (_09252_, _08719_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _60917_ (_09253_, _08718_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor _60918_ (_09254_, _09253_, _08734_);
  and _60919_ (_09255_, _09254_, _09252_);
  nand _60920_ (_09256_, _08719_, \oc8051_golden_model_1.IRAM[1] [4]);
  nand _60921_ (_09257_, _08718_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _60922_ (_09258_, _09257_, _08734_);
  and _60923_ (_09259_, _09258_, _09256_);
  or _60924_ (_09260_, _09259_, _09255_);
  and _60925_ (_09261_, _09260_, _09126_);
  or _60926_ (_09262_, _09261_, _09251_);
  nand _60927_ (_09263_, _09262_, _08708_);
  and _60928_ (_09264_, _09263_, _09241_);
  not _60929_ (_09265_, _09264_);
  or _60930_ (_09266_, _09126_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _60931_ (_09267_, _08726_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _60932_ (_09268_, _09267_, _09266_);
  nand _60933_ (_09269_, _09268_, _08734_);
  or _60934_ (_09270_, _09126_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _60935_ (_09271_, _08726_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _60936_ (_09272_, _09271_, _09270_);
  nand _60937_ (_09273_, _09272_, _09131_);
  nand _60938_ (_09274_, _09273_, _09269_);
  nand _60939_ (_09275_, _09274_, _08718_);
  or _60940_ (_09276_, _09126_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _60941_ (_09277_, _08726_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _60942_ (_09278_, _09277_, _09276_);
  nand _60943_ (_09279_, _09278_, _08734_);
  or _60944_ (_09280_, _09126_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _60945_ (_09281_, _08726_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _60946_ (_09282_, _09281_, _09280_);
  nand _60947_ (_09283_, _09282_, _09131_);
  nand _60948_ (_09284_, _09283_, _09279_);
  nand _60949_ (_09285_, _09284_, _08719_);
  nand _60950_ (_09286_, _09285_, _09275_);
  nand _60951_ (_09287_, _09286_, _08709_);
  nand _60952_ (_09288_, _08719_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _60953_ (_09289_, _08718_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor _60954_ (_09290_, _09289_, _08734_);
  and _60955_ (_09291_, _09290_, _09288_);
  nand _60956_ (_09292_, _08719_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand _60957_ (_09293_, _08718_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _60958_ (_09294_, _09293_, _08734_);
  and _60959_ (_09295_, _09294_, _09292_);
  or _60960_ (_09296_, _09295_, _09291_);
  and _60961_ (_09297_, _09296_, _08726_);
  nand _60962_ (_09298_, _08719_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _60963_ (_09299_, _08718_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor _60964_ (_09300_, _09299_, _08734_);
  and _60965_ (_09301_, _09300_, _09298_);
  nand _60966_ (_09302_, _08719_, \oc8051_golden_model_1.IRAM[1] [3]);
  nand _60967_ (_09303_, _08718_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _60968_ (_09304_, _09303_, _08734_);
  and _60969_ (_09305_, _09304_, _09302_);
  or _60970_ (_09306_, _09305_, _09301_);
  and _60971_ (_09307_, _09306_, _09126_);
  or _60972_ (_09308_, _09307_, _09297_);
  nand _60973_ (_09309_, _09308_, _08708_);
  and _60974_ (_09310_, _09309_, _09287_);
  not _60975_ (_09311_, _09310_);
  or _60976_ (_09312_, _09126_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _60977_ (_09313_, _08726_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _60978_ (_09314_, _09313_, _09312_);
  nand _60979_ (_09315_, _09314_, _08734_);
  or _60980_ (_09316_, _09126_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _60981_ (_09317_, _08726_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _60982_ (_09318_, _09317_, _09316_);
  nand _60983_ (_09319_, _09318_, _09131_);
  nand _60984_ (_09320_, _09319_, _09315_);
  nand _60985_ (_09321_, _09320_, _08718_);
  or _60986_ (_09322_, _09126_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _60987_ (_09323_, _08726_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _60988_ (_09324_, _09323_, _09322_);
  nand _60989_ (_09325_, _09324_, _08734_);
  or _60990_ (_09326_, _09126_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _60991_ (_09327_, _08726_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _60992_ (_09328_, _09327_, _09326_);
  nand _60993_ (_09329_, _09328_, _09131_);
  nand _60994_ (_09330_, _09329_, _09325_);
  nand _60995_ (_09331_, _09330_, _08719_);
  nand _60996_ (_09332_, _09331_, _09321_);
  nand _60997_ (_09333_, _09332_, _08709_);
  nand _60998_ (_09334_, _08719_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _60999_ (_09335_, _08718_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor _61000_ (_09336_, _09335_, _08734_);
  and _61001_ (_09337_, _09336_, _09334_);
  nand _61002_ (_09338_, _08719_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand _61003_ (_09339_, _08718_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _61004_ (_09340_, _09339_, _08734_);
  and _61005_ (_09341_, _09340_, _09338_);
  or _61006_ (_09342_, _09341_, _09337_);
  and _61007_ (_09343_, _09342_, _08726_);
  nand _61008_ (_09344_, _08719_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _61009_ (_09345_, _08718_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor _61010_ (_09346_, _09345_, _08734_);
  and _61011_ (_09347_, _09346_, _09344_);
  nand _61012_ (_09348_, _08719_, \oc8051_golden_model_1.IRAM[1] [2]);
  nand _61013_ (_09349_, _08718_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _61014_ (_09350_, _09349_, _08734_);
  and _61015_ (_09351_, _09350_, _09348_);
  or _61016_ (_09352_, _09351_, _09347_);
  and _61017_ (_09353_, _09352_, _09126_);
  or _61018_ (_09354_, _09353_, _09343_);
  nand _61019_ (_09355_, _09354_, _08708_);
  and _61020_ (_09356_, _09355_, _09333_);
  not _61021_ (_09357_, _09356_);
  or _61022_ (_09358_, _09126_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _61023_ (_09359_, _08726_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _61024_ (_09360_, _09359_, _09358_);
  nand _61025_ (_09361_, _09360_, _08734_);
  nand _61026_ (_09362_, _08726_, _07436_);
  or _61027_ (_09363_, _08726_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _61028_ (_09364_, _09363_, _09362_);
  nand _61029_ (_09365_, _09364_, _09131_);
  nand _61030_ (_09366_, _09365_, _09361_);
  nand _61031_ (_09367_, _09366_, _08718_);
  or _61032_ (_09368_, _09126_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _61033_ (_09369_, _08726_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _61034_ (_09370_, _09369_, _09368_);
  nand _61035_ (_09371_, _09370_, _08734_);
  nand _61036_ (_09372_, _08726_, _07424_);
  or _61037_ (_09373_, _08726_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _61038_ (_09374_, _09373_, _09372_);
  nand _61039_ (_09375_, _09374_, _09131_);
  nand _61040_ (_09376_, _09375_, _09371_);
  nand _61041_ (_09377_, _09376_, _08719_);
  nand _61042_ (_09378_, _09377_, _09367_);
  nand _61043_ (_09379_, _09378_, _08709_);
  or _61044_ (_09380_, _08718_, _07402_);
  and _61045_ (_09381_, _08718_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor _61046_ (_09382_, _09381_, _08734_);
  and _61047_ (_09383_, _09382_, _09380_);
  nand _61048_ (_09384_, _08719_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand _61049_ (_09385_, _08718_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _61050_ (_09386_, _09385_, _08734_);
  and _61051_ (_09387_, _09386_, _09384_);
  or _61052_ (_09388_, _09387_, _09383_);
  and _61053_ (_09389_, _09388_, _08726_);
  or _61054_ (_09390_, _08718_, _07400_);
  and _61055_ (_09391_, _08718_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor _61056_ (_09392_, _09391_, _08734_);
  and _61057_ (_09393_, _09392_, _09390_);
  nand _61058_ (_09394_, _08719_, \oc8051_golden_model_1.IRAM[1] [1]);
  nand _61059_ (_09395_, _08718_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _61060_ (_09396_, _09395_, _08734_);
  and _61061_ (_09397_, _09396_, _09394_);
  or _61062_ (_09398_, _09397_, _09393_);
  and _61063_ (_09399_, _09398_, _09126_);
  or _61064_ (_09400_, _09399_, _09389_);
  nand _61065_ (_09401_, _09400_, _08708_);
  and _61066_ (_09402_, _09401_, _09379_);
  nand _61067_ (_09403_, _08726_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _61068_ (_09404_, _08726_, _07242_);
  and _61069_ (_09405_, _09404_, _09403_);
  nand _61070_ (_09406_, _09405_, _08734_);
  nand _61071_ (_09407_, _08726_, _07237_);
  or _61072_ (_09408_, _08726_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _61073_ (_09409_, _09408_, _09407_);
  nand _61074_ (_09410_, _09409_, _09131_);
  nand _61075_ (_09411_, _09410_, _09406_);
  nand _61076_ (_09412_, _09411_, _08718_);
  or _61077_ (_09413_, _09126_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _61078_ (_09414_, _08726_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _61079_ (_09415_, _09414_, _09413_);
  nand _61080_ (_09416_, _09415_, _08734_);
  or _61081_ (_09417_, _09126_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _61082_ (_09418_, _08726_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _61083_ (_09419_, _09418_, _09417_);
  nand _61084_ (_09420_, _09419_, _09131_);
  nand _61085_ (_09421_, _09420_, _09416_);
  nand _61086_ (_09422_, _09421_, _08719_);
  nand _61087_ (_09423_, _09422_, _09412_);
  nand _61088_ (_09424_, _09423_, _08709_);
  nand _61089_ (_09425_, _08719_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _61090_ (_09426_, _08718_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor _61091_ (_09427_, _09426_, _08734_);
  and _61092_ (_09428_, _09427_, _09425_);
  nand _61093_ (_09429_, _08719_, \oc8051_golden_model_1.IRAM[0] [0]);
  nand _61094_ (_09430_, _08718_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _61095_ (_09431_, _09430_, _08734_);
  and _61096_ (_09432_, _09431_, _09429_);
  or _61097_ (_09433_, _09432_, _09428_);
  and _61098_ (_09434_, _09433_, _08726_);
  nand _61099_ (_09435_, _08719_, \oc8051_golden_model_1.IRAM[3] [0]);
  and _61100_ (_09436_, _08718_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor _61101_ (_09437_, _09436_, _08734_);
  and _61102_ (_09438_, _09437_, _09435_);
  nand _61103_ (_09439_, _08719_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand _61104_ (_09440_, _08718_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _61105_ (_09441_, _09440_, _08734_);
  and _61106_ (_09442_, _09441_, _09439_);
  or _61107_ (_09443_, _09442_, _09438_);
  and _61108_ (_09444_, _09443_, _09126_);
  or _61109_ (_09445_, _09444_, _09434_);
  nand _61110_ (_09446_, _09445_, _08708_);
  and _61111_ (_09447_, _09446_, _09424_);
  nor _61112_ (_09448_, _09447_, _09402_);
  and _61113_ (_09449_, _09448_, _09357_);
  and _61114_ (_09450_, _09449_, _09311_);
  and _61115_ (_09451_, _09450_, _09265_);
  and _61116_ (_09452_, _09451_, _09219_);
  and _61117_ (_09453_, _09452_, _09173_);
  or _61118_ (_09454_, _09453_, _08778_);
  nand _61119_ (_09455_, _09453_, _08778_);
  and _61120_ (_09456_, _09455_, _09454_);
  or _61121_ (_09457_, _09456_, _07361_);
  not _61122_ (_09458_, _07359_);
  nand _61123_ (_09459_, _05985_, _05848_);
  or _61124_ (_09460_, _09459_, _08683_);
  and _61125_ (_09461_, _09460_, _09458_);
  and _61126_ (_09462_, _09461_, _09457_);
  and _61127_ (_09463_, _09462_, _09125_);
  and _61128_ (_09464_, _08791_, _07359_);
  or _61129_ (_09465_, _09464_, _06503_);
  or _61130_ (_09466_, _09465_, _09463_);
  and _61131_ (_09467_, _09466_, _08616_);
  or _61132_ (_09468_, _09467_, _05998_);
  and _61133_ (_09469_, _08814_, _05998_);
  nor _61134_ (_09470_, _09469_, _06272_);
  and _61135_ (_09471_, _09470_, _09468_);
  and _61136_ (_09472_, _08668_, _06272_);
  nor _61137_ (_09473_, _07591_, _07581_);
  not _61138_ (_09474_, _09473_);
  or _61139_ (_09475_, _09474_, _09472_);
  or _61140_ (_09476_, _09475_, _09471_);
  not _61141_ (_09477_, _08209_);
  not _61142_ (_09478_, _08305_);
  not _61143_ (_09479_, _08596_);
  not _61144_ (_09480_, _07680_);
  not _61145_ (_09481_, _07854_);
  not _61146_ (_09482_, _07448_);
  and _61147_ (_09483_, _09482_, _07250_);
  and _61148_ (_09484_, _09483_, _09481_);
  and _61149_ (_09485_, _09484_, _09480_);
  and _61150_ (_09486_, _09485_, _09479_);
  and _61151_ (_09487_, _09486_, _09478_);
  and _61152_ (_09488_, _09487_, _09477_);
  nor _61153_ (_09489_, _09488_, _08107_);
  and _61154_ (_09490_, _09488_, _08107_);
  or _61155_ (_09491_, _09490_, _09489_);
  or _61156_ (_09492_, _09491_, _09473_);
  and _61157_ (_09493_, _09492_, _09476_);
  or _61158_ (_09494_, _09493_, _07055_);
  not _61159_ (_09495_, _07379_);
  not _61160_ (_09496_, _08778_);
  and _61161_ (_09497_, _09447_, _09402_);
  and _61162_ (_09498_, _09497_, _09356_);
  and _61163_ (_09499_, _09498_, _09310_);
  and _61164_ (_09500_, _09499_, _09264_);
  and _61165_ (_09501_, _09500_, _09218_);
  and _61166_ (_09502_, _09501_, _09172_);
  nor _61167_ (_09503_, _09502_, _09496_);
  and _61168_ (_09504_, _09502_, _09496_);
  or _61169_ (_09505_, _09504_, _09503_);
  or _61170_ (_09507_, _09505_, _07375_);
  and _61171_ (_09508_, _09507_, _09495_);
  and _61172_ (_09509_, _09508_, _09494_);
  or _61173_ (_09510_, _09509_, _08606_);
  and _61174_ (_09511_, _09510_, _07631_);
  and _61175_ (_09512_, _09511_, _07944_);
  or _61176_ (_09513_, _09512_, _07945_);
  not _61177_ (_09514_, _07386_);
  and _61178_ (_09515_, _07688_, _06342_);
  and _61179_ (_09516_, _07687_, _06342_);
  nor _61180_ (_09517_, _09516_, _07690_);
  nor _61181_ (_09518_, _09517_, _09515_);
  not _61182_ (_09519_, _09516_);
  or _61183_ (_09520_, _07803_, _07387_);
  and _61184_ (_09521_, _09520_, _09519_);
  and _61185_ (_09522_, _07367_, _07564_);
  and _61186_ (_09523_, _09522_, _06019_);
  and _61187_ (_09524_, _09523_, _07598_);
  nor _61188_ (_09525_, _09524_, _07543_);
  and _61189_ (_09526_, _09525_, _09521_);
  nand _61190_ (_09528_, _09526_, _09518_);
  or _61191_ (_09529_, _09528_, _09514_);
  and _61192_ (_09530_, _09529_, _09513_);
  and _61193_ (_09531_, _09525_, _09518_);
  and _61194_ (_09532_, _09531_, _09521_);
  and _61195_ (_09533_, _09532_, _07386_);
  not _61196_ (_09534_, _06503_);
  and _61197_ (_09535_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _61198_ (_09536_, _09535_, \oc8051_golden_model_1.PC [10]);
  and _61199_ (_09537_, _09536_, _08618_);
  and _61200_ (_09538_, _09537_, \oc8051_golden_model_1.PC [11]);
  and _61201_ (_09539_, _09538_, \oc8051_golden_model_1.PC [12]);
  and _61202_ (_09540_, _09539_, \oc8051_golden_model_1.PC [13]);
  and _61203_ (_09541_, _09540_, \oc8051_golden_model_1.PC [14]);
  nor _61204_ (_09542_, _09541_, \oc8051_golden_model_1.PC [15]);
  and _61205_ (_09543_, _09535_, _08618_);
  and _61206_ (_09544_, _09543_, \oc8051_golden_model_1.PC [10]);
  and _61207_ (_09545_, _09544_, \oc8051_golden_model_1.PC [11]);
  and _61208_ (_09546_, _09545_, \oc8051_golden_model_1.PC [12]);
  and _61209_ (_09547_, _09546_, \oc8051_golden_model_1.PC [13]);
  and _61210_ (_09548_, _09547_, \oc8051_golden_model_1.PC [14]);
  and _61211_ (_09549_, _09548_, \oc8051_golden_model_1.PC [15]);
  nor _61212_ (_09550_, _09549_, _09542_);
  and _61213_ (_09551_, _09550_, _09534_);
  and _61214_ (_09552_, _09536_, _08612_);
  and _61215_ (_09553_, _09552_, \oc8051_golden_model_1.PC [11]);
  and _61216_ (_09554_, _09553_, \oc8051_golden_model_1.PC [12]);
  and _61217_ (_09555_, _09554_, \oc8051_golden_model_1.PC [13]);
  and _61218_ (_09556_, _09555_, \oc8051_golden_model_1.PC [14]);
  nor _61219_ (_09557_, _09556_, \oc8051_golden_model_1.PC [15]);
  and _61220_ (_09558_, _09535_, _08612_);
  and _61221_ (_09559_, _09558_, \oc8051_golden_model_1.PC [10]);
  and _61222_ (_09560_, _09559_, \oc8051_golden_model_1.PC [11]);
  and _61223_ (_09561_, _09560_, \oc8051_golden_model_1.PC [12]);
  and _61224_ (_09562_, _09561_, \oc8051_golden_model_1.PC [13]);
  and _61225_ (_09563_, _09562_, \oc8051_golden_model_1.PC [14]);
  and _61226_ (_09564_, _09563_, \oc8051_golden_model_1.PC [15]);
  nor _61227_ (_09565_, _09564_, _09557_);
  and _61228_ (_09566_, _09565_, _06503_);
  or _61229_ (_09567_, _09566_, _09551_);
  and _61230_ (_09568_, _09567_, _09525_);
  and _61231_ (_09569_, _09568_, _09533_);
  or _61232_ (_41495_, _09569_, _09530_);
  not _61233_ (_09570_, \oc8051_golden_model_1.B [7]);
  nor _61234_ (_09571_, _01442_, _09570_);
  not _61235_ (_09572_, _06333_);
  nor _61236_ (_09573_, _08025_, _09570_);
  not _61237_ (_09574_, _08025_);
  nor _61238_ (_09575_, _08107_, _09574_);
  or _61239_ (_09576_, _09575_, _09573_);
  or _61240_ (_09577_, _09576_, _06327_);
  nor _61241_ (_09578_, _08637_, _09570_);
  and _61242_ (_09579_, _08668_, _08637_);
  or _61243_ (_09580_, _09579_, _09578_);
  and _61244_ (_09581_, _09580_, _06352_);
  and _61245_ (_09582_, _08791_, _08025_);
  or _61246_ (_09583_, _09582_, _09573_);
  or _61247_ (_09584_, _09583_, _07275_);
  and _61248_ (_09585_, _08025_, \oc8051_golden_model_1.ACC [7]);
  or _61249_ (_09586_, _09585_, _09573_);
  and _61250_ (_09587_, _09586_, _07259_);
  nor _61251_ (_09588_, _07259_, _09570_);
  or _61252_ (_09589_, _09588_, _06474_);
  or _61253_ (_09590_, _09589_, _09587_);
  and _61254_ (_09591_, _09590_, _06357_);
  and _61255_ (_09592_, _09591_, _09584_);
  and _61256_ (_09593_, _08672_, _08637_);
  or _61257_ (_09594_, _09593_, _09578_);
  and _61258_ (_09595_, _09594_, _06356_);
  or _61259_ (_09596_, _09595_, _06410_);
  or _61260_ (_09597_, _09596_, _09592_);
  or _61261_ (_09598_, _09576_, _06772_);
  and _61262_ (_09599_, _09598_, _09597_);
  or _61263_ (_09600_, _09599_, _06417_);
  or _61264_ (_09601_, _09586_, _06426_);
  and _61265_ (_09602_, _09601_, _06353_);
  and _61266_ (_09603_, _09602_, _09600_);
  or _61267_ (_09604_, _09603_, _09581_);
  and _61268_ (_09605_, _09604_, _06346_);
  and _61269_ (_09606_, _06489_, _06443_);
  or _61270_ (_09607_, _09578_, _08809_);
  and _61271_ (_09608_, _09594_, _06345_);
  and _61272_ (_09609_, _09608_, _09607_);
  or _61273_ (_09610_, _09609_, _09606_);
  or _61274_ (_09611_, _09610_, _09605_);
  not _61275_ (_09612_, _09606_);
  and _61276_ (_09613_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _61277_ (_09614_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _61278_ (_09615_, _09614_, _09613_);
  and _61279_ (_09616_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and _61280_ (_09617_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and _61281_ (_09618_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _61282_ (_09619_, _09618_, _09617_);
  nor _61283_ (_09620_, _09619_, _09615_);
  and _61284_ (_09621_, _09620_, _09616_);
  nor _61285_ (_09622_, _09621_, _09615_);
  and _61286_ (_09623_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _61287_ (_09624_, _09623_, _09617_);
  and _61288_ (_09625_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _61289_ (_09626_, _09625_, _09613_);
  nor _61290_ (_09627_, _09626_, _09624_);
  not _61291_ (_09628_, _09627_);
  nor _61292_ (_09629_, _09628_, _09622_);
  and _61293_ (_09630_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _61294_ (_09631_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and _61295_ (_09632_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and _61296_ (_09633_, _09632_, _09631_);
  nor _61297_ (_09634_, _09632_, _09631_);
  nor _61298_ (_09635_, _09634_, _09633_);
  and _61299_ (_09636_, _09635_, _09630_);
  nor _61300_ (_09637_, _09635_, _09630_);
  nor _61301_ (_09638_, _09637_, _09636_);
  and _61302_ (_09639_, _09628_, _09622_);
  nor _61303_ (_09640_, _09639_, _09629_);
  and _61304_ (_09641_, _09640_, _09638_);
  nor _61305_ (_09642_, _09641_, _09629_);
  not _61306_ (_09643_, _09617_);
  and _61307_ (_09644_, _09623_, _09643_);
  and _61308_ (_09645_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and _61309_ (_09646_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _61310_ (_09647_, _09646_, _09631_);
  and _61311_ (_09648_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and _61312_ (_09649_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor _61313_ (_09650_, _09649_, _09648_);
  nor _61314_ (_09651_, _09650_, _09647_);
  and _61315_ (_09652_, _09651_, _09645_);
  nor _61316_ (_09653_, _09651_, _09645_);
  nor _61317_ (_09654_, _09653_, _09652_);
  and _61318_ (_09655_, _09654_, _09644_);
  nor _61319_ (_09656_, _09654_, _09644_);
  nor _61320_ (_09657_, _09656_, _09655_);
  not _61321_ (_09658_, _09657_);
  nor _61322_ (_09659_, _09658_, _09642_);
  and _61323_ (_09660_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _61324_ (_09661_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and _61325_ (_09662_, _09661_, _09660_);
  nor _61326_ (_09663_, _09636_, _09633_);
  and _61327_ (_09664_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and _61328_ (_09665_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _61329_ (_09666_, _09665_, _09664_);
  nor _61330_ (_09667_, _09665_, _09664_);
  nor _61331_ (_09668_, _09667_, _09666_);
  not _61332_ (_09669_, _09668_);
  nor _61333_ (_09670_, _09669_, _09663_);
  and _61334_ (_09671_, _09669_, _09663_);
  nor _61335_ (_09672_, _09671_, _09670_);
  and _61336_ (_09673_, _09672_, _09662_);
  nor _61337_ (_09674_, _09672_, _09662_);
  nor _61338_ (_09675_, _09674_, _09673_);
  and _61339_ (_09676_, _09658_, _09642_);
  nor _61340_ (_09677_, _09676_, _09659_);
  and _61341_ (_09678_, _09677_, _09675_);
  nor _61342_ (_09679_, _09678_, _09659_);
  nor _61343_ (_09680_, _09652_, _09647_);
  and _61344_ (_09682_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and _61345_ (_09683_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and _61346_ (_09685_, _09683_, _09682_);
  nor _61347_ (_09686_, _09683_, _09682_);
  nor _61348_ (_09688_, _09686_, _09685_);
  not _61349_ (_09689_, _09688_);
  nor _61350_ (_09691_, _09689_, _09680_);
  and _61351_ (_09692_, _09689_, _09680_);
  nor _61352_ (_09694_, _09692_, _09691_);
  and _61353_ (_09695_, _09694_, _09666_);
  nor _61354_ (_09697_, _09694_, _09666_);
  nor _61355_ (_09698_, _09697_, _09695_);
  nor _61356_ (_09700_, _09655_, _09624_);
  and _61357_ (_09701_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and _61358_ (_09703_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _61359_ (_09704_, _09703_, _09646_);
  nor _61360_ (_09706_, _09703_, _09646_);
  nor _61361_ (_09707_, _09706_, _09704_);
  and _61362_ (_09709_, _09707_, _09701_);
  nor _61363_ (_09710_, _09707_, _09701_);
  nor _61364_ (_09712_, _09710_, _09709_);
  not _61365_ (_09713_, _09712_);
  nor _61366_ (_09715_, _09713_, _09700_);
  and _61367_ (_09716_, _09713_, _09700_);
  nor _61368_ (_09718_, _09716_, _09715_);
  and _61369_ (_09719_, _09718_, _09698_);
  nor _61370_ (_09720_, _09718_, _09698_);
  nor _61371_ (_09721_, _09720_, _09719_);
  not _61372_ (_09722_, _09721_);
  nor _61373_ (_09723_, _09722_, _09679_);
  nor _61374_ (_09724_, _09673_, _09670_);
  not _61375_ (_09725_, _09724_);
  and _61376_ (_09726_, _09722_, _09679_);
  nor _61377_ (_09727_, _09726_, _09723_);
  and _61378_ (_09728_, _09727_, _09725_);
  nor _61379_ (_09729_, _09728_, _09723_);
  nor _61380_ (_09730_, _09695_, _09691_);
  not _61381_ (_09731_, _09730_);
  nor _61382_ (_09732_, _09719_, _09715_);
  not _61383_ (_09733_, _09732_);
  and _61384_ (_09734_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _61385_ (_09735_, _09734_, _09646_);
  and _61386_ (_09736_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _61387_ (_09737_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _61388_ (_09738_, _09737_, _09736_);
  nor _61389_ (_09739_, _09738_, _09735_);
  nor _61390_ (_09740_, _09709_, _09704_);
  and _61391_ (_09741_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and _61392_ (_09742_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and _61393_ (_09743_, _09742_, _09741_);
  nor _61394_ (_09744_, _09742_, _09741_);
  nor _61395_ (_09745_, _09744_, _09743_);
  not _61396_ (_09746_, _09745_);
  nor _61397_ (_09747_, _09746_, _09740_);
  and _61398_ (_09748_, _09746_, _09740_);
  nor _61399_ (_09749_, _09748_, _09747_);
  and _61400_ (_09750_, _09749_, _09685_);
  nor _61401_ (_09751_, _09749_, _09685_);
  nor _61402_ (_09752_, _09751_, _09750_);
  and _61403_ (_09753_, _09752_, _09739_);
  nor _61404_ (_09754_, _09752_, _09739_);
  nor _61405_ (_09755_, _09754_, _09753_);
  and _61406_ (_09756_, _09755_, _09733_);
  nor _61407_ (_09757_, _09755_, _09733_);
  nor _61408_ (_09758_, _09757_, _09756_);
  and _61409_ (_09759_, _09758_, _09731_);
  nor _61410_ (_09760_, _09758_, _09731_);
  nor _61411_ (_09761_, _09760_, _09759_);
  not _61412_ (_09762_, _09761_);
  nor _61413_ (_09763_, _09762_, _09729_);
  nor _61414_ (_09764_, _09759_, _09756_);
  nor _61415_ (_09765_, _09750_, _09747_);
  not _61416_ (_09766_, _09765_);
  and _61417_ (_09767_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and _61418_ (_09768_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _61419_ (_09769_, _09768_, _09767_);
  nor _61420_ (_09770_, _09768_, _09767_);
  nor _61421_ (_09771_, _09770_, _09769_);
  and _61422_ (_09772_, _09771_, _09735_);
  nor _61423_ (_09773_, _09771_, _09735_);
  nor _61424_ (_09774_, _09773_, _09772_);
  and _61425_ (_09775_, _09774_, _09743_);
  nor _61426_ (_09777_, _09774_, _09743_);
  nor _61427_ (_09779_, _09777_, _09775_);
  and _61428_ (_09780_, _09779_, _09734_);
  nor _61429_ (_09782_, _09779_, _09734_);
  nor _61430_ (_09783_, _09782_, _09780_);
  and _61431_ (_09785_, _09783_, _09753_);
  nor _61432_ (_09786_, _09783_, _09753_);
  nor _61433_ (_09788_, _09786_, _09785_);
  and _61434_ (_09789_, _09788_, _09766_);
  nor _61435_ (_09791_, _09788_, _09766_);
  nor _61436_ (_09792_, _09791_, _09789_);
  not _61437_ (_09794_, _09792_);
  nor _61438_ (_09795_, _09794_, _09764_);
  and _61439_ (_09797_, _09794_, _09764_);
  nor _61440_ (_09798_, _09797_, _09795_);
  and _61441_ (_09800_, _09798_, _09763_);
  nor _61442_ (_09801_, _09789_, _09785_);
  nor _61443_ (_09803_, _09775_, _09772_);
  not _61444_ (_09804_, _09803_);
  and _61445_ (_09806_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and _61446_ (_09807_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _61447_ (_09809_, _09807_, _09806_);
  nor _61448_ (_09810_, _09807_, _09806_);
  nor _61449_ (_09812_, _09810_, _09809_);
  and _61450_ (_09813_, _09812_, _09769_);
  nor _61451_ (_09814_, _09812_, _09769_);
  nor _61452_ (_09815_, _09814_, _09813_);
  and _61453_ (_09816_, _09815_, _09780_);
  nor _61454_ (_09817_, _09815_, _09780_);
  nor _61455_ (_09818_, _09817_, _09816_);
  and _61456_ (_09819_, _09818_, _09804_);
  nor _61457_ (_09820_, _09818_, _09804_);
  nor _61458_ (_09821_, _09820_, _09819_);
  not _61459_ (_09822_, _09821_);
  nor _61460_ (_09823_, _09822_, _09801_);
  and _61461_ (_09824_, _09822_, _09801_);
  nor _61462_ (_09825_, _09824_, _09823_);
  and _61463_ (_09826_, _09825_, _09795_);
  nor _61464_ (_09827_, _09825_, _09795_);
  nor _61465_ (_09828_, _09827_, _09826_);
  and _61466_ (_09829_, _09828_, _09800_);
  nor _61467_ (_09830_, _09828_, _09800_);
  nor _61468_ (_09831_, _09830_, _09829_);
  and _61469_ (_09832_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and _61470_ (_09833_, _09832_, _09617_);
  and _61471_ (_09834_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and _61472_ (_09835_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor _61473_ (_09836_, _09835_, _09614_);
  nor _61474_ (_09837_, _09836_, _09833_);
  and _61475_ (_09838_, _09837_, _09834_);
  nor _61476_ (_09839_, _09838_, _09833_);
  not _61477_ (_09840_, _09839_);
  nor _61478_ (_09841_, _09620_, _09616_);
  nor _61479_ (_09842_, _09841_, _09621_);
  and _61480_ (_09843_, _09842_, _09840_);
  and _61481_ (_09844_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _61482_ (_09845_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and _61483_ (_09846_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _61484_ (_09847_, _09846_, _09845_);
  nor _61485_ (_09848_, _09846_, _09845_);
  nor _61486_ (_09849_, _09848_, _09847_);
  and _61487_ (_09850_, _09849_, _09844_);
  nor _61488_ (_09851_, _09849_, _09844_);
  nor _61489_ (_09852_, _09851_, _09850_);
  nor _61490_ (_09853_, _09842_, _09840_);
  nor _61491_ (_09854_, _09853_, _09843_);
  and _61492_ (_09855_, _09854_, _09852_);
  nor _61493_ (_09856_, _09855_, _09843_);
  nor _61494_ (_09857_, _09640_, _09638_);
  nor _61495_ (_09858_, _09857_, _09641_);
  not _61496_ (_09859_, _09858_);
  nor _61497_ (_09860_, _09859_, _09856_);
  and _61498_ (_09861_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _61499_ (_09862_, _09861_, _09661_);
  nor _61500_ (_09863_, _09850_, _09847_);
  nor _61501_ (_09864_, _09661_, _09660_);
  nor _61502_ (_09865_, _09864_, _09662_);
  not _61503_ (_09866_, _09865_);
  nor _61504_ (_09867_, _09866_, _09863_);
  and _61505_ (_09868_, _09866_, _09863_);
  nor _61506_ (_09869_, _09868_, _09867_);
  and _61507_ (_09870_, _09869_, _09862_);
  nor _61508_ (_09871_, _09869_, _09862_);
  nor _61509_ (_09872_, _09871_, _09870_);
  and _61510_ (_09873_, _09859_, _09856_);
  nor _61511_ (_09874_, _09873_, _09860_);
  and _61512_ (_09875_, _09874_, _09872_);
  nor _61513_ (_09876_, _09875_, _09860_);
  nor _61514_ (_09877_, _09677_, _09675_);
  nor _61515_ (_09878_, _09877_, _09678_);
  not _61516_ (_09879_, _09878_);
  nor _61517_ (_09880_, _09879_, _09876_);
  nor _61518_ (_09881_, _09870_, _09867_);
  not _61519_ (_09882_, _09881_);
  and _61520_ (_09883_, _09879_, _09876_);
  nor _61521_ (_09884_, _09883_, _09880_);
  and _61522_ (_09885_, _09884_, _09882_);
  nor _61523_ (_09886_, _09885_, _09880_);
  nor _61524_ (_09887_, _09727_, _09725_);
  nor _61525_ (_09888_, _09887_, _09728_);
  not _61526_ (_09889_, _09888_);
  nor _61527_ (_09890_, _09889_, _09886_);
  and _61528_ (_09891_, _09762_, _09729_);
  nor _61529_ (_09892_, _09891_, _09763_);
  and _61530_ (_09893_, _09892_, _09890_);
  nor _61531_ (_09894_, _09798_, _09763_);
  nor _61532_ (_09895_, _09894_, _09800_);
  nand _61533_ (_09896_, _09895_, _09893_);
  and _61534_ (_09897_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and _61535_ (_09898_, _09897_, _09832_);
  and _61536_ (_09899_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _61537_ (_09900_, _09897_, _09832_);
  nor _61538_ (_09901_, _09900_, _09898_);
  and _61539_ (_09902_, _09901_, _09899_);
  nor _61540_ (_09903_, _09902_, _09898_);
  not _61541_ (_09904_, _09903_);
  nor _61542_ (_09905_, _09837_, _09834_);
  nor _61543_ (_09906_, _09905_, _09838_);
  and _61544_ (_09907_, _09906_, _09904_);
  and _61545_ (_09908_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and _61546_ (_09909_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _61547_ (_09910_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _61548_ (_09911_, _09910_, _09909_);
  nor _61549_ (_09912_, _09910_, _09909_);
  nor _61550_ (_09913_, _09912_, _09911_);
  and _61551_ (_09914_, _09913_, _09908_);
  nor _61552_ (_09915_, _09913_, _09908_);
  nor _61553_ (_09916_, _09915_, _09914_);
  nor _61554_ (_09917_, _09906_, _09904_);
  nor _61555_ (_09918_, _09917_, _09907_);
  and _61556_ (_09919_, _09918_, _09916_);
  nor _61557_ (_09920_, _09919_, _09907_);
  not _61558_ (_09921_, _09920_);
  nor _61559_ (_09922_, _09854_, _09852_);
  nor _61560_ (_09923_, _09922_, _09855_);
  and _61561_ (_09924_, _09923_, _09921_);
  nor _61562_ (_09925_, _09914_, _09911_);
  and _61563_ (_09926_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and _61564_ (_09927_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor _61565_ (_09928_, _09927_, _09926_);
  nor _61566_ (_09929_, _09928_, _09862_);
  not _61567_ (_09930_, _09929_);
  nor _61568_ (_09931_, _09930_, _09925_);
  and _61569_ (_09932_, _09930_, _09925_);
  nor _61570_ (_09933_, _09932_, _09931_);
  nor _61571_ (_09934_, _09923_, _09921_);
  nor _61572_ (_09935_, _09934_, _09924_);
  and _61573_ (_09936_, _09935_, _09933_);
  nor _61574_ (_09937_, _09936_, _09924_);
  nor _61575_ (_09938_, _09874_, _09872_);
  nor _61576_ (_09939_, _09938_, _09875_);
  not _61577_ (_09940_, _09939_);
  nor _61578_ (_09941_, _09940_, _09937_);
  and _61579_ (_09942_, _09940_, _09937_);
  nor _61580_ (_09943_, _09942_, _09941_);
  and _61581_ (_09944_, _09943_, _09931_);
  nor _61582_ (_09945_, _09944_, _09941_);
  nor _61583_ (_09946_, _09884_, _09882_);
  nor _61584_ (_09947_, _09946_, _09885_);
  not _61585_ (_09948_, _09947_);
  nor _61586_ (_09949_, _09948_, _09945_);
  and _61587_ (_09950_, _09889_, _09886_);
  nor _61588_ (_09951_, _09950_, _09890_);
  and _61589_ (_09952_, _09951_, _09949_);
  nor _61590_ (_09953_, _09892_, _09890_);
  nor _61591_ (_09954_, _09953_, _09893_);
  and _61592_ (_09955_, _09954_, _09952_);
  nor _61593_ (_09956_, _09954_, _09952_);
  nor _61594_ (_09957_, _09956_, _09955_);
  and _61595_ (_09958_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and _61596_ (_09959_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _61597_ (_09960_, _09959_, _09958_);
  and _61598_ (_09961_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _61599_ (_09962_, _09959_, _09958_);
  nor _61600_ (_09963_, _09962_, _09960_);
  and _61601_ (_09964_, _09963_, _09961_);
  nor _61602_ (_09965_, _09964_, _09960_);
  not _61603_ (_09966_, _09965_);
  nor _61604_ (_09967_, _09901_, _09899_);
  nor _61605_ (_09968_, _09967_, _09902_);
  and _61606_ (_09969_, _09968_, _09966_);
  and _61607_ (_09970_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _61608_ (_09971_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _61609_ (_09972_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and _61610_ (_09973_, _09972_, _09971_);
  nor _61611_ (_09974_, _09972_, _09971_);
  nor _61612_ (_09975_, _09974_, _09973_);
  and _61613_ (_09976_, _09975_, _09970_);
  nor _61614_ (_09977_, _09975_, _09970_);
  nor _61615_ (_09978_, _09977_, _09976_);
  nor _61616_ (_09979_, _09968_, _09966_);
  nor _61617_ (_09980_, _09979_, _09969_);
  and _61618_ (_09981_, _09980_, _09978_);
  nor _61619_ (_09982_, _09981_, _09969_);
  not _61620_ (_09983_, _09982_);
  nor _61621_ (_09984_, _09918_, _09916_);
  nor _61622_ (_09985_, _09984_, _09919_);
  and _61623_ (_09986_, _09985_, _09983_);
  not _61624_ (_09987_, _09861_);
  nor _61625_ (_09988_, _09976_, _09973_);
  nor _61626_ (_09989_, _09988_, _09987_);
  and _61627_ (_09990_, _09988_, _09987_);
  nor _61628_ (_09991_, _09990_, _09989_);
  nor _61629_ (_09992_, _09985_, _09983_);
  nor _61630_ (_09993_, _09992_, _09986_);
  and _61631_ (_09994_, _09993_, _09991_);
  nor _61632_ (_09995_, _09994_, _09986_);
  not _61633_ (_09996_, _09995_);
  nor _61634_ (_09997_, _09935_, _09933_);
  nor _61635_ (_09998_, _09997_, _09936_);
  and _61636_ (_09999_, _09998_, _09996_);
  nor _61637_ (_10000_, _09998_, _09996_);
  nor _61638_ (_10001_, _10000_, _09999_);
  and _61639_ (_10002_, _10001_, _09989_);
  nor _61640_ (_10003_, _10002_, _09999_);
  nor _61641_ (_10004_, _09943_, _09931_);
  nor _61642_ (_10005_, _10004_, _09944_);
  not _61643_ (_10006_, _10005_);
  nor _61644_ (_10007_, _10006_, _10003_);
  and _61645_ (_10008_, _09948_, _09945_);
  nor _61646_ (_10009_, _10008_, _09949_);
  and _61647_ (_10010_, _10009_, _10007_);
  nor _61648_ (_10011_, _09951_, _09949_);
  nor _61649_ (_10012_, _10011_, _09952_);
  nand _61650_ (_10013_, _10012_, _10010_);
  or _61651_ (_10014_, _10012_, _10010_);
  and _61652_ (_10015_, _10014_, _10013_);
  and _61653_ (_10016_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _61654_ (_10017_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _61655_ (_10018_, _10017_, _10016_);
  and _61656_ (_10019_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor _61657_ (_10020_, _10017_, _10016_);
  nor _61658_ (_10021_, _10020_, _10018_);
  and _61659_ (_10022_, _10021_, _10019_);
  nor _61660_ (_10023_, _10022_, _10018_);
  not _61661_ (_10024_, _10023_);
  nor _61662_ (_10025_, _09963_, _09961_);
  nor _61663_ (_10026_, _10025_, _09964_);
  and _61664_ (_10027_, _10026_, _10024_);
  and _61665_ (_10028_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _61666_ (_10029_, _10028_, _09972_);
  and _61667_ (_10030_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and _61668_ (_10031_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _61669_ (_10032_, _10031_, _10030_);
  nor _61670_ (_10033_, _10032_, _10029_);
  nor _61671_ (_10034_, _10026_, _10024_);
  nor _61672_ (_10035_, _10034_, _10027_);
  and _61673_ (_10036_, _10035_, _10033_);
  nor _61674_ (_10037_, _10036_, _10027_);
  not _61675_ (_10038_, _10037_);
  nor _61676_ (_10039_, _09980_, _09978_);
  nor _61677_ (_10040_, _10039_, _09981_);
  and _61678_ (_10041_, _10040_, _10038_);
  nor _61679_ (_10042_, _10040_, _10038_);
  nor _61680_ (_10043_, _10042_, _10041_);
  and _61681_ (_10044_, _10043_, _10029_);
  nor _61682_ (_10045_, _10044_, _10041_);
  not _61683_ (_10046_, _10045_);
  nor _61684_ (_10047_, _09993_, _09991_);
  nor _61685_ (_10048_, _10047_, _09994_);
  and _61686_ (_10049_, _10048_, _10046_);
  nor _61687_ (_10050_, _10001_, _09989_);
  nor _61688_ (_10051_, _10050_, _10002_);
  and _61689_ (_10052_, _10051_, _10049_);
  and _61690_ (_10053_, _10006_, _10003_);
  nor _61691_ (_10054_, _10053_, _10007_);
  and _61692_ (_10055_, _10054_, _10052_);
  nor _61693_ (_10056_, _10009_, _10007_);
  nor _61694_ (_10057_, _10056_, _10010_);
  and _61695_ (_10058_, _10057_, _10055_);
  nor _61696_ (_10059_, _10057_, _10055_);
  nor _61697_ (_10060_, _10059_, _10058_);
  and _61698_ (_10061_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _61699_ (_10062_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and _61700_ (_10063_, _10062_, _10061_);
  and _61701_ (_10064_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _61702_ (_10065_, _10062_, _10061_);
  nor _61703_ (_10066_, _10065_, _10063_);
  and _61704_ (_10067_, _10066_, _10064_);
  nor _61705_ (_10068_, _10067_, _10063_);
  not _61706_ (_10069_, _10068_);
  nor _61707_ (_10070_, _10021_, _10019_);
  nor _61708_ (_10071_, _10070_, _10022_);
  and _61709_ (_10072_, _10071_, _10069_);
  nor _61710_ (_10073_, _10071_, _10069_);
  nor _61711_ (_10074_, _10073_, _10072_);
  and _61712_ (_10075_, _10074_, _10028_);
  nor _61713_ (_10076_, _10075_, _10072_);
  not _61714_ (_10077_, _10076_);
  nor _61715_ (_10078_, _10035_, _10033_);
  nor _61716_ (_10079_, _10078_, _10036_);
  and _61717_ (_10080_, _10079_, _10077_);
  nor _61718_ (_10081_, _10043_, _10029_);
  nor _61719_ (_10082_, _10081_, _10044_);
  and _61720_ (_10083_, _10082_, _10080_);
  nor _61721_ (_10084_, _10048_, _10046_);
  nor _61722_ (_10085_, _10084_, _10049_);
  and _61723_ (_10086_, _10085_, _10083_);
  nor _61724_ (_10087_, _10051_, _10049_);
  nor _61725_ (_10088_, _10087_, _10052_);
  and _61726_ (_10089_, _10088_, _10086_);
  nor _61727_ (_10090_, _10054_, _10052_);
  nor _61728_ (_10091_, _10090_, _10055_);
  and _61729_ (_10092_, _10091_, _10089_);
  and _61730_ (_10093_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and _61731_ (_10094_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and _61732_ (_10095_, _10094_, _10093_);
  nor _61733_ (_10096_, _10066_, _10064_);
  nor _61734_ (_10097_, _10096_, _10067_);
  and _61735_ (_10098_, _10097_, _10095_);
  nor _61736_ (_10099_, _10074_, _10028_);
  nor _61737_ (_10100_, _10099_, _10075_);
  and _61738_ (_10101_, _10100_, _10098_);
  nor _61739_ (_10102_, _10079_, _10077_);
  nor _61740_ (_10103_, _10102_, _10080_);
  and _61741_ (_10104_, _10103_, _10101_);
  nor _61742_ (_10105_, _10082_, _10080_);
  nor _61743_ (_10106_, _10105_, _10083_);
  and _61744_ (_10107_, _10106_, _10104_);
  nor _61745_ (_10108_, _10085_, _10083_);
  nor _61746_ (_10109_, _10108_, _10086_);
  and _61747_ (_10110_, _10109_, _10107_);
  nor _61748_ (_10111_, _10088_, _10086_);
  nor _61749_ (_10112_, _10111_, _10089_);
  and _61750_ (_10113_, _10112_, _10110_);
  nor _61751_ (_10114_, _10091_, _10089_);
  nor _61752_ (_10115_, _10114_, _10092_);
  and _61753_ (_10116_, _10115_, _10113_);
  nor _61754_ (_10117_, _10116_, _10092_);
  not _61755_ (_10118_, _10117_);
  and _61756_ (_10119_, _10118_, _10060_);
  or _61757_ (_10120_, _10119_, _10058_);
  nand _61758_ (_10121_, _10120_, _10015_);
  and _61759_ (_10122_, _10121_, _10013_);
  not _61760_ (_10123_, _10122_);
  and _61761_ (_10124_, _10123_, _09957_);
  or _61762_ (_10125_, _10124_, _09955_);
  or _61763_ (_10126_, _09895_, _09893_);
  and _61764_ (_10127_, _10126_, _09896_);
  nand _61765_ (_10128_, _10127_, _10125_);
  and _61766_ (_10129_, _10128_, _09896_);
  not _61767_ (_10130_, _10129_);
  and _61768_ (_10131_, _10130_, _09831_);
  or _61769_ (_10132_, _10131_, _09829_);
  and _61770_ (_10133_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not _61771_ (_10134_, _10133_);
  nor _61772_ (_10135_, _10134_, _09768_);
  nor _61773_ (_10136_, _10135_, _09813_);
  nor _61774_ (_10137_, _09819_, _09816_);
  nor _61775_ (_10138_, _10137_, _10136_);
  and _61776_ (_10139_, _10137_, _10136_);
  nor _61777_ (_10140_, _10139_, _10138_);
  nor _61778_ (_10141_, _09826_, _09823_);
  not _61779_ (_10142_, _10141_);
  and _61780_ (_10143_, _10142_, _10140_);
  nor _61781_ (_10144_, _10142_, _10140_);
  nor _61782_ (_10145_, _10144_, _10143_);
  and _61783_ (_10146_, _10145_, _10132_);
  or _61784_ (_10147_, _10138_, _09809_);
  or _61785_ (_10148_, _10147_, _10143_);
  or _61786_ (_10149_, _10148_, _10146_);
  or _61787_ (_10150_, _10149_, _09612_);
  and _61788_ (_10151_, _10150_, _06340_);
  and _61789_ (_10152_, _10151_, _09611_);
  not _61790_ (_10153_, _06327_);
  and _61791_ (_10154_, _08828_, _08637_);
  or _61792_ (_10155_, _10154_, _09578_);
  and _61793_ (_10156_, _10155_, _06339_);
  or _61794_ (_10157_, _10156_, _10153_);
  or _61795_ (_10158_, _10157_, _10152_);
  and _61796_ (_10159_, _10158_, _09577_);
  or _61797_ (_10160_, _10159_, _09572_);
  and _61798_ (_10161_, _08778_, _08025_);
  or _61799_ (_10162_, _09573_, _06333_);
  or _61800_ (_10163_, _10162_, _10161_);
  and _61801_ (_10164_, _10163_, _06313_);
  and _61802_ (_10165_, _10164_, _10160_);
  and _61803_ (_10166_, _06489_, _06002_);
  and _61804_ (_10167_, _09076_, _08025_);
  or _61805_ (_10168_, _10167_, _09573_);
  and _61806_ (_10169_, _10168_, _06037_);
  or _61807_ (_10170_, _10169_, _10166_);
  or _61808_ (_10171_, _10170_, _10165_);
  not _61809_ (_10172_, _10166_);
  not _61810_ (_10173_, \oc8051_golden_model_1.B [1]);
  nor _61811_ (_10174_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor _61812_ (_10175_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and _61813_ (_10176_, _10175_, _10174_);
  and _61814_ (_10177_, _10176_, _10173_);
  nor _61815_ (_10178_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not _61816_ (_10179_, \oc8051_golden_model_1.B [0]);
  and _61817_ (_10180_, _10179_, \oc8051_golden_model_1.ACC [7]);
  and _61818_ (_10181_, _10180_, _10178_);
  and _61819_ (_10182_, _10181_, _10177_);
  and _61820_ (_10183_, _10178_, _10177_);
  nor _61821_ (_10184_, _10183_, _08688_);
  or _61822_ (_10185_, _10179_, \oc8051_golden_model_1.ACC [6]);
  and _61823_ (_10186_, _10185_, \oc8051_golden_model_1.ACC [7]);
  or _61824_ (_10187_, _10186_, _10173_);
  and _61825_ (_10188_, _10178_, _10176_);
  and _61826_ (_10189_, _10188_, _10187_);
  not _61827_ (_10190_, _10189_);
  and _61828_ (_10191_, _10190_, _10184_);
  nor _61829_ (_10192_, _10191_, _10182_);
  not _61830_ (_10193_, \oc8051_golden_model_1.ACC [6]);
  and _61831_ (_10194_, _10189_, \oc8051_golden_model_1.B [0]);
  nor _61832_ (_10195_, _10194_, _10193_);
  and _61833_ (_10196_, _10195_, _10173_);
  nor _61834_ (_10197_, _10195_, _10173_);
  nor _61835_ (_10198_, _10197_, _10196_);
  nor _61836_ (_10199_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor _61837_ (_10200_, _10199_, _09832_);
  nor _61838_ (_10201_, _10200_, \oc8051_golden_model_1.ACC [4]);
  and _61839_ (_10202_, \oc8051_golden_model_1.ACC [4], _10179_);
  nor _61840_ (_10203_, _10202_, \oc8051_golden_model_1.ACC [5]);
  not _61841_ (_10204_, \oc8051_golden_model_1.ACC [4]);
  and _61842_ (_10205_, _10204_, \oc8051_golden_model_1.B [0]);
  nor _61843_ (_10206_, _10205_, _10203_);
  nor _61844_ (_10207_, _10206_, _10201_);
  not _61845_ (_10208_, _10207_);
  and _61846_ (_10209_, _10208_, _10198_);
  not _61847_ (_10210_, _10209_);
  nor _61848_ (_10211_, _10192_, \oc8051_golden_model_1.B [2]);
  nor _61849_ (_10212_, _10211_, _10196_);
  and _61850_ (_10213_, _10212_, _10210_);
  not _61851_ (_10214_, _10213_);
  not _61852_ (_10215_, \oc8051_golden_model_1.B [3]);
  nor _61853_ (_10216_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _61854_ (_10217_, _10216_, _10174_);
  and _61855_ (_10218_, _10217_, _10215_);
  and _61856_ (_10219_, \oc8051_golden_model_1.B [2], _08688_);
  not _61857_ (_10220_, _10219_);
  and _61858_ (_10221_, _10220_, _10218_);
  and _61859_ (_10222_, _10221_, _10214_);
  nor _61860_ (_10223_, _10222_, _10192_);
  nor _61861_ (_10224_, _10223_, _10182_);
  and _61862_ (_10225_, _10217_, \oc8051_golden_model_1.ACC [7]);
  nor _61863_ (_10226_, _10225_, _10218_);
  nor _61864_ (_10227_, _10224_, \oc8051_golden_model_1.B [3]);
  nor _61865_ (_10228_, _10208_, _10198_);
  nor _61866_ (_10229_, _10228_, _10209_);
  and _61867_ (_10230_, _10229_, _10222_);
  not _61868_ (_10231_, _10195_);
  nor _61869_ (_10232_, _10222_, _10231_);
  nor _61870_ (_10233_, _10232_, _10230_);
  nor _61871_ (_10234_, _10233_, \oc8051_golden_model_1.B [2]);
  and _61872_ (_10235_, _10233_, \oc8051_golden_model_1.B [2]);
  nor _61873_ (_10236_, _10235_, _10234_);
  not _61874_ (_10237_, \oc8051_golden_model_1.ACC [5]);
  nor _61875_ (_10238_, _10222_, _10237_);
  and _61876_ (_10239_, _10222_, _10200_);
  or _61877_ (_10240_, _10239_, _10238_);
  and _61878_ (_10241_, _10240_, _10173_);
  nor _61879_ (_10242_, _10240_, _10173_);
  nor _61880_ (_10243_, _10242_, _10205_);
  nor _61881_ (_10244_, _10243_, _10241_);
  not _61882_ (_10245_, _10244_);
  and _61883_ (_10246_, _10245_, _10236_);
  or _61884_ (_10247_, _10246_, _10234_);
  nor _61885_ (_10248_, _10247_, _10227_);
  nor _61886_ (_10249_, _10248_, _10226_);
  nor _61887_ (_10250_, _10249_, _10224_);
  nor _61888_ (_10251_, _10250_, _10182_);
  nor _61889_ (_10252_, _10249_, _10233_);
  nor _61890_ (_10253_, _10245_, _10236_);
  nor _61891_ (_10254_, _10253_, _10246_);
  and _61892_ (_10255_, _10254_, _10249_);
  or _61893_ (_10256_, _10255_, _10252_);
  and _61894_ (_10257_, _10256_, _10215_);
  nor _61895_ (_10258_, _10256_, _10215_);
  nor _61896_ (_10259_, _10258_, _10257_);
  not _61897_ (_10260_, _10259_);
  nor _61898_ (_10261_, _10249_, _10240_);
  nor _61899_ (_10262_, _10242_, _10241_);
  and _61900_ (_10263_, _10262_, _10205_);
  nor _61901_ (_10264_, _10262_, _10205_);
  nor _61902_ (_10265_, _10264_, _10263_);
  and _61903_ (_10266_, _10265_, _10249_);
  or _61904_ (_10267_, _10266_, _10261_);
  nor _61905_ (_10268_, _10267_, \oc8051_golden_model_1.B [2]);
  and _61906_ (_10269_, _10267_, \oc8051_golden_model_1.B [2]);
  nor _61907_ (_10270_, _10205_, _10202_);
  and _61908_ (_10271_, _10249_, _10270_);
  nor _61909_ (_10272_, _10249_, \oc8051_golden_model_1.ACC [4]);
  nor _61910_ (_10273_, _10272_, _10271_);
  and _61911_ (_10274_, _10273_, _10173_);
  nor _61912_ (_10275_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _61913_ (_10276_, _10275_, _10016_);
  nor _61914_ (_10277_, _10276_, \oc8051_golden_model_1.ACC [2]);
  and _61915_ (_10278_, _10179_, \oc8051_golden_model_1.ACC [2]);
  nor _61916_ (_10279_, _10278_, \oc8051_golden_model_1.ACC [3]);
  not _61917_ (_10280_, \oc8051_golden_model_1.ACC [2]);
  and _61918_ (_10281_, \oc8051_golden_model_1.B [0], _10280_);
  nor _61919_ (_10282_, _10281_, _10279_);
  nor _61920_ (_10283_, _10282_, _10277_);
  not _61921_ (_10284_, _10283_);
  nor _61922_ (_10285_, _10273_, _10173_);
  nor _61923_ (_10286_, _10285_, _10274_);
  and _61924_ (_10287_, _10286_, _10284_);
  nor _61925_ (_10288_, _10287_, _10274_);
  nor _61926_ (_10289_, _10288_, _10269_);
  nor _61927_ (_10290_, _10289_, _10268_);
  nor _61928_ (_10291_, _10290_, _10260_);
  nor _61929_ (_10292_, _10251_, \oc8051_golden_model_1.B [4]);
  nor _61930_ (_10293_, _10292_, _10257_);
  not _61931_ (_10294_, _10293_);
  nor _61932_ (_10295_, _10294_, _10291_);
  not _61933_ (_10296_, \oc8051_golden_model_1.B [5]);
  and _61934_ (_10297_, _10216_, _10296_);
  and _61935_ (_10298_, \oc8051_golden_model_1.B [4], _08688_);
  not _61936_ (_10299_, _10298_);
  and _61937_ (_10300_, _10299_, _10297_);
  not _61938_ (_10301_, _10300_);
  nor _61939_ (_10302_, _10301_, _10295_);
  nor _61940_ (_10303_, _10302_, _10251_);
  nor _61941_ (_10304_, _10303_, _10182_);
  not _61942_ (_10305_, \oc8051_golden_model_1.B [4]);
  and _61943_ (_10306_, _10290_, _10260_);
  nor _61944_ (_10307_, _10306_, _10291_);
  not _61945_ (_10308_, _10307_);
  and _61946_ (_10309_, _10308_, _10302_);
  nor _61947_ (_10310_, _10302_, _10256_);
  nor _61948_ (_10311_, _10310_, _10309_);
  and _61949_ (_10312_, _10311_, _10305_);
  nor _61950_ (_10313_, _10311_, _10305_);
  nor _61951_ (_10314_, _10313_, _10312_);
  not _61952_ (_10315_, _10314_);
  nor _61953_ (_10316_, _10302_, _10267_);
  nor _61954_ (_10317_, _10269_, _10268_);
  and _61955_ (_10318_, _10317_, _10288_);
  nor _61956_ (_10319_, _10317_, _10288_);
  nor _61957_ (_10320_, _10319_, _10318_);
  not _61958_ (_10321_, _10320_);
  and _61959_ (_10322_, _10321_, _10302_);
  nor _61960_ (_10323_, _10322_, _10316_);
  nor _61961_ (_10324_, _10323_, \oc8051_golden_model_1.B [3]);
  and _61962_ (_10325_, _10323_, \oc8051_golden_model_1.B [3]);
  not _61963_ (_10326_, \oc8051_golden_model_1.B [2]);
  nor _61964_ (_10327_, _10286_, _10284_);
  nor _61965_ (_10328_, _10327_, _10287_);
  not _61966_ (_10329_, _10328_);
  and _61967_ (_10330_, _10329_, _10302_);
  nor _61968_ (_10331_, _10302_, _10273_);
  nor _61969_ (_10332_, _10331_, _10330_);
  and _61970_ (_10333_, _10332_, _10326_);
  not _61971_ (_10334_, \oc8051_golden_model_1.ACC [3]);
  nor _61972_ (_10335_, _10302_, _10334_);
  and _61973_ (_10336_, _10302_, _10276_);
  or _61974_ (_10337_, _10336_, _10335_);
  and _61975_ (_10338_, _10337_, _10173_);
  nor _61976_ (_10339_, _10337_, _10173_);
  nor _61977_ (_10340_, _10339_, _10281_);
  nor _61978_ (_10341_, _10340_, _10338_);
  nor _61979_ (_10342_, _10332_, _10326_);
  nor _61980_ (_10343_, _10342_, _10333_);
  not _61981_ (_10344_, _10343_);
  nor _61982_ (_10345_, _10344_, _10341_);
  nor _61983_ (_10346_, _10345_, _10333_);
  nor _61984_ (_10347_, _10346_, _10325_);
  nor _61985_ (_10348_, _10347_, _10324_);
  nor _61986_ (_10349_, _10348_, _10315_);
  nor _61987_ (_10350_, _10304_, \oc8051_golden_model_1.B [5]);
  nor _61988_ (_10351_, _10350_, _10312_);
  not _61989_ (_10352_, _10351_);
  nor _61990_ (_10353_, _10352_, _10349_);
  not _61991_ (_10354_, _10353_);
  not _61992_ (_10355_, _10216_);
  and _61993_ (_10356_, \oc8051_golden_model_1.B [5], _08688_);
  nor _61994_ (_10357_, _10356_, _10355_);
  and _61995_ (_10358_, _10357_, _10354_);
  nor _61996_ (_10359_, _10358_, _10304_);
  not _61997_ (_10360_, _10358_);
  and _61998_ (_10361_, _10348_, _10315_);
  nor _61999_ (_10362_, _10361_, _10349_);
  nor _62000_ (_10363_, _10362_, _10360_);
  nor _62001_ (_10364_, _10358_, _10311_);
  nor _62002_ (_10365_, _10364_, _10363_);
  and _62003_ (_10366_, _10365_, _10296_);
  nor _62004_ (_10367_, _10365_, _10296_);
  nor _62005_ (_10368_, _10367_, _10366_);
  not _62006_ (_10369_, _10368_);
  nor _62007_ (_10370_, _10358_, _10323_);
  nor _62008_ (_10371_, _10325_, _10324_);
  nor _62009_ (_10372_, _10371_, _10346_);
  and _62010_ (_10373_, _10371_, _10346_);
  or _62011_ (_10374_, _10373_, _10372_);
  and _62012_ (_10375_, _10374_, _10358_);
  or _62013_ (_10376_, _10375_, _10370_);
  and _62014_ (_10377_, _10376_, _10305_);
  nor _62015_ (_10378_, _10376_, _10305_);
  and _62016_ (_10379_, _10344_, _10341_);
  nor _62017_ (_10380_, _10379_, _10345_);
  nor _62018_ (_10381_, _10380_, _10360_);
  nor _62019_ (_10382_, _10358_, _10332_);
  nor _62020_ (_10383_, _10382_, _10381_);
  and _62021_ (_10384_, _10383_, _10215_);
  nor _62022_ (_10385_, _10339_, _10338_);
  nor _62023_ (_10386_, _10385_, _10281_);
  and _62024_ (_10387_, _10385_, _10281_);
  or _62025_ (_10388_, _10387_, _10386_);
  nor _62026_ (_10389_, _10388_, _10360_);
  nor _62027_ (_10390_, _10358_, _10337_);
  nor _62028_ (_10391_, _10390_, _10389_);
  and _62029_ (_10392_, _10391_, _10326_);
  nor _62030_ (_10393_, _10391_, _10326_);
  nor _62031_ (_10394_, _10281_, _10278_);
  and _62032_ (_10395_, _10358_, _10394_);
  nor _62033_ (_10396_, _10358_, \oc8051_golden_model_1.ACC [2]);
  nor _62034_ (_10397_, _10396_, _10395_);
  and _62035_ (_10398_, _10397_, _10173_);
  and _62036_ (_10399_, _06097_, \oc8051_golden_model_1.B [0]);
  not _62037_ (_10400_, _10399_);
  nor _62038_ (_10401_, _10397_, _10173_);
  nor _62039_ (_10402_, _10401_, _10398_);
  and _62040_ (_10403_, _10402_, _10400_);
  nor _62041_ (_10404_, _10403_, _10398_);
  nor _62042_ (_10405_, _10404_, _10393_);
  nor _62043_ (_10406_, _10405_, _10392_);
  nor _62044_ (_10407_, _10383_, _10215_);
  nor _62045_ (_10408_, _10407_, _10384_);
  not _62046_ (_10409_, _10408_);
  nor _62047_ (_10410_, _10409_, _10406_);
  nor _62048_ (_10411_, _10410_, _10384_);
  nor _62049_ (_10412_, _10411_, _10378_);
  nor _62050_ (_10413_, _10412_, _10377_);
  nor _62051_ (_10414_, _10413_, _10369_);
  nor _62052_ (_10415_, _10414_, _10366_);
  and _62053_ (_10416_, \oc8051_golden_model_1.ACC [7], _09570_);
  nor _62054_ (_10417_, _10416_, _10216_);
  nor _62055_ (_10418_, _10417_, _10415_);
  nor _62056_ (_10419_, _10359_, _10182_);
  nor _62057_ (_10420_, _10419_, _10355_);
  nor _62058_ (_10421_, _10420_, _10418_);
  and _62059_ (_10422_, _10421_, _10359_);
  or _62060_ (_10423_, _10422_, _10182_);
  nor _62061_ (_10424_, _10423_, _09570_);
  and _62062_ (_10425_, _10421_, _10391_);
  nor _62063_ (_10426_, _10393_, _10392_);
  and _62064_ (_10427_, _10426_, _10404_);
  nor _62065_ (_10428_, _10426_, _10404_);
  nor _62066_ (_10429_, _10428_, _10427_);
  nor _62067_ (_10430_, _10429_, _10421_);
  or _62068_ (_10431_, _10430_, _10425_);
  and _62069_ (_10432_, _10431_, _10215_);
  nor _62070_ (_10433_, _10431_, _10215_);
  nor _62071_ (_10434_, _10433_, _10432_);
  nor _62072_ (_10435_, _10402_, _10400_);
  nor _62073_ (_10436_, _10435_, _10403_);
  nor _62074_ (_10437_, _10436_, _10421_);
  not _62075_ (_10438_, _10421_);
  nor _62076_ (_10439_, _10438_, _10397_);
  nor _62077_ (_10440_, _10439_, _10437_);
  nor _62078_ (_10441_, _10440_, _10326_);
  and _62079_ (_10442_, _10440_, _10326_);
  nor _62080_ (_10443_, _10442_, _10441_);
  and _62081_ (_10444_, _10443_, _10434_);
  and _62082_ (_10445_, _10421_, _06097_);
  nor _62083_ (_10446_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  nor _62084_ (_10447_, _10446_, _10093_);
  nor _62085_ (_10448_, _10421_, _10447_);
  nor _62086_ (_10449_, _10448_, _10445_);
  and _62087_ (_10450_, _10449_, _10173_);
  nor _62088_ (_10451_, _10449_, _10173_);
  and _62089_ (_10452_, _10179_, \oc8051_golden_model_1.ACC [0]);
  not _62090_ (_10453_, _10452_);
  nor _62091_ (_10454_, _10453_, _10451_);
  nor _62092_ (_10455_, _10454_, _10450_);
  and _62093_ (_10456_, _10455_, _10444_);
  and _62094_ (_10457_, _10441_, _10434_);
  nor _62095_ (_10458_, _10457_, _10433_);
  not _62096_ (_10459_, _10458_);
  nor _62097_ (_10460_, _10459_, _10456_);
  and _62098_ (_10461_, _10409_, _10406_);
  nor _62099_ (_10462_, _10461_, _10410_);
  nor _62100_ (_10463_, _10462_, _10421_);
  nor _62101_ (_10464_, _10438_, _10383_);
  nor _62102_ (_10465_, _10464_, _10463_);
  nor _62103_ (_10466_, _10465_, _10305_);
  and _62104_ (_10467_, _10465_, _10305_);
  nor _62105_ (_10468_, _10467_, _10466_);
  nor _62106_ (_10469_, _10378_, _10377_);
  nor _62107_ (_10470_, _10469_, _10411_);
  and _62108_ (_10471_, _10469_, _10411_);
  or _62109_ (_10472_, _10471_, _10470_);
  nor _62110_ (_10473_, _10472_, _10421_);
  nor _62111_ (_10474_, _10438_, _10376_);
  nor _62112_ (_10475_, _10474_, _10473_);
  nor _62113_ (_10476_, _10475_, _10296_);
  and _62114_ (_10477_, _10475_, _10296_);
  nor _62115_ (_10478_, _10477_, _10476_);
  and _62116_ (_10479_, _10478_, _10468_);
  nor _62117_ (_10480_, _10423_, \oc8051_golden_model_1.B [7]);
  nor _62118_ (_10481_, _10480_, _10133_);
  not _62119_ (_10482_, _10481_);
  not _62120_ (_10483_, \oc8051_golden_model_1.B [6]);
  and _62121_ (_10484_, _10413_, _10369_);
  nor _62122_ (_10485_, _10484_, _10414_);
  nor _62123_ (_10486_, _10485_, _10421_);
  nor _62124_ (_10487_, _10438_, _10365_);
  nor _62125_ (_10488_, _10487_, _10486_);
  nor _62126_ (_10489_, _10488_, _10483_);
  and _62127_ (_10490_, _10488_, _10483_);
  nor _62128_ (_10491_, _10490_, _10489_);
  and _62129_ (_10492_, _10491_, _10482_);
  and _62130_ (_10493_, _10492_, _10479_);
  not _62131_ (_10494_, _10493_);
  nor _62132_ (_10495_, _10494_, _10460_);
  not _62133_ (_10496_, _10492_);
  and _62134_ (_10497_, _10478_, _10466_);
  nor _62135_ (_10498_, _10497_, _10476_);
  nor _62136_ (_10499_, _10498_, _10496_);
  and _62137_ (_10500_, _10489_, _10482_);
  or _62138_ (_10501_, _10500_, _10499_);
  or _62139_ (_10502_, _10501_, _10495_);
  nor _62140_ (_10503_, _10502_, _10424_);
  nor _62141_ (_10504_, _10451_, _10450_);
  and _62142_ (_10505_, \oc8051_golden_model_1.B [0], _06071_);
  not _62143_ (_10506_, _10505_);
  and _62144_ (_10507_, _10506_, _10504_);
  and _62145_ (_10508_, _10507_, _10453_);
  and _62146_ (_10509_, _10508_, _10444_);
  and _62147_ (_10510_, _10509_, _10493_);
  nor _62148_ (_10511_, _10510_, _10503_);
  or _62149_ (_10512_, _10511_, _10182_);
  and _62150_ (_10513_, _10512_, _10423_);
  or _62151_ (_10514_, _10513_, _10172_);
  and _62152_ (_10515_, _10514_, _10171_);
  or _62153_ (_10516_, _10515_, _06277_);
  and _62154_ (_10517_, _08880_, _08025_);
  or _62155_ (_10518_, _10517_, _09573_);
  or _62156_ (_10519_, _10518_, _06278_);
  and _62157_ (_10520_, _10519_, _07334_);
  and _62158_ (_10521_, _10520_, _10516_);
  and _62159_ (_10522_, _09090_, _08025_);
  or _62160_ (_10523_, _10522_, _09573_);
  and _62161_ (_10524_, _10523_, _06502_);
  or _62162_ (_10525_, _10524_, _06615_);
  or _62163_ (_10526_, _10525_, _10521_);
  and _62164_ (_10527_, _09096_, _08025_);
  or _62165_ (_10528_, _09573_, _07337_);
  or _62166_ (_10529_, _10528_, _10527_);
  and _62167_ (_10530_, _10529_, _07339_);
  and _62168_ (_10531_, _10530_, _10526_);
  or _62169_ (_10532_, _09573_, _08110_);
  and _62170_ (_10533_, _10518_, _06507_);
  and _62171_ (_10534_, _10533_, _10532_);
  or _62172_ (_10535_, _10534_, _10531_);
  and _62173_ (_10536_, _10535_, _07331_);
  and _62174_ (_10537_, _09586_, _06610_);
  and _62175_ (_10538_, _10537_, _10532_);
  or _62176_ (_10539_, _10538_, _06509_);
  or _62177_ (_10540_, _10539_, _10536_);
  and _62178_ (_10541_, _09087_, _08025_);
  or _62179_ (_10542_, _09573_, _09107_);
  or _62180_ (_10543_, _10542_, _10541_);
  and _62181_ (_10544_, _10543_, _09112_);
  and _62182_ (_10545_, _10544_, _10540_);
  nor _62183_ (_10546_, _09095_, _09574_);
  or _62184_ (_10547_, _10546_, _09573_);
  and _62185_ (_10548_, _10547_, _06602_);
  or _62186_ (_10549_, _10548_, _06639_);
  or _62187_ (_10550_, _10549_, _10545_);
  or _62188_ (_10551_, _09583_, _07048_);
  and _62189_ (_10552_, _10551_, _05990_);
  and _62190_ (_10553_, _10552_, _10550_);
  and _62191_ (_10554_, _09580_, _05989_);
  or _62192_ (_10555_, _10554_, _06646_);
  or _62193_ (_10556_, _10555_, _10553_);
  and _62194_ (_10557_, _08605_, _08025_);
  or _62195_ (_10558_, _09573_, _06651_);
  or _62196_ (_10559_, _10558_, _10557_);
  and _62197_ (_10560_, _10559_, _01442_);
  and _62198_ (_10561_, _10560_, _10556_);
  or _62199_ (_10562_, _10561_, _09571_);
  and _62200_ (_41496_, _10562_, _43634_);
  nor _62201_ (_10563_, _01442_, _08688_);
  and _62202_ (_10564_, _06030_, _06360_);
  nand _62203_ (_10565_, _10564_, _10193_);
  and _62204_ (_10566_, _06489_, _06360_);
  not _62205_ (_10567_, _10566_);
  nor _62206_ (_10568_, _08211_, _10193_);
  nor _62207_ (_10569_, _08307_, _10237_);
  and _62208_ (_10570_, _08307_, _10237_);
  nor _62209_ (_10571_, _08598_, _10204_);
  not _62210_ (_10572_, _10571_);
  nor _62211_ (_10573_, _08358_, _10334_);
  and _62212_ (_10574_, _08358_, _10334_);
  nor _62213_ (_10575_, _08502_, _10280_);
  nor _62214_ (_10576_, _08403_, _06097_);
  and _62215_ (_10577_, _08453_, \oc8051_golden_model_1.ACC [0]);
  and _62216_ (_10578_, _08403_, _06097_);
  nor _62217_ (_10579_, _10578_, _10576_);
  and _62218_ (_10580_, _10579_, _10577_);
  nor _62219_ (_10581_, _10580_, _10576_);
  and _62220_ (_10582_, _08502_, _10280_);
  nor _62221_ (_10583_, _10582_, _10575_);
  not _62222_ (_10584_, _10583_);
  nor _62223_ (_10585_, _10584_, _10581_);
  nor _62224_ (_10586_, _10585_, _10575_);
  nor _62225_ (_10587_, _10586_, _10574_);
  or _62226_ (_10588_, _10587_, _10573_);
  and _62227_ (_10589_, _08598_, _10204_);
  nor _62228_ (_10590_, _10589_, _10571_);
  nand _62229_ (_10591_, _10590_, _10588_);
  and _62230_ (_10592_, _10591_, _10572_);
  nor _62231_ (_10593_, _10592_, _10570_);
  or _62232_ (_10594_, _10593_, _10569_);
  and _62233_ (_10595_, _08211_, _10193_);
  nor _62234_ (_10596_, _10595_, _10568_);
  and _62235_ (_10597_, _10596_, _10594_);
  nor _62236_ (_10598_, _10597_, _10568_);
  nor _62237_ (_10599_, _10598_, _09096_);
  and _62238_ (_10600_, _10598_, _09096_);
  or _62239_ (_10601_, _10600_, _10599_);
  and _62240_ (_10602_, _10601_, _06363_);
  nor _62241_ (_10603_, _08017_, _08688_);
  and _62242_ (_10604_, _09087_, _08017_);
  or _62243_ (_10605_, _10604_, _10603_);
  and _62244_ (_10606_, _10605_, _06509_);
  and _62245_ (_10607_, _08107_, _08688_);
  nor _62246_ (_10608_, _06318_, _07167_);
  nor _62247_ (_10609_, _10608_, _06022_);
  nand _62248_ (_10610_, _10609_, _10607_);
  not _62249_ (_10611_, _06976_);
  nor _62250_ (_10612_, _08107_, _08688_);
  nor _62251_ (_10613_, _10608_, _06017_);
  or _62252_ (_10614_, _06903_, _06480_);
  and _62253_ (_10615_, _10614_, _06506_);
  nor _62254_ (_10616_, _10615_, _10613_);
  not _62255_ (_10617_, _10616_);
  and _62256_ (_10618_, _10617_, _10612_);
  not _62257_ (_10619_, _08017_);
  nor _62258_ (_10620_, _08107_, _10619_);
  or _62259_ (_10621_, _10620_, _10603_);
  or _62260_ (_10622_, _10621_, _06327_);
  and _62261_ (_10623_, _06489_, _06038_);
  not _62262_ (_10624_, _10623_);
  and _62263_ (_10625_, _08602_, \oc8051_golden_model_1.PSW [7]);
  nor _62264_ (_10626_, _10625_, _08109_);
  and _62265_ (_10627_, _10625_, _08109_);
  nor _62266_ (_10628_, _10627_, _10626_);
  and _62267_ (_10629_, _10628_, \oc8051_golden_model_1.ACC [7]);
  nor _62268_ (_10630_, _10628_, \oc8051_golden_model_1.ACC [7]);
  nor _62269_ (_10631_, _10630_, _10629_);
  not _62270_ (_10632_, _10631_);
  and _62271_ (_10633_, _08505_, \oc8051_golden_model_1.PSW [7]);
  and _62272_ (_10634_, _10633_, _08599_);
  and _62273_ (_10635_, _10634_, _08308_);
  nor _62274_ (_10636_, _10635_, _08212_);
  nor _62275_ (_10637_, _10636_, _10625_);
  nor _62276_ (_10638_, _10637_, _10193_);
  nor _62277_ (_10639_, _10634_, _08308_);
  nor _62278_ (_10640_, _10639_, _10635_);
  and _62279_ (_10641_, _10640_, _10237_);
  nor _62280_ (_10642_, _10640_, _10237_);
  nor _62281_ (_10643_, _10633_, _08599_);
  nor _62282_ (_10644_, _10643_, _10634_);
  nor _62283_ (_10645_, _10644_, _10204_);
  nor _62284_ (_10646_, _10645_, _10642_);
  nor _62285_ (_10647_, _10646_, _10641_);
  nor _62286_ (_10648_, _10642_, _10641_);
  not _62287_ (_10649_, _10648_);
  and _62288_ (_10650_, _10644_, _10204_);
  or _62289_ (_10651_, _10650_, _10645_);
  or _62290_ (_10652_, _10651_, _10649_);
  and _62291_ (_10653_, _08504_, \oc8051_golden_model_1.PSW [7]);
  nor _62292_ (_10654_, _10653_, _08359_);
  nor _62293_ (_10655_, _10654_, _10633_);
  nor _62294_ (_10656_, _10655_, _10334_);
  and _62295_ (_10657_, _10655_, _10334_);
  nor _62296_ (_10658_, _10657_, _10656_);
  and _62297_ (_10659_, _08454_, \oc8051_golden_model_1.PSW [7]);
  nor _62298_ (_10660_, _10659_, _08503_);
  nor _62299_ (_10661_, _10660_, _10653_);
  nor _62300_ (_10662_, _10661_, _10280_);
  and _62301_ (_10663_, _10661_, _10280_);
  nor _62302_ (_10664_, _10663_, _10662_);
  and _62303_ (_10665_, _10664_, _10658_);
  and _62304_ (_10666_, _08453_, \oc8051_golden_model_1.PSW [7]);
  nor _62305_ (_10667_, _10666_, _08404_);
  nor _62306_ (_10668_, _10667_, _10659_);
  nor _62307_ (_10669_, _10668_, _06097_);
  and _62308_ (_10670_, _10668_, _06097_);
  nor _62309_ (_10671_, _08453_, \oc8051_golden_model_1.PSW [7]);
  nor _62310_ (_10672_, _10671_, _10666_);
  and _62311_ (_10673_, _10672_, _06071_);
  nor _62312_ (_10674_, _10673_, _10670_);
  or _62313_ (_10675_, _10674_, _10669_);
  nand _62314_ (_10676_, _10675_, _10665_);
  and _62315_ (_10677_, _10662_, _10658_);
  nor _62316_ (_10678_, _10677_, _10656_);
  and _62317_ (_10679_, _10678_, _10676_);
  nor _62318_ (_10680_, _10679_, _10652_);
  nor _62319_ (_10681_, _10680_, _10647_);
  and _62320_ (_10683_, _10637_, _10193_);
  nor _62321_ (_10684_, _10638_, _10683_);
  not _62322_ (_10685_, _10684_);
  nor _62323_ (_10686_, _10685_, _10681_);
  or _62324_ (_10687_, _10686_, _10638_);
  and _62325_ (_10688_, _10687_, _10632_);
  nor _62326_ (_10689_, _10687_, _10632_);
  or _62327_ (_10690_, _10689_, _10688_);
  or _62328_ (_10691_, _10690_, _06458_);
  and _62329_ (_10692_, _10691_, _10624_);
  and _62330_ (_10694_, _06489_, _06350_);
  nand _62331_ (_10695_, _10694_, _10334_);
  nor _62332_ (_10696_, _06056_, _06034_);
  nand _62333_ (_10697_, _10696_, _08107_);
  nor _62334_ (_10698_, _08645_, _08688_);
  and _62335_ (_10699_, _08672_, _08645_);
  or _62336_ (_10700_, _10699_, _10698_);
  or _62337_ (_10701_, _10700_, _06357_);
  and _62338_ (_10702_, _10701_, _06772_);
  and _62339_ (_10703_, _06489_, _06815_);
  and _62340_ (_10705_, _10703_, _08778_);
  and _62341_ (_10706_, _06035_, _07583_);
  not _62342_ (_10707_, _10706_);
  nor _62343_ (_10708_, _06850_, _06315_);
  and _62344_ (_10709_, _10708_, _07545_);
  and _62345_ (_10710_, _10709_, _10707_);
  nor _62346_ (_10711_, _10710_, _06061_);
  not _62347_ (_10712_, _10711_);
  nor _62348_ (_10713_, _10712_, _08107_);
  nor _62349_ (_10714_, _10711_, _10703_);
  nor _62350_ (_10716_, _06855_, _08688_);
  and _62351_ (_10717_, _06855_, _08688_);
  or _62352_ (_10718_, _10717_, _10716_);
  and _62353_ (_10719_, _10718_, _10714_);
  or _62354_ (_10720_, _10719_, _10713_);
  or _62355_ (_10721_, _10720_, _10705_);
  and _62356_ (_10722_, _07275_, _06062_);
  and _62357_ (_10723_, _10722_, _10721_);
  and _62358_ (_10724_, _08791_, _08017_);
  or _62359_ (_10725_, _10724_, _10603_);
  and _62360_ (_10727_, _10725_, _06474_);
  or _62361_ (_10728_, _10727_, _10723_);
  and _62362_ (_10729_, _06489_, _06355_);
  not _62363_ (_10730_, _10729_);
  and _62364_ (_10731_, _10730_, _10728_);
  nor _62365_ (_10732_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor _62366_ (_10733_, _10732_, _10334_);
  and _62367_ (_10734_, _10733_, \oc8051_golden_model_1.ACC [4]);
  and _62368_ (_10735_, _10734_, \oc8051_golden_model_1.ACC [5]);
  and _62369_ (_10736_, _10735_, \oc8051_golden_model_1.ACC [6]);
  and _62370_ (_10738_, _10736_, \oc8051_golden_model_1.ACC [7]);
  nor _62371_ (_10739_, _10736_, \oc8051_golden_model_1.ACC [7]);
  nor _62372_ (_10740_, _10739_, _10738_);
  nor _62373_ (_10741_, _10734_, \oc8051_golden_model_1.ACC [5]);
  nor _62374_ (_10742_, _10741_, _10735_);
  nor _62375_ (_10743_, _10735_, \oc8051_golden_model_1.ACC [6]);
  nor _62376_ (_10744_, _10743_, _10736_);
  nor _62377_ (_10745_, _10744_, _10742_);
  not _62378_ (_10746_, _10745_);
  nand _62379_ (_10747_, _10746_, _10740_);
  nor _62380_ (_10749_, _10738_, \oc8051_golden_model_1.PSW [7]);
  and _62381_ (_10750_, _10749_, _10747_);
  nor _62382_ (_10751_, _10750_, _10745_);
  or _62383_ (_10752_, _10751_, _10740_);
  and _62384_ (_10753_, _10747_, _10729_);
  and _62385_ (_10754_, _10753_, _10752_);
  or _62386_ (_10755_, _10754_, _06356_);
  or _62387_ (_10756_, _10755_, _10731_);
  and _62388_ (_10757_, _10756_, _10702_);
  and _62389_ (_10758_, _10621_, _06410_);
  or _62390_ (_10759_, _10758_, _10696_);
  or _62391_ (_10760_, _10759_, _10757_);
  and _62392_ (_10761_, _10760_, _10697_);
  or _62393_ (_10762_, _10761_, _07289_);
  or _62394_ (_10763_, _08778_, _07290_);
  and _62395_ (_10764_, _10763_, _06426_);
  and _62396_ (_10765_, _10764_, _10762_);
  nor _62397_ (_10766_, _08109_, _06426_);
  or _62398_ (_10767_, _10766_, _10694_);
  or _62399_ (_10768_, _10767_, _10765_);
  and _62400_ (_10769_, _10768_, _10695_);
  or _62401_ (_10770_, _10769_, _06352_);
  and _62402_ (_10771_, _08668_, _08645_);
  or _62403_ (_10772_, _10771_, _10698_);
  or _62404_ (_10773_, _10772_, _06353_);
  and _62405_ (_10774_, _10773_, _06346_);
  and _62406_ (_10775_, _10774_, _10770_);
  or _62407_ (_10776_, _10698_, _08809_);
  and _62408_ (_10777_, _10700_, _06345_);
  and _62409_ (_10778_, _10777_, _10776_);
  or _62410_ (_10779_, _10778_, _09606_);
  or _62411_ (_10780_, _10779_, _10775_);
  nor _62412_ (_10781_, _10112_, _10110_);
  nor _62413_ (_10782_, _10781_, _10113_);
  or _62414_ (_10783_, _10782_, _09612_);
  nand _62415_ (_10784_, _06038_, _05985_);
  and _62416_ (_10785_, _10784_, _10783_);
  and _62417_ (_10786_, _10785_, _10780_);
  and _62418_ (_10787_, _07250_, \oc8051_golden_model_1.PSW [7]);
  and _62419_ (_10788_, _10787_, _09482_);
  and _62420_ (_10789_, _10788_, _09481_);
  and _62421_ (_10790_, _10789_, _09480_);
  and _62422_ (_10791_, _10790_, _09479_);
  and _62423_ (_10792_, _10791_, _09478_);
  and _62424_ (_10793_, _10792_, _09477_);
  and _62425_ (_10794_, _10793_, _08674_);
  nor _62426_ (_10795_, _10793_, _08674_);
  or _62427_ (_10796_, _10795_, _10794_);
  and _62428_ (_10797_, _10796_, \oc8051_golden_model_1.ACC [7]);
  nor _62429_ (_10798_, _10796_, \oc8051_golden_model_1.ACC [7]);
  nor _62430_ (_10799_, _10798_, _10797_);
  not _62431_ (_10800_, _10799_);
  nor _62432_ (_10801_, _10792_, _09477_);
  nor _62433_ (_10802_, _10801_, _10793_);
  nor _62434_ (_10803_, _10802_, _10193_);
  nor _62435_ (_10804_, _10791_, _09478_);
  nor _62436_ (_10805_, _10804_, _10792_);
  and _62437_ (_10806_, _10805_, _10237_);
  nor _62438_ (_10807_, _10805_, _10237_);
  nor _62439_ (_10808_, _10790_, _09479_);
  nor _62440_ (_10809_, _10808_, _10791_);
  nor _62441_ (_10810_, _10809_, _10204_);
  nor _62442_ (_10811_, _10810_, _10807_);
  nor _62443_ (_10812_, _10811_, _10806_);
  nor _62444_ (_10813_, _10807_, _10806_);
  not _62445_ (_10814_, _10813_);
  and _62446_ (_10815_, _10809_, _10204_);
  or _62447_ (_10816_, _10815_, _10810_);
  or _62448_ (_10817_, _10816_, _10814_);
  nor _62449_ (_10818_, _10789_, _09480_);
  nor _62450_ (_10819_, _10818_, _10790_);
  nor _62451_ (_10820_, _10819_, _10334_);
  and _62452_ (_10821_, _10819_, _10334_);
  nor _62453_ (_10822_, _10821_, _10820_);
  nor _62454_ (_10823_, _10788_, _09481_);
  nor _62455_ (_10824_, _10823_, _10789_);
  nor _62456_ (_10825_, _10824_, _10280_);
  and _62457_ (_10826_, _10824_, _10280_);
  nor _62458_ (_10827_, _10826_, _10825_);
  and _62459_ (_10828_, _10827_, _10822_);
  nor _62460_ (_10829_, _10787_, _09482_);
  nor _62461_ (_10830_, _10829_, _10788_);
  nor _62462_ (_10831_, _10830_, _06097_);
  and _62463_ (_10832_, _10830_, _06097_);
  nor _62464_ (_10833_, _07250_, \oc8051_golden_model_1.PSW [7]);
  nor _62465_ (_10834_, _10833_, _10787_);
  and _62466_ (_10835_, _10834_, _06071_);
  nor _62467_ (_10836_, _10835_, _10832_);
  or _62468_ (_10837_, _10836_, _10831_);
  and _62469_ (_10838_, _10837_, _10828_);
  and _62470_ (_10839_, _10825_, _10822_);
  or _62471_ (_10840_, _10839_, _10820_);
  nor _62472_ (_10841_, _10840_, _10838_);
  nor _62473_ (_10842_, _10841_, _10817_);
  nor _62474_ (_10843_, _10842_, _10812_);
  and _62475_ (_10844_, _10802_, _10193_);
  nor _62476_ (_10845_, _10803_, _10844_);
  not _62477_ (_10846_, _10845_);
  nor _62478_ (_10847_, _10846_, _10843_);
  or _62479_ (_10848_, _10847_, _10803_);
  and _62480_ (_10849_, _10848_, _10800_);
  nor _62481_ (_10850_, _10848_, _10800_);
  nor _62482_ (_10851_, _10850_, _10849_);
  or _62483_ (_10852_, _10851_, _10784_);
  and _62484_ (_10853_, _06471_, _06038_);
  not _62485_ (_10854_, _10853_);
  nand _62486_ (_10855_, _10854_, _10852_);
  or _62487_ (_10856_, _10855_, _10786_);
  and _62488_ (_10857_, _09502_, \oc8051_golden_model_1.PSW [7]);
  nor _62489_ (_10858_, _10857_, _09496_);
  and _62490_ (_10859_, _10857_, _09496_);
  nor _62491_ (_10860_, _10859_, _10858_);
  and _62492_ (_10861_, _10860_, \oc8051_golden_model_1.ACC [7]);
  nor _62493_ (_10862_, _10860_, \oc8051_golden_model_1.ACC [7]);
  nor _62494_ (_10863_, _10862_, _10861_);
  not _62495_ (_10864_, _10863_);
  and _62496_ (_10865_, _09501_, \oc8051_golden_model_1.PSW [7]);
  nor _62497_ (_10866_, _10865_, _09172_);
  nor _62498_ (_10867_, _10866_, _10857_);
  nor _62499_ (_10868_, _10867_, _10193_);
  and _62500_ (_10869_, _09500_, \oc8051_golden_model_1.PSW [7]);
  nor _62501_ (_10870_, _10869_, _09218_);
  nor _62502_ (_10871_, _10870_, _10865_);
  and _62503_ (_10872_, _10871_, _10237_);
  nor _62504_ (_10873_, _10871_, _10237_);
  nor _62505_ (_10874_, _10873_, _10872_);
  not _62506_ (_10875_, _10874_);
  and _62507_ (_10876_, _09499_, \oc8051_golden_model_1.PSW [7]);
  nor _62508_ (_10877_, _10876_, _09264_);
  nor _62509_ (_10878_, _10877_, _10869_);
  nor _62510_ (_10879_, _10878_, _10204_);
  and _62511_ (_10880_, _10878_, _10204_);
  or _62512_ (_10881_, _10880_, _10879_);
  or _62513_ (_10882_, _10881_, _10875_);
  and _62514_ (_10883_, _09498_, \oc8051_golden_model_1.PSW [7]);
  nor _62515_ (_10884_, _10883_, _09310_);
  nor _62516_ (_10885_, _10884_, _10876_);
  nor _62517_ (_10886_, _10885_, _10334_);
  and _62518_ (_10887_, _10885_, _10334_);
  nor _62519_ (_10888_, _10887_, _10886_);
  and _62520_ (_10889_, _09497_, \oc8051_golden_model_1.PSW [7]);
  nor _62521_ (_10890_, _10889_, _09356_);
  nor _62522_ (_10891_, _10890_, _10883_);
  nor _62523_ (_10892_, _10891_, _10280_);
  and _62524_ (_10893_, _10891_, _10280_);
  nor _62525_ (_10894_, _10893_, _10892_);
  and _62526_ (_10895_, _10894_, _10888_);
  and _62527_ (_10896_, _09447_, \oc8051_golden_model_1.PSW [7]);
  nor _62528_ (_10897_, _10896_, _09402_);
  nor _62529_ (_10898_, _10897_, _10889_);
  nor _62530_ (_10899_, _10898_, _06097_);
  and _62531_ (_10900_, _10898_, _06097_);
  nor _62532_ (_10901_, _09447_, \oc8051_golden_model_1.PSW [7]);
  nor _62533_ (_10902_, _10901_, _10896_);
  and _62534_ (_10903_, _10902_, _06071_);
  nor _62535_ (_10904_, _10903_, _10900_);
  or _62536_ (_10905_, _10904_, _10899_);
  nand _62537_ (_10906_, _10905_, _10895_);
  and _62538_ (_10907_, _10892_, _10888_);
  nor _62539_ (_10908_, _10907_, _10886_);
  and _62540_ (_10909_, _10908_, _10906_);
  nor _62541_ (_10910_, _10909_, _10882_);
  and _62542_ (_10911_, _10879_, _10874_);
  nor _62543_ (_10912_, _10911_, _10873_);
  not _62544_ (_10913_, _10912_);
  nor _62545_ (_10914_, _10913_, _10910_);
  and _62546_ (_10915_, _10867_, _10193_);
  nor _62547_ (_10916_, _10868_, _10915_);
  not _62548_ (_10917_, _10916_);
  nor _62549_ (_10918_, _10917_, _10914_);
  or _62550_ (_10919_, _10918_, _10868_);
  and _62551_ (_10920_, _10919_, _10864_);
  nor _62552_ (_10921_, _10919_, _10864_);
  nor _62553_ (_10922_, _10921_, _10920_);
  nand _62554_ (_10923_, _10922_, _10853_);
  and _62555_ (_10924_, _10923_, _10856_);
  or _62556_ (_10925_, _10924_, _06453_);
  and _62557_ (_10926_, _10925_, _10692_);
  and _62558_ (_10927_, _08827_, _06622_);
  and _62559_ (_10928_, _10927_, _08020_);
  and _62560_ (_10929_, _10928_, _07741_);
  nor _62561_ (_10930_, _10929_, _06366_);
  and _62562_ (_10931_, _10929_, _06366_);
  nor _62563_ (_10932_, _10931_, _10930_);
  and _62564_ (_10933_, _10932_, \oc8051_golden_model_1.ACC [7]);
  nor _62565_ (_10934_, _10932_, \oc8051_golden_model_1.ACC [7]);
  nor _62566_ (_10935_, _10934_, _10933_);
  not _62567_ (_10936_, _10935_);
  nor _62568_ (_10937_, _10928_, _07741_);
  nor _62569_ (_10938_, _10937_, _10929_);
  nor _62570_ (_10939_, _10938_, _10193_);
  and _62571_ (_10940_, _10927_, _07959_);
  nor _62572_ (_10941_, _10940_, _07983_);
  nor _62573_ (_10942_, _10941_, _10928_);
  and _62574_ (_10943_, _10942_, _10237_);
  nor _62575_ (_10944_, _10942_, _10237_);
  nor _62576_ (_10945_, _10927_, _07959_);
  nor _62577_ (_10946_, _10945_, _10940_);
  nor _62578_ (_10947_, _10946_, _10204_);
  nor _62579_ (_10948_, _10947_, _10944_);
  nor _62580_ (_10949_, _10948_, _10943_);
  nor _62581_ (_10950_, _10944_, _10943_);
  and _62582_ (_10951_, _10946_, _10204_);
  nor _62583_ (_10952_, _10951_, _10947_);
  and _62584_ (_10953_, _10952_, _10950_);
  not _62585_ (_10954_, _10953_);
  nor _62586_ (_10955_, _08827_, _06622_);
  nor _62587_ (_10956_, _10955_, _10927_);
  and _62588_ (_10957_, _10956_, _10334_);
  nor _62589_ (_10958_, _10956_, _10334_);
  nor _62590_ (_10959_, _10958_, _10957_);
  and _62591_ (_10960_, _07990_, \oc8051_golden_model_1.PSW [7]);
  nor _62592_ (_10961_, _10960_, _07799_);
  nor _62593_ (_10962_, _10961_, _08827_);
  nor _62594_ (_10963_, _10962_, _10280_);
  and _62595_ (_10964_, _10962_, _10280_);
  nor _62596_ (_10965_, _10964_, _10963_);
  and _62597_ (_10966_, _10965_, _10959_);
  not _62598_ (_10967_, \oc8051_golden_model_1.PSW [7]);
  nor _62599_ (_10968_, _06310_, _10967_);
  nor _62600_ (_10969_, _10968_, _07383_);
  nor _62601_ (_10970_, _10969_, _10960_);
  nor _62602_ (_10971_, _10970_, _06097_);
  and _62603_ (_10972_, _10970_, _06097_);
  nor _62604_ (_10973_, _10972_, _10971_);
  not _62605_ (_10974_, _10973_);
  nor _62606_ (_10975_, _06310_, \oc8051_golden_model_1.PSW [7]);
  and _62607_ (_10976_, _06310_, \oc8051_golden_model_1.PSW [7]);
  nor _62608_ (_10977_, _10976_, _10975_);
  nor _62609_ (_10978_, _10977_, \oc8051_golden_model_1.ACC [0]);
  nor _62610_ (_10979_, _10978_, _10974_);
  or _62611_ (_10980_, _10979_, _10971_);
  and _62612_ (_10981_, _10980_, _10966_);
  not _62613_ (_10982_, _10981_);
  not _62614_ (_10983_, _10963_);
  nor _62615_ (_10984_, _10983_, _10957_);
  nor _62616_ (_10985_, _10984_, _10958_);
  and _62617_ (_10986_, _10985_, _10982_);
  nor _62618_ (_10987_, _10986_, _10954_);
  nor _62619_ (_10988_, _10987_, _10949_);
  and _62620_ (_10989_, _10938_, _10193_);
  nor _62621_ (_10990_, _10939_, _10989_);
  not _62622_ (_10991_, _10990_);
  nor _62623_ (_10992_, _10991_, _10988_);
  or _62624_ (_10993_, _10992_, _10939_);
  and _62625_ (_10994_, _10993_, _10936_);
  nor _62626_ (_10995_, _10993_, _10936_);
  or _62627_ (_10996_, _10995_, _10994_);
  and _62628_ (_10997_, _10996_, _10623_);
  or _62629_ (_10998_, _10997_, _06042_);
  or _62630_ (_10999_, _10998_, _10926_);
  or _62631_ (_11000_, _06238_, _06043_);
  and _62632_ (_11001_, _11000_, _06340_);
  and _62633_ (_11002_, _11001_, _10999_);
  and _62634_ (_11003_, _08828_, _08645_);
  or _62635_ (_11004_, _11003_, _10698_);
  and _62636_ (_11005_, _11004_, _06339_);
  or _62637_ (_11006_, _11005_, _10153_);
  or _62638_ (_11007_, _11006_, _11002_);
  and _62639_ (_11008_, _11007_, _10622_);
  or _62640_ (_11009_, _11008_, _09572_);
  and _62641_ (_11010_, _08778_, _08017_);
  or _62642_ (_11011_, _10603_, _06333_);
  or _62643_ (_11012_, _11011_, _11010_);
  and _62644_ (_11013_, _11012_, _06313_);
  and _62645_ (_11014_, _11013_, _11009_);
  and _62646_ (_11015_, _09076_, _08017_);
  or _62647_ (_11016_, _11015_, _10603_);
  and _62648_ (_11017_, _11016_, _06037_);
  or _62649_ (_11018_, _11017_, _10166_);
  or _62650_ (_11019_, _11018_, _11014_);
  or _62651_ (_11020_, _10179_, \oc8051_golden_model_1.ACC [7]);
  nand _62652_ (_11021_, _11020_, _10183_);
  nand _62653_ (_11022_, _11021_, _10166_);
  and _62654_ (_11023_, _11022_, _11019_);
  or _62655_ (_11024_, _11023_, _06031_);
  or _62656_ (_11025_, _06238_, _06032_);
  and _62657_ (_11026_, _11025_, _11024_);
  or _62658_ (_11027_, _11026_, _06277_);
  and _62659_ (_11028_, _06489_, _06276_);
  not _62660_ (_11029_, _11028_);
  and _62661_ (_11030_, _08880_, _08017_);
  or _62662_ (_11031_, _11030_, _10603_);
  or _62663_ (_11032_, _11031_, _06278_);
  and _62664_ (_11033_, _11032_, _11029_);
  and _62665_ (_11034_, _11033_, _11027_);
  and _62666_ (_11035_, _11028_, _06238_);
  nor _62667_ (_11036_, _06320_, _06011_);
  or _62668_ (_11037_, _11036_, _11035_);
  or _62669_ (_11038_, _11037_, _11034_);
  nor _62670_ (_11039_, _10612_, _10607_);
  not _62671_ (_11040_, _11036_);
  or _62672_ (_11041_, _11040_, _11039_);
  and _62673_ (_11042_, _06315_, _06501_);
  not _62674_ (_11043_, _11042_);
  not _62675_ (_11044_, _06802_);
  and _62676_ (_11045_, _06903_, _06501_);
  and _62677_ (_11046_, _07167_, _06501_);
  nor _62678_ (_11047_, _11046_, _11045_);
  and _62679_ (_11048_, _11047_, _11044_);
  and _62680_ (_11049_, _11048_, _11043_);
  and _62681_ (_11050_, _11049_, _11041_);
  and _62682_ (_11051_, _11050_, _11038_);
  and _62683_ (_11052_, _06471_, _06501_);
  not _62684_ (_11053_, _11049_);
  and _62685_ (_11054_, _11053_, _11039_);
  or _62686_ (_11055_, _11054_, _11052_);
  or _62687_ (_11056_, _11055_, _11051_);
  nor _62688_ (_11057_, _08778_, \oc8051_golden_model_1.ACC [7]);
  and _62689_ (_11058_, _08778_, \oc8051_golden_model_1.ACC [7]);
  nor _62690_ (_11059_, _11058_, _11057_);
  not _62691_ (_11060_, _11052_);
  or _62692_ (_11061_, _11060_, _11059_);
  and _62693_ (_11062_, _11061_, _06614_);
  and _62694_ (_11063_, _11062_, _11056_);
  and _62695_ (_11064_, _06489_, _06501_);
  and _62696_ (_11065_, _09096_, _06613_);
  or _62697_ (_11066_, _11065_, _11064_);
  or _62698_ (_11067_, _11066_, _11063_);
  nor _62699_ (_11068_, _06238_, \oc8051_golden_model_1.ACC [7]);
  and _62700_ (_11069_, _06238_, \oc8051_golden_model_1.ACC [7]);
  nor _62701_ (_11070_, _11069_, _11068_);
  not _62702_ (_11071_, _11064_);
  or _62703_ (_11072_, _11071_, _11070_);
  nand _62704_ (_11073_, _11072_, _11067_);
  nand _62705_ (_11074_, _11073_, _06616_);
  and _62706_ (_11075_, _09090_, _08017_);
  or _62707_ (_11076_, _11075_, _07334_);
  and _62708_ (_11077_, _11076_, _07337_);
  or _62709_ (_11078_, _11077_, _10603_);
  and _62710_ (_11079_, _11078_, _10616_);
  and _62711_ (_11080_, _11079_, _11074_);
  or _62712_ (_11081_, _11080_, _10618_);
  and _62713_ (_11082_, _11081_, _06973_);
  and _62714_ (_11083_, _10612_, _06972_);
  or _62715_ (_11084_, _11083_, _11082_);
  and _62716_ (_11085_, _11084_, _10611_);
  and _62717_ (_11086_, _11058_, _06976_);
  or _62718_ (_11087_, _11086_, _06608_);
  or _62719_ (_11088_, _11087_, _11085_);
  and _62720_ (_11089_, _06489_, _06506_);
  not _62721_ (_11090_, _11089_);
  or _62722_ (_11091_, _09094_, _06609_);
  and _62723_ (_11092_, _11091_, _11090_);
  and _62724_ (_11093_, _11092_, _11088_);
  and _62725_ (_11094_, _11089_, _11069_);
  or _62726_ (_11095_, _11094_, _11093_);
  and _62727_ (_11096_, _11095_, _07339_);
  nand _62728_ (_11097_, _11031_, _06507_);
  nor _62729_ (_11098_, _11097_, _09095_);
  or _62730_ (_11099_, _11098_, _10609_);
  or _62731_ (_11100_, _11099_, _11096_);
  and _62732_ (_11101_, _11100_, _10610_);
  and _62733_ (_11102_, _10614_, _06508_);
  or _62734_ (_11103_, _11102_, _11101_);
  or _62735_ (_11104_, _10708_, _06022_);
  nor _62736_ (_11105_, _10607_, _06984_);
  or _62737_ (_11106_, _11105_, _11104_);
  and _62738_ (_11107_, _11106_, _11103_);
  nor _62739_ (_11108_, _10607_, _06985_);
  or _62740_ (_11109_, _11108_, _06987_);
  or _62741_ (_11110_, _11109_, _11107_);
  nand _62742_ (_11111_, _11057_, _06987_);
  and _62743_ (_11112_, _11111_, _06605_);
  and _62744_ (_11113_, _11112_, _11110_);
  and _62745_ (_11114_, _06489_, _06508_);
  nor _62746_ (_11115_, _09095_, _06605_);
  or _62747_ (_11116_, _11115_, _11114_);
  or _62748_ (_11117_, _11116_, _11113_);
  nand _62749_ (_11118_, _11114_, _11068_);
  and _62750_ (_11119_, _11118_, _09107_);
  and _62751_ (_11120_, _11119_, _11117_);
  or _62752_ (_11121_, _11120_, _10606_);
  nor _62753_ (_11122_, _06320_, _06015_);
  not _62754_ (_11123_, _11122_);
  and _62755_ (_11124_, _06315_, _06511_);
  nor _62756_ (_11125_, _06324_, _06015_);
  nor _62757_ (_11126_, _11125_, _11124_);
  and _62758_ (_11127_, _11126_, _11123_);
  and _62759_ (_11128_, _11127_, _11121_);
  and _62760_ (_11129_, _06471_, _06511_);
  not _62761_ (_11130_, _11127_);
  and _62762_ (_11131_, _10802_, \oc8051_golden_model_1.ACC [6]);
  and _62763_ (_11132_, _10805_, \oc8051_golden_model_1.ACC [5]);
  nand _62764_ (_11133_, _10809_, \oc8051_golden_model_1.ACC [4]);
  and _62765_ (_11134_, _10819_, \oc8051_golden_model_1.ACC [3]);
  and _62766_ (_11135_, _10824_, \oc8051_golden_model_1.ACC [2]);
  and _62767_ (_11136_, _10830_, \oc8051_golden_model_1.ACC [1]);
  nor _62768_ (_11137_, _10832_, _10831_);
  not _62769_ (_11138_, _11137_);
  and _62770_ (_11139_, _10834_, \oc8051_golden_model_1.ACC [0]);
  and _62771_ (_11140_, _11139_, _11138_);
  nor _62772_ (_11141_, _11140_, _11136_);
  nor _62773_ (_11142_, _11141_, _10827_);
  nor _62774_ (_11143_, _11142_, _11135_);
  nor _62775_ (_11144_, _11143_, _10822_);
  or _62776_ (_11145_, _11144_, _11134_);
  nand _62777_ (_11146_, _11145_, _10816_);
  and _62778_ (_11147_, _11146_, _11133_);
  nor _62779_ (_11148_, _11147_, _10813_);
  or _62780_ (_11149_, _11148_, _11132_);
  and _62781_ (_11150_, _11149_, _10846_);
  nor _62782_ (_11151_, _11150_, _11131_);
  nor _62783_ (_11152_, _11151_, _10799_);
  and _62784_ (_11153_, _11151_, _10799_);
  nor _62785_ (_11154_, _11153_, _11152_);
  and _62786_ (_11155_, _11154_, _11130_);
  or _62787_ (_11156_, _11155_, _11129_);
  or _62788_ (_11157_, _11156_, _11128_);
  not _62789_ (_11158_, _11129_);
  nand _62790_ (_11159_, _10867_, \oc8051_golden_model_1.ACC [6]);
  and _62791_ (_11160_, _10871_, \oc8051_golden_model_1.ACC [5]);
  nand _62792_ (_11161_, _10878_, \oc8051_golden_model_1.ACC [4]);
  and _62793_ (_11162_, _10885_, \oc8051_golden_model_1.ACC [3]);
  and _62794_ (_11163_, _10891_, \oc8051_golden_model_1.ACC [2]);
  and _62795_ (_11164_, _10898_, \oc8051_golden_model_1.ACC [1]);
  nor _62796_ (_11165_, _10900_, _10899_);
  not _62797_ (_11166_, _11165_);
  and _62798_ (_11167_, _10902_, \oc8051_golden_model_1.ACC [0]);
  and _62799_ (_11168_, _11167_, _11166_);
  nor _62800_ (_11169_, _11168_, _11164_);
  nor _62801_ (_11170_, _11169_, _10894_);
  nor _62802_ (_11171_, _11170_, _11163_);
  nor _62803_ (_11172_, _11171_, _10888_);
  or _62804_ (_11173_, _11172_, _11162_);
  nand _62805_ (_11174_, _11173_, _10881_);
  and _62806_ (_11175_, _11174_, _11161_);
  nor _62807_ (_11176_, _11175_, _10874_);
  or _62808_ (_11177_, _11176_, _11160_);
  nand _62809_ (_11178_, _11177_, _10917_);
  and _62810_ (_11179_, _11178_, _11159_);
  nor _62811_ (_11180_, _11179_, _10863_);
  and _62812_ (_11181_, _11179_, _10863_);
  nor _62813_ (_11182_, _11181_, _11180_);
  or _62814_ (_11183_, _11182_, _11158_);
  and _62815_ (_11184_, _11183_, _06601_);
  and _62816_ (_11185_, _11184_, _11157_);
  and _62817_ (_11186_, _06489_, _06511_);
  nor _62818_ (_11187_, _11186_, _06600_);
  not _62819_ (_11188_, _11187_);
  nand _62820_ (_11189_, _10637_, \oc8051_golden_model_1.ACC [6]);
  and _62821_ (_11190_, _10640_, \oc8051_golden_model_1.ACC [5]);
  nand _62822_ (_11191_, _10644_, \oc8051_golden_model_1.ACC [4]);
  and _62823_ (_11192_, _10655_, \oc8051_golden_model_1.ACC [3]);
  and _62824_ (_11193_, _10661_, \oc8051_golden_model_1.ACC [2]);
  and _62825_ (_11194_, _10668_, \oc8051_golden_model_1.ACC [1]);
  nor _62826_ (_11195_, _10670_, _10669_);
  not _62827_ (_11196_, _11195_);
  and _62828_ (_11197_, _10672_, \oc8051_golden_model_1.ACC [0]);
  and _62829_ (_11198_, _11197_, _11196_);
  nor _62830_ (_11199_, _11198_, _11194_);
  nor _62831_ (_11200_, _11199_, _10664_);
  nor _62832_ (_11201_, _11200_, _11193_);
  nor _62833_ (_11202_, _11201_, _10658_);
  or _62834_ (_11203_, _11202_, _11192_);
  nand _62835_ (_11204_, _11203_, _10651_);
  and _62836_ (_11205_, _11204_, _11191_);
  nor _62837_ (_11206_, _11205_, _10648_);
  or _62838_ (_11207_, _11206_, _11190_);
  nand _62839_ (_11208_, _11207_, _10685_);
  and _62840_ (_11209_, _11208_, _11189_);
  nor _62841_ (_11210_, _11209_, _10631_);
  and _62842_ (_11211_, _11209_, _10631_);
  nor _62843_ (_11212_, _11211_, _11210_);
  or _62844_ (_11213_, _11212_, _11186_);
  and _62845_ (_11214_, _11213_, _11188_);
  or _62846_ (_11215_, _11214_, _11185_);
  and _62847_ (_11216_, _06030_, _06511_);
  not _62848_ (_11217_, _11216_);
  not _62849_ (_11218_, _11186_);
  nand _62850_ (_11219_, _10938_, \oc8051_golden_model_1.ACC [6]);
  and _62851_ (_11220_, _10942_, \oc8051_golden_model_1.ACC [5]);
  nand _62852_ (_11221_, _10946_, \oc8051_golden_model_1.ACC [4]);
  not _62853_ (_11222_, _10952_);
  and _62854_ (_11223_, _10956_, \oc8051_golden_model_1.ACC [3]);
  and _62855_ (_11224_, _10962_, \oc8051_golden_model_1.ACC [2]);
  and _62856_ (_11225_, _10970_, \oc8051_golden_model_1.ACC [1]);
  nor _62857_ (_11226_, _10977_, _06071_);
  and _62858_ (_11227_, _11226_, _10974_);
  nor _62859_ (_11228_, _11227_, _11225_);
  nor _62860_ (_11229_, _11228_, _10965_);
  nor _62861_ (_11230_, _11229_, _11224_);
  nor _62862_ (_11231_, _11230_, _10959_);
  or _62863_ (_11232_, _11231_, _11223_);
  nand _62864_ (_11233_, _11232_, _11222_);
  and _62865_ (_11234_, _11233_, _11221_);
  nor _62866_ (_11235_, _11234_, _10950_);
  or _62867_ (_11236_, _11235_, _11220_);
  nand _62868_ (_11237_, _11236_, _10991_);
  and _62869_ (_11238_, _11237_, _11219_);
  nor _62870_ (_11239_, _11238_, _10935_);
  and _62871_ (_11240_, _11238_, _10935_);
  nor _62872_ (_11241_, _11240_, _11239_);
  or _62873_ (_11242_, _11241_, _11218_);
  and _62874_ (_11243_, _11242_, _11217_);
  and _62875_ (_11244_, _11243_, _11215_);
  nand _62876_ (_11245_, _11216_, \oc8051_golden_model_1.ACC [6]);
  nor _62877_ (_11246_, _10608_, _06020_);
  nor _62878_ (_11247_, _10708_, _06020_);
  nor _62879_ (_11248_, _11247_, _11246_);
  nand _62880_ (_11249_, _11248_, _11245_);
  or _62881_ (_11250_, _11249_, _11244_);
  nor _62882_ (_11251_, _08209_, _10193_);
  not _62883_ (_11252_, _11251_);
  nand _62884_ (_11253_, _08209_, _10193_);
  and _62885_ (_11254_, _11253_, _11252_);
  nor _62886_ (_11255_, _08305_, _10237_);
  and _62887_ (_11256_, _08305_, _10237_);
  nor _62888_ (_11257_, _11256_, _11255_);
  nor _62889_ (_11258_, _08596_, _10204_);
  not _62890_ (_11259_, _11258_);
  nand _62891_ (_11260_, _08596_, _10204_);
  and _62892_ (_11261_, _11260_, _11259_);
  nor _62893_ (_11262_, _07680_, _10334_);
  and _62894_ (_11263_, _07680_, _10334_);
  nor _62895_ (_11264_, _07854_, _10280_);
  and _62896_ (_11265_, _07854_, _10280_);
  nor _62897_ (_11266_, _11265_, _11264_);
  not _62898_ (_11267_, _11266_);
  nor _62899_ (_11268_, _07448_, _06097_);
  and _62900_ (_11269_, _07448_, _06097_);
  nor _62901_ (_11270_, _11269_, _11268_);
  and _62902_ (_11271_, _07250_, \oc8051_golden_model_1.ACC [0]);
  and _62903_ (_11272_, _11271_, _11270_);
  nor _62904_ (_11273_, _11272_, _11268_);
  nor _62905_ (_11274_, _11273_, _11267_);
  nor _62906_ (_11275_, _11274_, _11264_);
  nor _62907_ (_11276_, _11275_, _11263_);
  or _62908_ (_11277_, _11276_, _11262_);
  and _62909_ (_11278_, _11277_, _11261_);
  nor _62910_ (_11279_, _11278_, _11258_);
  not _62911_ (_11280_, _11279_);
  and _62912_ (_11281_, _11280_, _11257_);
  or _62913_ (_11282_, _11281_, _11255_);
  and _62914_ (_11283_, _11282_, _11254_);
  nor _62915_ (_11284_, _11283_, _11251_);
  and _62916_ (_11285_, _11284_, _11039_);
  nor _62917_ (_11286_, _11284_, _11039_);
  or _62918_ (_11287_, _11286_, _11285_);
  or _62919_ (_11288_, _11287_, _11248_);
  and _62920_ (_11289_, _11288_, _11250_);
  and _62921_ (_11290_, _06471_, _06360_);
  or _62922_ (_11291_, _11290_, _11289_);
  not _62923_ (_11292_, _11290_);
  and _62924_ (_11293_, _09172_, \oc8051_golden_model_1.ACC [6]);
  or _62925_ (_11294_, _09172_, \oc8051_golden_model_1.ACC [6]);
  not _62926_ (_11295_, _11293_);
  and _62927_ (_11296_, _11295_, _11294_);
  and _62928_ (_11297_, _09218_, \oc8051_golden_model_1.ACC [5]);
  nor _62929_ (_11298_, _09218_, \oc8051_golden_model_1.ACC [5]);
  or _62930_ (_11299_, _11298_, _11297_);
  and _62931_ (_11300_, _09264_, \oc8051_golden_model_1.ACC [4]);
  not _62932_ (_11301_, _11300_);
  or _62933_ (_11302_, _09264_, \oc8051_golden_model_1.ACC [4]);
  and _62934_ (_11303_, _11301_, _11302_);
  and _62935_ (_11304_, _09310_, \oc8051_golden_model_1.ACC [3]);
  nor _62936_ (_11305_, _09310_, \oc8051_golden_model_1.ACC [3]);
  and _62937_ (_11306_, _09356_, \oc8051_golden_model_1.ACC [2]);
  nor _62938_ (_11307_, _09356_, \oc8051_golden_model_1.ACC [2]);
  nor _62939_ (_11308_, _11306_, _11307_);
  and _62940_ (_11309_, _09402_, \oc8051_golden_model_1.ACC [1]);
  nand _62941_ (_11310_, _09401_, _09379_);
  and _62942_ (_11311_, _11310_, _06097_);
  nor _62943_ (_11312_, _11309_, _11311_);
  and _62944_ (_11313_, _09447_, \oc8051_golden_model_1.ACC [0]);
  and _62945_ (_11314_, _11313_, _11312_);
  nor _62946_ (_11315_, _11314_, _11309_);
  not _62947_ (_11316_, _11315_);
  and _62948_ (_11317_, _11316_, _11308_);
  nor _62949_ (_11318_, _11317_, _11306_);
  nor _62950_ (_11319_, _11318_, _11305_);
  or _62951_ (_11320_, _11319_, _11304_);
  nand _62952_ (_11321_, _11320_, _11303_);
  and _62953_ (_11322_, _11321_, _11301_);
  nor _62954_ (_11323_, _11322_, _11299_);
  or _62955_ (_11324_, _11323_, _11297_);
  and _62956_ (_11325_, _11324_, _11296_);
  nor _62957_ (_11326_, _11325_, _11293_);
  and _62958_ (_11327_, _11326_, _11059_);
  nor _62959_ (_11328_, _11326_, _11059_);
  or _62960_ (_11329_, _11328_, _11327_);
  or _62961_ (_11330_, _11329_, _11292_);
  and _62962_ (_11331_, _11330_, _06364_);
  and _62963_ (_11332_, _11331_, _11291_);
  or _62964_ (_11333_, _11332_, _10602_);
  and _62965_ (_11334_, _11333_, _10567_);
  nor _62966_ (_11335_, _06397_, _10193_);
  not _62967_ (_11336_, _11335_);
  and _62968_ (_11337_, _06397_, _10193_);
  nor _62969_ (_11338_, _11335_, _11337_);
  nor _62970_ (_11339_, _06685_, _10237_);
  and _62971_ (_11340_, _06685_, _10237_);
  nor _62972_ (_11341_, _07093_, _10204_);
  not _62973_ (_11342_, _11341_);
  and _62974_ (_11343_, _07093_, _10204_);
  nor _62975_ (_11344_, _11341_, _11343_);
  nor _62976_ (_11345_, _06269_, _10334_);
  and _62977_ (_11346_, _06269_, _10334_);
  nor _62978_ (_11347_, _06727_, _10280_);
  and _62979_ (_11348_, _06727_, _10280_);
  nor _62980_ (_11349_, _11347_, _11348_);
  nor _62981_ (_11350_, _07127_, _06097_);
  nor _62982_ (_11351_, _06310_, _06071_);
  and _62983_ (_11352_, _07127_, \oc8051_golden_model_1.ACC [1]);
  nor _62984_ (_11353_, _07127_, \oc8051_golden_model_1.ACC [1]);
  nor _62985_ (_11354_, _11353_, _11352_);
  not _62986_ (_11355_, _11354_);
  and _62987_ (_11356_, _11355_, _11351_);
  nor _62988_ (_11357_, _11356_, _11350_);
  not _62989_ (_11358_, _11357_);
  and _62990_ (_11359_, _11358_, _11349_);
  nor _62991_ (_11360_, _11359_, _11347_);
  nor _62992_ (_11361_, _11360_, _11346_);
  or _62993_ (_11362_, _11361_, _11345_);
  nand _62994_ (_11363_, _11362_, _11344_);
  and _62995_ (_11364_, _11363_, _11342_);
  nor _62996_ (_11365_, _11364_, _11340_);
  or _62997_ (_11366_, _11365_, _11339_);
  nand _62998_ (_11367_, _11366_, _11338_);
  and _62999_ (_11368_, _11367_, _11336_);
  nor _63000_ (_11369_, _11368_, _11070_);
  and _63001_ (_11370_, _11368_, _11070_);
  or _63002_ (_11371_, _11370_, _11369_);
  and _63003_ (_11372_, _11371_, _10566_);
  or _63004_ (_11373_, _11372_, _10564_);
  or _63005_ (_11374_, _11373_, _11334_);
  and _63006_ (_11375_, _11374_, _10565_);
  or _63007_ (_11376_, _11375_, _06639_);
  and _63008_ (_11377_, _06489_, _05848_);
  not _63009_ (_11378_, _11377_);
  or _63010_ (_11379_, _10725_, _07048_);
  and _63011_ (_11380_, _11379_, _11378_);
  and _63012_ (_11381_, _11380_, _11376_);
  and _63013_ (_11382_, _06030_, _05848_);
  and _63014_ (_11383_, _10732_, _06071_);
  and _63015_ (_11384_, _11383_, _10334_);
  and _63016_ (_11385_, _11384_, _10204_);
  and _63017_ (_11386_, _11385_, _10237_);
  and _63018_ (_11387_, _11386_, _10193_);
  nor _63019_ (_11388_, _11387_, _08688_);
  and _63020_ (_11389_, _11387_, _08688_);
  or _63021_ (_11390_, _11389_, _11388_);
  and _63022_ (_11391_, _11390_, _11377_);
  or _63023_ (_11392_, _11391_, _11382_);
  or _63024_ (_11393_, _11392_, _11381_);
  nand _63025_ (_11394_, _11382_, _10967_);
  and _63026_ (_11395_, _11394_, _05990_);
  and _63027_ (_11396_, _11395_, _11393_);
  and _63028_ (_11397_, _10772_, _05989_);
  or _63029_ (_11398_, _11397_, _06646_);
  or _63030_ (_11399_, _11398_, _11396_);
  and _63031_ (_11400_, _06489_, _05996_);
  not _63032_ (_11401_, _11400_);
  and _63033_ (_11402_, _08605_, _08017_);
  or _63034_ (_11403_, _10603_, _06651_);
  or _63035_ (_11404_, _11403_, _11402_);
  and _63036_ (_11405_, _11404_, _11401_);
  and _63037_ (_11406_, _11405_, _11399_);
  and _63038_ (_11407_, _06030_, _05996_);
  and _63039_ (_11408_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and _63040_ (_11409_, _11408_, \oc8051_golden_model_1.ACC [2]);
  and _63041_ (_11410_, _11409_, \oc8051_golden_model_1.ACC [3]);
  and _63042_ (_11411_, _11410_, \oc8051_golden_model_1.ACC [4]);
  and _63043_ (_11412_, _11411_, \oc8051_golden_model_1.ACC [5]);
  and _63044_ (_11413_, _11412_, \oc8051_golden_model_1.ACC [6]);
  nor _63045_ (_11414_, _11413_, _08688_);
  and _63046_ (_11415_, _11413_, _08688_);
  or _63047_ (_11416_, _11415_, _11414_);
  and _63048_ (_11417_, _11416_, _11400_);
  or _63049_ (_11418_, _11417_, _11407_);
  or _63050_ (_11419_, _11418_, _11406_);
  nand _63051_ (_11420_, _11407_, _06071_);
  and _63052_ (_11421_, _11420_, _01442_);
  and _63053_ (_11422_, _11421_, _11419_);
  or _63054_ (_11423_, _11422_, _10563_);
  and _63055_ (_41497_, _11423_, _43634_);
  not _63056_ (_11424_, _08042_);
  and _63057_ (_11425_, _11424_, \oc8051_golden_model_1.PCON [7]);
  and _63058_ (_11426_, _09096_, _08042_);
  or _63059_ (_11427_, _11426_, _11425_);
  and _63060_ (_11428_, _11427_, _06615_);
  nor _63061_ (_11429_, _08107_, _11424_);
  or _63062_ (_11430_, _11429_, _11425_);
  or _63063_ (_11431_, _11430_, _06327_);
  and _63064_ (_11432_, _08791_, _08042_);
  or _63065_ (_11433_, _11432_, _11425_);
  or _63066_ (_11434_, _11433_, _07275_);
  and _63067_ (_11435_, _08042_, \oc8051_golden_model_1.ACC [7]);
  or _63068_ (_11436_, _11435_, _11425_);
  and _63069_ (_11437_, _11436_, _07259_);
  and _63070_ (_11438_, _07260_, \oc8051_golden_model_1.PCON [7]);
  or _63071_ (_11439_, _11438_, _06474_);
  or _63072_ (_11440_, _11439_, _11437_);
  and _63073_ (_11441_, _11440_, _06772_);
  and _63074_ (_11442_, _11441_, _11434_);
  and _63075_ (_11443_, _11430_, _06410_);
  or _63076_ (_11444_, _11443_, _11442_);
  and _63077_ (_11445_, _11444_, _06426_);
  and _63078_ (_11446_, _11436_, _06417_);
  or _63079_ (_11447_, _11446_, _10153_);
  or _63080_ (_11448_, _11447_, _11445_);
  and _63081_ (_11449_, _11448_, _11431_);
  or _63082_ (_11450_, _11449_, _09572_);
  and _63083_ (_11451_, _08778_, _08042_);
  or _63084_ (_11452_, _11425_, _06333_);
  or _63085_ (_11453_, _11452_, _11451_);
  and _63086_ (_11454_, _11453_, _06313_);
  and _63087_ (_11455_, _11454_, _11450_);
  and _63088_ (_11456_, _09076_, _08042_);
  or _63089_ (_11457_, _11456_, _11425_);
  and _63090_ (_11458_, _11457_, _06037_);
  or _63091_ (_11459_, _11458_, _06277_);
  or _63092_ (_11460_, _11459_, _11455_);
  and _63093_ (_11461_, _08880_, _08042_);
  or _63094_ (_11462_, _11461_, _11425_);
  or _63095_ (_11463_, _11462_, _06278_);
  and _63096_ (_11464_, _11463_, _11460_);
  or _63097_ (_11465_, _11464_, _06502_);
  and _63098_ (_11466_, _09090_, _08042_);
  or _63099_ (_11467_, _11425_, _07334_);
  or _63100_ (_11468_, _11467_, _11466_);
  and _63101_ (_11469_, _11468_, _07337_);
  and _63102_ (_11470_, _11469_, _11465_);
  or _63103_ (_11471_, _11470_, _11428_);
  and _63104_ (_11472_, _11471_, _07339_);
  or _63105_ (_11473_, _11425_, _08110_);
  and _63106_ (_11474_, _11462_, _06507_);
  and _63107_ (_11475_, _11474_, _11473_);
  or _63108_ (_11476_, _11475_, _11472_);
  and _63109_ (_11477_, _11476_, _07331_);
  and _63110_ (_11478_, _11436_, _06610_);
  and _63111_ (_11479_, _11478_, _11473_);
  or _63112_ (_11480_, _11479_, _06509_);
  or _63113_ (_11481_, _11480_, _11477_);
  and _63114_ (_11482_, _09087_, _08042_);
  or _63115_ (_11483_, _11425_, _09107_);
  or _63116_ (_11484_, _11483_, _11482_);
  and _63117_ (_11485_, _11484_, _09112_);
  and _63118_ (_11486_, _11485_, _11481_);
  nor _63119_ (_11487_, _09095_, _11424_);
  or _63120_ (_11488_, _11487_, _11425_);
  and _63121_ (_11489_, _11488_, _06602_);
  or _63122_ (_11490_, _11489_, _06639_);
  or _63123_ (_11491_, _11490_, _11486_);
  or _63124_ (_11492_, _11433_, _07048_);
  and _63125_ (_11493_, _11492_, _06651_);
  and _63126_ (_11494_, _11493_, _11491_);
  and _63127_ (_11495_, _08605_, _08042_);
  or _63128_ (_11496_, _11495_, _11425_);
  and _63129_ (_11497_, _11496_, _06646_);
  or _63130_ (_11498_, _11497_, _01446_);
  or _63131_ (_11499_, _11498_, _11494_);
  or _63132_ (_11500_, _01442_, \oc8051_golden_model_1.PCON [7]);
  and _63133_ (_11501_, _11500_, _43634_);
  and _63134_ (_41498_, _11501_, _11499_);
  not _63135_ (_11502_, _07965_);
  and _63136_ (_11503_, _11502_, \oc8051_golden_model_1.TMOD [7]);
  and _63137_ (_11504_, _09096_, _07965_);
  or _63138_ (_11505_, _11504_, _11503_);
  and _63139_ (_11506_, _11505_, _06615_);
  nor _63140_ (_11507_, _08107_, _11502_);
  or _63141_ (_11508_, _11507_, _11503_);
  or _63142_ (_11509_, _11508_, _06327_);
  and _63143_ (_11510_, _08791_, _07965_);
  or _63144_ (_11511_, _11510_, _11503_);
  or _63145_ (_11512_, _11511_, _07275_);
  and _63146_ (_11513_, _07965_, \oc8051_golden_model_1.ACC [7]);
  or _63147_ (_11514_, _11513_, _11503_);
  and _63148_ (_11515_, _11514_, _07259_);
  and _63149_ (_11516_, _07260_, \oc8051_golden_model_1.TMOD [7]);
  or _63150_ (_11517_, _11516_, _06474_);
  or _63151_ (_11518_, _11517_, _11515_);
  and _63152_ (_11519_, _11518_, _06772_);
  and _63153_ (_11520_, _11519_, _11512_);
  and _63154_ (_11521_, _11508_, _06410_);
  or _63155_ (_11522_, _11521_, _11520_);
  and _63156_ (_11523_, _11522_, _06426_);
  and _63157_ (_11524_, _11514_, _06417_);
  or _63158_ (_11525_, _11524_, _10153_);
  or _63159_ (_11526_, _11525_, _11523_);
  and _63160_ (_11527_, _11526_, _11509_);
  or _63161_ (_11528_, _11527_, _09572_);
  and _63162_ (_11529_, _08778_, _07965_);
  or _63163_ (_11530_, _11503_, _06333_);
  or _63164_ (_11531_, _11530_, _11529_);
  and _63165_ (_11532_, _11531_, _06313_);
  and _63166_ (_11533_, _11532_, _11528_);
  and _63167_ (_11534_, _09076_, _07965_);
  or _63168_ (_11535_, _11534_, _11503_);
  and _63169_ (_11536_, _11535_, _06037_);
  or _63170_ (_11537_, _11536_, _06277_);
  or _63171_ (_11538_, _11537_, _11533_);
  and _63172_ (_11539_, _08880_, _07965_);
  or _63173_ (_11540_, _11539_, _11503_);
  or _63174_ (_11541_, _11540_, _06278_);
  and _63175_ (_11542_, _11541_, _11538_);
  or _63176_ (_11543_, _11542_, _06502_);
  and _63177_ (_11544_, _09090_, _07965_);
  or _63178_ (_11545_, _11503_, _07334_);
  or _63179_ (_11546_, _11545_, _11544_);
  and _63180_ (_11547_, _11546_, _07337_);
  and _63181_ (_11548_, _11547_, _11543_);
  or _63182_ (_11549_, _11548_, _11506_);
  and _63183_ (_11550_, _11549_, _07339_);
  or _63184_ (_11551_, _11503_, _08110_);
  and _63185_ (_11552_, _11540_, _06507_);
  and _63186_ (_11553_, _11552_, _11551_);
  or _63187_ (_11554_, _11553_, _11550_);
  and _63188_ (_11555_, _11554_, _07331_);
  and _63189_ (_11556_, _11514_, _06610_);
  and _63190_ (_11557_, _11556_, _11551_);
  or _63191_ (_11558_, _11557_, _06509_);
  or _63192_ (_11559_, _11558_, _11555_);
  and _63193_ (_11560_, _09087_, _07965_);
  or _63194_ (_11561_, _11503_, _09107_);
  or _63195_ (_11562_, _11561_, _11560_);
  and _63196_ (_11563_, _11562_, _09112_);
  and _63197_ (_11564_, _11563_, _11559_);
  nor _63198_ (_11565_, _09095_, _11502_);
  or _63199_ (_11566_, _11565_, _11503_);
  and _63200_ (_11567_, _11566_, _06602_);
  or _63201_ (_11568_, _11567_, _06639_);
  or _63202_ (_11569_, _11568_, _11564_);
  or _63203_ (_11570_, _11511_, _07048_);
  and _63204_ (_11571_, _11570_, _06651_);
  and _63205_ (_11572_, _11571_, _11569_);
  and _63206_ (_11573_, _08605_, _07965_);
  or _63207_ (_11574_, _11573_, _11503_);
  and _63208_ (_11575_, _11574_, _06646_);
  or _63209_ (_11576_, _11575_, _01446_);
  or _63210_ (_11577_, _11576_, _11572_);
  or _63211_ (_11578_, _01442_, \oc8051_golden_model_1.TMOD [7]);
  and _63212_ (_11579_, _11578_, _43634_);
  and _63213_ (_41499_, _11579_, _11577_);
  not _63214_ (_11580_, \oc8051_golden_model_1.DPL [7]);
  nor _63215_ (_11581_, _08001_, _11580_);
  and _63216_ (_11582_, _09096_, _08001_);
  or _63217_ (_11583_, _11582_, _11581_);
  and _63218_ (_11584_, _11583_, _06615_);
  not _63219_ (_11585_, _08001_);
  nor _63220_ (_11586_, _08107_, _11585_);
  or _63221_ (_11587_, _11586_, _11581_);
  or _63222_ (_11588_, _11587_, _06327_);
  and _63223_ (_11589_, _08791_, _08001_);
  or _63224_ (_11590_, _11589_, _11581_);
  or _63225_ (_11591_, _11590_, _07275_);
  and _63226_ (_11592_, _08158_, \oc8051_golden_model_1.ACC [7]);
  or _63227_ (_11593_, _11592_, _11581_);
  and _63228_ (_11594_, _11593_, _07259_);
  nor _63229_ (_11595_, _07259_, _11580_);
  or _63230_ (_11596_, _11595_, _06474_);
  or _63231_ (_11597_, _11596_, _11594_);
  and _63232_ (_11598_, _11597_, _06772_);
  and _63233_ (_11599_, _11598_, _11591_);
  and _63234_ (_11600_, _11587_, _06410_);
  or _63235_ (_11601_, _11600_, _06417_);
  or _63236_ (_11602_, _11601_, _11599_);
  and _63237_ (_11603_, _06443_, _06030_);
  not _63238_ (_11604_, _11603_);
  or _63239_ (_11605_, _11593_, _06426_);
  and _63240_ (_11606_, _11605_, _11604_);
  and _63241_ (_11607_, _11606_, _11602_);
  and _63242_ (_11608_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _63243_ (_11609_, _11608_, \oc8051_golden_model_1.DPL [2]);
  and _63244_ (_11610_, _11609_, \oc8051_golden_model_1.DPL [3]);
  and _63245_ (_11611_, _11610_, \oc8051_golden_model_1.DPL [4]);
  and _63246_ (_11612_, _11611_, \oc8051_golden_model_1.DPL [5]);
  and _63247_ (_11613_, _11612_, \oc8051_golden_model_1.DPL [6]);
  nor _63248_ (_11614_, _11613_, \oc8051_golden_model_1.DPL [7]);
  and _63249_ (_11615_, _11613_, \oc8051_golden_model_1.DPL [7]);
  nor _63250_ (_11616_, _11615_, _11614_);
  and _63251_ (_11617_, _11616_, _11603_);
  or _63252_ (_11618_, _11617_, _11607_);
  and _63253_ (_11619_, _11618_, _06487_);
  nor _63254_ (_11620_, _08879_, _06487_);
  or _63255_ (_11621_, _11620_, _10153_);
  or _63256_ (_11622_, _11621_, _11619_);
  and _63257_ (_11623_, _11622_, _11588_);
  or _63258_ (_11624_, _11623_, _09572_);
  and _63259_ (_11625_, _08778_, _08158_);
  or _63260_ (_11626_, _11581_, _06333_);
  or _63261_ (_11627_, _11626_, _11625_);
  and _63262_ (_11628_, _11627_, _06313_);
  and _63263_ (_11629_, _11628_, _11624_);
  and _63264_ (_11630_, _09076_, _08158_);
  or _63265_ (_11631_, _11630_, _11581_);
  and _63266_ (_11632_, _11631_, _06037_);
  or _63267_ (_11633_, _11632_, _06277_);
  or _63268_ (_11634_, _11633_, _11629_);
  and _63269_ (_11635_, _08880_, _08158_);
  or _63270_ (_11636_, _11635_, _11581_);
  or _63271_ (_11637_, _11636_, _06278_);
  and _63272_ (_11638_, _11637_, _11634_);
  or _63273_ (_11639_, _11638_, _06502_);
  and _63274_ (_11640_, _09090_, _08001_);
  or _63275_ (_11641_, _11581_, _07334_);
  or _63276_ (_11642_, _11641_, _11640_);
  and _63277_ (_11643_, _11642_, _07337_);
  and _63278_ (_11644_, _11643_, _11639_);
  or _63279_ (_11645_, _11644_, _11584_);
  and _63280_ (_11646_, _11645_, _07339_);
  or _63281_ (_11647_, _11581_, _08110_);
  and _63282_ (_11648_, _11636_, _06507_);
  and _63283_ (_11649_, _11648_, _11647_);
  or _63284_ (_11650_, _11649_, _11646_);
  and _63285_ (_11651_, _11650_, _07331_);
  and _63286_ (_11652_, _11593_, _06610_);
  and _63287_ (_11653_, _11652_, _11647_);
  or _63288_ (_11654_, _11653_, _06509_);
  or _63289_ (_11655_, _11654_, _11651_);
  and _63290_ (_11656_, _09087_, _08001_);
  or _63291_ (_11657_, _11581_, _09107_);
  or _63292_ (_11658_, _11657_, _11656_);
  and _63293_ (_11659_, _11658_, _09112_);
  and _63294_ (_11660_, _11659_, _11655_);
  nor _63295_ (_11661_, _09095_, _11585_);
  or _63296_ (_11662_, _11661_, _11581_);
  and _63297_ (_11663_, _11662_, _06602_);
  or _63298_ (_11664_, _11663_, _06639_);
  or _63299_ (_11665_, _11664_, _11660_);
  or _63300_ (_11666_, _11590_, _07048_);
  and _63301_ (_11667_, _11666_, _06651_);
  and _63302_ (_11668_, _11667_, _11665_);
  and _63303_ (_11669_, _08605_, _08001_);
  or _63304_ (_11670_, _11669_, _11581_);
  and _63305_ (_11671_, _11670_, _06646_);
  or _63306_ (_11672_, _11671_, _01446_);
  or _63307_ (_11673_, _11672_, _11668_);
  or _63308_ (_11674_, _01442_, \oc8051_golden_model_1.DPL [7]);
  and _63309_ (_11675_, _11674_, _43634_);
  and _63310_ (_41501_, _11675_, _11673_);
  not _63311_ (_11676_, \oc8051_golden_model_1.DPH [7]);
  nor _63312_ (_11677_, _08153_, _11676_);
  and _63313_ (_11678_, _09096_, _07995_);
  or _63314_ (_11679_, _11678_, _11677_);
  and _63315_ (_11680_, _11679_, _06615_);
  not _63316_ (_11681_, _07995_);
  nor _63317_ (_11682_, _08107_, _11681_);
  or _63318_ (_11683_, _11682_, _11677_);
  or _63319_ (_11684_, _11683_, _06327_);
  and _63320_ (_11685_, _08791_, _07995_);
  or _63321_ (_11686_, _11685_, _11677_);
  or _63322_ (_11687_, _11686_, _07275_);
  and _63323_ (_11688_, _08153_, \oc8051_golden_model_1.ACC [7]);
  or _63324_ (_11689_, _11688_, _11677_);
  and _63325_ (_11690_, _11689_, _07259_);
  nor _63326_ (_11691_, _07259_, _11676_);
  or _63327_ (_11692_, _11691_, _06474_);
  or _63328_ (_11693_, _11692_, _11690_);
  and _63329_ (_11694_, _11693_, _06772_);
  and _63330_ (_11695_, _11694_, _11687_);
  and _63331_ (_11696_, _11683_, _06410_);
  or _63332_ (_11697_, _11696_, _06417_);
  or _63333_ (_11698_, _11697_, _11695_);
  or _63334_ (_11699_, _11689_, _06426_);
  and _63335_ (_11700_, _11699_, _11604_);
  and _63336_ (_11701_, _11700_, _11698_);
  and _63337_ (_11702_, _11615_, \oc8051_golden_model_1.DPH [0]);
  and _63338_ (_11703_, _11702_, \oc8051_golden_model_1.DPH [1]);
  and _63339_ (_11704_, _11703_, \oc8051_golden_model_1.DPH [2]);
  and _63340_ (_11705_, _11704_, \oc8051_golden_model_1.DPH [3]);
  and _63341_ (_11706_, _11705_, \oc8051_golden_model_1.DPH [4]);
  and _63342_ (_11707_, _11706_, \oc8051_golden_model_1.DPH [5]);
  and _63343_ (_11708_, _11707_, \oc8051_golden_model_1.DPH [6]);
  nand _63344_ (_11709_, _11708_, \oc8051_golden_model_1.DPH [7]);
  or _63345_ (_11710_, _11708_, \oc8051_golden_model_1.DPH [7]);
  and _63346_ (_11711_, _11710_, _11709_);
  and _63347_ (_11712_, _11711_, _11603_);
  or _63348_ (_11713_, _11712_, _11701_);
  and _63349_ (_11714_, _11713_, _06487_);
  and _63350_ (_11715_, _06486_, _06238_);
  or _63351_ (_11716_, _11715_, _10153_);
  or _63352_ (_11717_, _11716_, _11714_);
  and _63353_ (_11718_, _11717_, _11684_);
  or _63354_ (_11719_, _11718_, _09572_);
  and _63355_ (_11720_, _08778_, _08153_);
  or _63356_ (_11721_, _11677_, _06333_);
  or _63357_ (_11722_, _11721_, _11720_);
  and _63358_ (_11723_, _11722_, _06313_);
  and _63359_ (_11724_, _11723_, _11719_);
  and _63360_ (_11725_, _09076_, _08153_);
  or _63361_ (_11726_, _11725_, _11677_);
  and _63362_ (_11727_, _11726_, _06037_);
  or _63363_ (_11728_, _11727_, _06277_);
  or _63364_ (_11729_, _11728_, _11724_);
  and _63365_ (_11730_, _08880_, _08153_);
  or _63366_ (_11731_, _11730_, _11677_);
  or _63367_ (_11732_, _11731_, _06278_);
  and _63368_ (_11733_, _11732_, _11729_);
  or _63369_ (_11734_, _11733_, _06502_);
  and _63370_ (_11735_, _09090_, _07995_);
  or _63371_ (_11736_, _11677_, _07334_);
  or _63372_ (_11737_, _11736_, _11735_);
  and _63373_ (_11738_, _11737_, _07337_);
  and _63374_ (_11739_, _11738_, _11734_);
  or _63375_ (_11740_, _11739_, _11680_);
  and _63376_ (_11741_, _11740_, _07339_);
  or _63377_ (_11742_, _11677_, _08110_);
  and _63378_ (_11743_, _11731_, _06507_);
  and _63379_ (_11744_, _11743_, _11742_);
  or _63380_ (_11745_, _11744_, _11741_);
  and _63381_ (_11746_, _11745_, _07331_);
  and _63382_ (_11747_, _11689_, _06610_);
  and _63383_ (_11748_, _11747_, _11742_);
  or _63384_ (_11749_, _11748_, _06509_);
  or _63385_ (_11750_, _11749_, _11746_);
  and _63386_ (_11751_, _09087_, _07995_);
  or _63387_ (_11752_, _11677_, _09107_);
  or _63388_ (_11753_, _11752_, _11751_);
  and _63389_ (_11754_, _11753_, _09112_);
  and _63390_ (_11755_, _11754_, _11750_);
  nor _63391_ (_11756_, _09095_, _11681_);
  or _63392_ (_11757_, _11756_, _11677_);
  and _63393_ (_11758_, _11757_, _06602_);
  or _63394_ (_11759_, _11758_, _06639_);
  or _63395_ (_11760_, _11759_, _11755_);
  or _63396_ (_11761_, _11686_, _07048_);
  and _63397_ (_11762_, _11761_, _06651_);
  and _63398_ (_11763_, _11762_, _11760_);
  and _63399_ (_11764_, _08605_, _07995_);
  or _63400_ (_11765_, _11764_, _11677_);
  and _63401_ (_11766_, _11765_, _06646_);
  or _63402_ (_11767_, _11766_, _01446_);
  or _63403_ (_11768_, _11767_, _11763_);
  or _63404_ (_11769_, _01442_, \oc8051_golden_model_1.DPH [7]);
  and _63405_ (_11770_, _11769_, _43634_);
  and _63406_ (_41502_, _11770_, _11768_);
  not _63407_ (_11771_, _07991_);
  and _63408_ (_11772_, _11771_, \oc8051_golden_model_1.TL1 [7]);
  and _63409_ (_11773_, _09096_, _07991_);
  or _63410_ (_11774_, _11773_, _11772_);
  and _63411_ (_11775_, _11774_, _06615_);
  nor _63412_ (_11776_, _08107_, _11771_);
  or _63413_ (_11777_, _11776_, _11772_);
  or _63414_ (_11778_, _11777_, _06327_);
  and _63415_ (_11779_, _08791_, _07991_);
  or _63416_ (_11780_, _11779_, _11772_);
  or _63417_ (_11781_, _11780_, _07275_);
  and _63418_ (_11782_, _07991_, \oc8051_golden_model_1.ACC [7]);
  or _63419_ (_11783_, _11782_, _11772_);
  and _63420_ (_11784_, _11783_, _07259_);
  and _63421_ (_11785_, _07260_, \oc8051_golden_model_1.TL1 [7]);
  or _63422_ (_11786_, _11785_, _06474_);
  or _63423_ (_11787_, _11786_, _11784_);
  and _63424_ (_11788_, _11787_, _06772_);
  and _63425_ (_11789_, _11788_, _11781_);
  and _63426_ (_11790_, _11777_, _06410_);
  or _63427_ (_11791_, _11790_, _11789_);
  and _63428_ (_11792_, _11791_, _06426_);
  and _63429_ (_11793_, _11783_, _06417_);
  or _63430_ (_11794_, _11793_, _10153_);
  or _63431_ (_11795_, _11794_, _11792_);
  and _63432_ (_11796_, _11795_, _11778_);
  or _63433_ (_11797_, _11796_, _09572_);
  and _63434_ (_11798_, _08778_, _07991_);
  or _63435_ (_11799_, _11772_, _06333_);
  or _63436_ (_11800_, _11799_, _11798_);
  and _63437_ (_11801_, _11800_, _06313_);
  and _63438_ (_11802_, _11801_, _11797_);
  and _63439_ (_11803_, _09076_, _07991_);
  or _63440_ (_11804_, _11803_, _11772_);
  and _63441_ (_11805_, _11804_, _06037_);
  or _63442_ (_11806_, _11805_, _06277_);
  or _63443_ (_11807_, _11806_, _11802_);
  and _63444_ (_11808_, _08880_, _07991_);
  or _63445_ (_11809_, _11808_, _11772_);
  or _63446_ (_11810_, _11809_, _06278_);
  and _63447_ (_11811_, _11810_, _11807_);
  or _63448_ (_11812_, _11811_, _06502_);
  and _63449_ (_11813_, _09090_, _07991_);
  or _63450_ (_11814_, _11772_, _07334_);
  or _63451_ (_11815_, _11814_, _11813_);
  and _63452_ (_11816_, _11815_, _07337_);
  and _63453_ (_11817_, _11816_, _11812_);
  or _63454_ (_11818_, _11817_, _11775_);
  and _63455_ (_11819_, _11818_, _07339_);
  or _63456_ (_11820_, _11772_, _08110_);
  and _63457_ (_11821_, _11809_, _06507_);
  and _63458_ (_11822_, _11821_, _11820_);
  or _63459_ (_11823_, _11822_, _11819_);
  and _63460_ (_11824_, _11823_, _07331_);
  and _63461_ (_11825_, _11783_, _06610_);
  and _63462_ (_11826_, _11825_, _11820_);
  or _63463_ (_11827_, _11826_, _06509_);
  or _63464_ (_11828_, _11827_, _11824_);
  and _63465_ (_11829_, _09087_, _07991_);
  or _63466_ (_11830_, _11772_, _09107_);
  or _63467_ (_11831_, _11830_, _11829_);
  and _63468_ (_11832_, _11831_, _09112_);
  and _63469_ (_11833_, _11832_, _11828_);
  nor _63470_ (_11834_, _09095_, _11771_);
  or _63471_ (_11835_, _11834_, _11772_);
  and _63472_ (_11836_, _11835_, _06602_);
  or _63473_ (_11837_, _11836_, _06639_);
  or _63474_ (_11838_, _11837_, _11833_);
  or _63475_ (_11839_, _11780_, _07048_);
  and _63476_ (_11840_, _11839_, _06651_);
  and _63477_ (_11841_, _11840_, _11838_);
  and _63478_ (_11842_, _08605_, _07991_);
  or _63479_ (_11843_, _11842_, _11772_);
  and _63480_ (_11844_, _11843_, _06646_);
  or _63481_ (_11845_, _11844_, _01446_);
  or _63482_ (_11846_, _11845_, _11841_);
  or _63483_ (_11847_, _01442_, \oc8051_golden_model_1.TL1 [7]);
  and _63484_ (_11848_, _11847_, _43634_);
  and _63485_ (_41503_, _11848_, _11846_);
  not _63486_ (_11849_, _08133_);
  and _63487_ (_11850_, _11849_, \oc8051_golden_model_1.TL0 [7]);
  and _63488_ (_11851_, _09096_, _07976_);
  or _63489_ (_11852_, _11851_, _11850_);
  and _63490_ (_11853_, _11852_, _06615_);
  not _63491_ (_11854_, _07976_);
  nor _63492_ (_11855_, _08107_, _11854_);
  or _63493_ (_11856_, _11855_, _11850_);
  or _63494_ (_11857_, _11856_, _06327_);
  and _63495_ (_11858_, _08791_, _07976_);
  or _63496_ (_11859_, _11858_, _11850_);
  or _63497_ (_11860_, _11859_, _07275_);
  and _63498_ (_11861_, _08133_, \oc8051_golden_model_1.ACC [7]);
  or _63499_ (_11862_, _11861_, _11850_);
  and _63500_ (_11863_, _11862_, _07259_);
  and _63501_ (_11864_, _07260_, \oc8051_golden_model_1.TL0 [7]);
  or _63502_ (_11865_, _11864_, _06474_);
  or _63503_ (_11866_, _11865_, _11863_);
  and _63504_ (_11867_, _11866_, _06772_);
  and _63505_ (_11868_, _11867_, _11860_);
  and _63506_ (_11869_, _11856_, _06410_);
  or _63507_ (_11870_, _11869_, _11868_);
  and _63508_ (_11871_, _11870_, _06426_);
  and _63509_ (_11872_, _11862_, _06417_);
  or _63510_ (_11873_, _11872_, _10153_);
  or _63511_ (_11874_, _11873_, _11871_);
  and _63512_ (_11875_, _11874_, _11857_);
  or _63513_ (_11876_, _11875_, _09572_);
  and _63514_ (_11877_, _08778_, _08133_);
  or _63515_ (_11878_, _11850_, _06333_);
  or _63516_ (_11879_, _11878_, _11877_);
  and _63517_ (_11880_, _11879_, _06313_);
  and _63518_ (_11881_, _11880_, _11876_);
  and _63519_ (_11882_, _09076_, _08133_);
  or _63520_ (_11883_, _11882_, _11850_);
  and _63521_ (_11884_, _11883_, _06037_);
  or _63522_ (_11885_, _11884_, _06277_);
  or _63523_ (_11886_, _11885_, _11881_);
  and _63524_ (_11887_, _08880_, _08133_);
  or _63525_ (_11888_, _11887_, _11850_);
  or _63526_ (_11889_, _11888_, _06278_);
  and _63527_ (_11890_, _11889_, _11886_);
  or _63528_ (_11891_, _11890_, _06502_);
  and _63529_ (_11892_, _09090_, _07976_);
  or _63530_ (_11893_, _11850_, _07334_);
  or _63531_ (_11894_, _11893_, _11892_);
  and _63532_ (_11895_, _11894_, _07337_);
  and _63533_ (_11896_, _11895_, _11891_);
  or _63534_ (_11897_, _11896_, _11853_);
  and _63535_ (_11898_, _11897_, _07339_);
  or _63536_ (_11899_, _11850_, _08110_);
  and _63537_ (_11900_, _11888_, _06507_);
  and _63538_ (_11901_, _11900_, _11899_);
  or _63539_ (_11902_, _11901_, _11898_);
  and _63540_ (_11903_, _11902_, _07331_);
  and _63541_ (_11904_, _11862_, _06610_);
  and _63542_ (_11905_, _11904_, _11899_);
  or _63543_ (_11906_, _11905_, _06509_);
  or _63544_ (_11907_, _11906_, _11903_);
  and _63545_ (_11908_, _09087_, _07976_);
  or _63546_ (_11909_, _11850_, _09107_);
  or _63547_ (_11910_, _11909_, _11908_);
  and _63548_ (_11911_, _11910_, _09112_);
  and _63549_ (_11912_, _11911_, _11907_);
  nor _63550_ (_11913_, _09095_, _11854_);
  or _63551_ (_11914_, _11913_, _11850_);
  and _63552_ (_11915_, _11914_, _06602_);
  or _63553_ (_11916_, _11915_, _06639_);
  or _63554_ (_11917_, _11916_, _11912_);
  or _63555_ (_11918_, _11859_, _07048_);
  and _63556_ (_11919_, _11918_, _06651_);
  and _63557_ (_11920_, _11919_, _11917_);
  and _63558_ (_11921_, _08605_, _07976_);
  or _63559_ (_11922_, _11921_, _11850_);
  and _63560_ (_11923_, _11922_, _06646_);
  or _63561_ (_11924_, _11923_, _01446_);
  or _63562_ (_11925_, _11924_, _11920_);
  or _63563_ (_11926_, _01442_, \oc8051_golden_model_1.TL0 [7]);
  and _63564_ (_11927_, _11926_, _43634_);
  and _63565_ (_41504_, _11927_, _11925_);
  and _63566_ (_11928_, _01446_, \oc8051_golden_model_1.TCON [7]);
  not _63567_ (_11929_, _08006_);
  and _63568_ (_11930_, _11929_, \oc8051_golden_model_1.TCON [7]);
  and _63569_ (_11931_, _09096_, _08006_);
  or _63570_ (_11932_, _11931_, _11930_);
  and _63571_ (_11933_, _11932_, _06615_);
  nor _63572_ (_11934_, _08107_, _11929_);
  or _63573_ (_11935_, _11934_, _11930_);
  or _63574_ (_11936_, _11935_, _06327_);
  not _63575_ (_11937_, _08633_);
  and _63576_ (_11938_, _11937_, \oc8051_golden_model_1.TCON [7]);
  and _63577_ (_11939_, _08668_, _08633_);
  or _63578_ (_11940_, _11939_, _11938_);
  and _63579_ (_11941_, _11940_, _06352_);
  and _63580_ (_11942_, _08791_, _08006_);
  or _63581_ (_11943_, _11942_, _11930_);
  or _63582_ (_11944_, _11943_, _07275_);
  and _63583_ (_11945_, _08006_, \oc8051_golden_model_1.ACC [7]);
  or _63584_ (_11946_, _11945_, _11930_);
  and _63585_ (_11947_, _11946_, _07259_);
  and _63586_ (_11948_, _07260_, \oc8051_golden_model_1.TCON [7]);
  or _63587_ (_11949_, _11948_, _06474_);
  or _63588_ (_11950_, _11949_, _11947_);
  and _63589_ (_11951_, _11950_, _06357_);
  and _63590_ (_11952_, _11951_, _11944_);
  and _63591_ (_11953_, _08672_, _08633_);
  or _63592_ (_11954_, _11953_, _11938_);
  and _63593_ (_11955_, _11954_, _06356_);
  or _63594_ (_11956_, _11955_, _06410_);
  or _63595_ (_11957_, _11956_, _11952_);
  or _63596_ (_11958_, _11935_, _06772_);
  and _63597_ (_11959_, _11958_, _11957_);
  or _63598_ (_11960_, _11959_, _06417_);
  or _63599_ (_11961_, _11946_, _06426_);
  and _63600_ (_11962_, _11961_, _06353_);
  and _63601_ (_11963_, _11962_, _11960_);
  or _63602_ (_11964_, _11963_, _11941_);
  and _63603_ (_11965_, _11964_, _06346_);
  and _63604_ (_11966_, _08810_, _08633_);
  or _63605_ (_11967_, _11966_, _11938_);
  and _63606_ (_11968_, _11967_, _06345_);
  or _63607_ (_11969_, _11968_, _11965_);
  and _63608_ (_11970_, _11969_, _06340_);
  and _63609_ (_11971_, _08828_, _08633_);
  or _63610_ (_11972_, _11971_, _11938_);
  and _63611_ (_11973_, _11972_, _06339_);
  or _63612_ (_11974_, _11973_, _10153_);
  or _63613_ (_11975_, _11974_, _11970_);
  and _63614_ (_11976_, _11975_, _11936_);
  or _63615_ (_11977_, _11976_, _09572_);
  and _63616_ (_11978_, _08778_, _08006_);
  or _63617_ (_11979_, _11930_, _06333_);
  or _63618_ (_11980_, _11979_, _11978_);
  and _63619_ (_11981_, _11980_, _06313_);
  and _63620_ (_11982_, _11981_, _11977_);
  and _63621_ (_11983_, _09076_, _08006_);
  or _63622_ (_11984_, _11983_, _11930_);
  and _63623_ (_11985_, _11984_, _06037_);
  or _63624_ (_11986_, _11985_, _06277_);
  or _63625_ (_11987_, _11986_, _11982_);
  and _63626_ (_11988_, _08880_, _08006_);
  or _63627_ (_11989_, _11988_, _11930_);
  or _63628_ (_11990_, _11989_, _06278_);
  and _63629_ (_11991_, _11990_, _11987_);
  or _63630_ (_11992_, _11991_, _06502_);
  and _63631_ (_11993_, _09090_, _08006_);
  or _63632_ (_11994_, _11930_, _07334_);
  or _63633_ (_11995_, _11994_, _11993_);
  and _63634_ (_11996_, _11995_, _07337_);
  and _63635_ (_11997_, _11996_, _11992_);
  or _63636_ (_11998_, _11997_, _11933_);
  and _63637_ (_11999_, _11998_, _07339_);
  or _63638_ (_12000_, _11930_, _08110_);
  and _63639_ (_12001_, _11989_, _06507_);
  and _63640_ (_12002_, _12001_, _12000_);
  or _63641_ (_12003_, _12002_, _11999_);
  and _63642_ (_12004_, _12003_, _07331_);
  and _63643_ (_12005_, _11946_, _06610_);
  and _63644_ (_12006_, _12005_, _12000_);
  or _63645_ (_12007_, _12006_, _06509_);
  or _63646_ (_12008_, _12007_, _12004_);
  and _63647_ (_12009_, _09087_, _08006_);
  or _63648_ (_12010_, _11930_, _09107_);
  or _63649_ (_12011_, _12010_, _12009_);
  and _63650_ (_12012_, _12011_, _09112_);
  and _63651_ (_12013_, _12012_, _12008_);
  nor _63652_ (_12014_, _09095_, _11929_);
  or _63653_ (_12015_, _12014_, _11930_);
  and _63654_ (_12016_, _12015_, _06602_);
  or _63655_ (_12017_, _12016_, _06639_);
  or _63656_ (_12018_, _12017_, _12013_);
  or _63657_ (_12019_, _11943_, _07048_);
  and _63658_ (_12020_, _12019_, _05990_);
  and _63659_ (_12021_, _12020_, _12018_);
  and _63660_ (_12022_, _11940_, _05989_);
  or _63661_ (_12023_, _12022_, _06646_);
  or _63662_ (_12024_, _12023_, _12021_);
  and _63663_ (_12025_, _08605_, _08006_);
  or _63664_ (_12026_, _11930_, _06651_);
  or _63665_ (_12027_, _12026_, _12025_);
  and _63666_ (_12028_, _12027_, _01442_);
  and _63667_ (_12029_, _12028_, _12024_);
  or _63668_ (_12030_, _12029_, _11928_);
  and _63669_ (_41505_, _12030_, _43634_);
  not _63670_ (_12031_, _07981_);
  and _63671_ (_12032_, _12031_, \oc8051_golden_model_1.TH1 [7]);
  and _63672_ (_12033_, _09096_, _07981_);
  or _63673_ (_12034_, _12033_, _12032_);
  and _63674_ (_12035_, _12034_, _06615_);
  and _63675_ (_12036_, _08791_, _07981_);
  or _63676_ (_12037_, _12036_, _12032_);
  or _63677_ (_12038_, _12037_, _07275_);
  and _63678_ (_12039_, _07981_, \oc8051_golden_model_1.ACC [7]);
  or _63679_ (_12040_, _12039_, _12032_);
  and _63680_ (_12041_, _12040_, _07259_);
  and _63681_ (_12042_, _07260_, \oc8051_golden_model_1.TH1 [7]);
  or _63682_ (_12043_, _12042_, _06474_);
  or _63683_ (_12044_, _12043_, _12041_);
  and _63684_ (_12045_, _12044_, _06772_);
  and _63685_ (_12046_, _12045_, _12038_);
  nor _63686_ (_12047_, _08107_, _12031_);
  or _63687_ (_12048_, _12047_, _12032_);
  and _63688_ (_12049_, _12048_, _06410_);
  or _63689_ (_12050_, _12049_, _12046_);
  and _63690_ (_12051_, _12050_, _06426_);
  and _63691_ (_12052_, _12040_, _06417_);
  or _63692_ (_12053_, _12052_, _10153_);
  or _63693_ (_12054_, _12053_, _12051_);
  or _63694_ (_12055_, _12048_, _06327_);
  and _63695_ (_12056_, _12055_, _12054_);
  or _63696_ (_12057_, _12056_, _09572_);
  and _63697_ (_12058_, _08778_, _07981_);
  or _63698_ (_12059_, _12032_, _06333_);
  or _63699_ (_12060_, _12059_, _12058_);
  and _63700_ (_12061_, _12060_, _06313_);
  and _63701_ (_12062_, _12061_, _12057_);
  and _63702_ (_12063_, _09076_, _07981_);
  or _63703_ (_12064_, _12063_, _12032_);
  and _63704_ (_12065_, _12064_, _06037_);
  or _63705_ (_12066_, _12065_, _06277_);
  or _63706_ (_12067_, _12066_, _12062_);
  and _63707_ (_12068_, _08880_, _07981_);
  or _63708_ (_12069_, _12068_, _12032_);
  or _63709_ (_12070_, _12069_, _06278_);
  and _63710_ (_12071_, _12070_, _12067_);
  or _63711_ (_12072_, _12071_, _06502_);
  and _63712_ (_12073_, _09090_, _07981_);
  or _63713_ (_12074_, _12032_, _07334_);
  or _63714_ (_12075_, _12074_, _12073_);
  and _63715_ (_12076_, _12075_, _07337_);
  and _63716_ (_12077_, _12076_, _12072_);
  or _63717_ (_12078_, _12077_, _12035_);
  and _63718_ (_12079_, _12078_, _07339_);
  or _63719_ (_12080_, _12032_, _08110_);
  and _63720_ (_12081_, _12069_, _06507_);
  and _63721_ (_12082_, _12081_, _12080_);
  or _63722_ (_12083_, _12082_, _12079_);
  and _63723_ (_12084_, _12083_, _07331_);
  and _63724_ (_12085_, _12040_, _06610_);
  and _63725_ (_12086_, _12085_, _12080_);
  or _63726_ (_12087_, _12086_, _06509_);
  or _63727_ (_12088_, _12087_, _12084_);
  and _63728_ (_12089_, _09087_, _07981_);
  or _63729_ (_12090_, _12032_, _09107_);
  or _63730_ (_12091_, _12090_, _12089_);
  and _63731_ (_12092_, _12091_, _09112_);
  and _63732_ (_12093_, _12092_, _12088_);
  nor _63733_ (_12094_, _09095_, _12031_);
  or _63734_ (_12095_, _12094_, _12032_);
  and _63735_ (_12096_, _12095_, _06602_);
  or _63736_ (_12097_, _12096_, _06639_);
  or _63737_ (_12098_, _12097_, _12093_);
  or _63738_ (_12099_, _12037_, _07048_);
  and _63739_ (_12100_, _12099_, _06651_);
  and _63740_ (_12101_, _12100_, _12098_);
  and _63741_ (_12102_, _08605_, _07981_);
  or _63742_ (_12103_, _12102_, _12032_);
  and _63743_ (_12104_, _12103_, _06646_);
  or _63744_ (_12105_, _12104_, _01446_);
  or _63745_ (_12106_, _12105_, _12101_);
  or _63746_ (_12107_, _01442_, \oc8051_golden_model_1.TH1 [7]);
  and _63747_ (_12108_, _12107_, _43634_);
  and _63748_ (_41507_, _12108_, _12106_);
  not _63749_ (_12109_, _07954_);
  and _63750_ (_12110_, _12109_, \oc8051_golden_model_1.TH0 [7]);
  and _63751_ (_12111_, _09096_, _07954_);
  or _63752_ (_12112_, _12111_, _12110_);
  and _63753_ (_12113_, _12112_, _06615_);
  nor _63754_ (_12114_, _08107_, _12109_);
  or _63755_ (_12115_, _12114_, _12110_);
  or _63756_ (_12116_, _12115_, _06327_);
  and _63757_ (_12117_, _08791_, _07954_);
  or _63758_ (_12118_, _12117_, _12110_);
  or _63759_ (_12119_, _12118_, _07275_);
  and _63760_ (_12120_, _07954_, \oc8051_golden_model_1.ACC [7]);
  or _63761_ (_12121_, _12120_, _12110_);
  and _63762_ (_12122_, _12121_, _07259_);
  and _63763_ (_12123_, _07260_, \oc8051_golden_model_1.TH0 [7]);
  or _63764_ (_12124_, _12123_, _06474_);
  or _63765_ (_12125_, _12124_, _12122_);
  and _63766_ (_12126_, _12125_, _06772_);
  and _63767_ (_12127_, _12126_, _12119_);
  and _63768_ (_12128_, _12115_, _06410_);
  or _63769_ (_12129_, _12128_, _12127_);
  and _63770_ (_12130_, _12129_, _06426_);
  and _63771_ (_12131_, _12121_, _06417_);
  or _63772_ (_12132_, _12131_, _10153_);
  or _63773_ (_12133_, _12132_, _12130_);
  and _63774_ (_12134_, _12133_, _12116_);
  or _63775_ (_12135_, _12134_, _09572_);
  and _63776_ (_12136_, _08778_, _07954_);
  or _63777_ (_12137_, _12110_, _06333_);
  or _63778_ (_12138_, _12137_, _12136_);
  and _63779_ (_12139_, _12138_, _06313_);
  and _63780_ (_12140_, _12139_, _12135_);
  and _63781_ (_12141_, _09076_, _07954_);
  or _63782_ (_12142_, _12141_, _12110_);
  and _63783_ (_12143_, _12142_, _06037_);
  or _63784_ (_12144_, _12143_, _06277_);
  or _63785_ (_12145_, _12144_, _12140_);
  and _63786_ (_12146_, _08880_, _07954_);
  or _63787_ (_12147_, _12146_, _12110_);
  or _63788_ (_12148_, _12147_, _06278_);
  and _63789_ (_12149_, _12148_, _12145_);
  or _63790_ (_12150_, _12149_, _06502_);
  and _63791_ (_12151_, _09090_, _07954_);
  or _63792_ (_12152_, _12110_, _07334_);
  or _63793_ (_12153_, _12152_, _12151_);
  and _63794_ (_12154_, _12153_, _07337_);
  and _63795_ (_12155_, _12154_, _12150_);
  or _63796_ (_12156_, _12155_, _12113_);
  and _63797_ (_12157_, _12156_, _07339_);
  or _63798_ (_12158_, _12110_, _08110_);
  and _63799_ (_12159_, _12147_, _06507_);
  and _63800_ (_12160_, _12159_, _12158_);
  or _63801_ (_12161_, _12160_, _12157_);
  and _63802_ (_12162_, _12161_, _07331_);
  and _63803_ (_12163_, _12121_, _06610_);
  and _63804_ (_12164_, _12163_, _12158_);
  or _63805_ (_12165_, _12164_, _06509_);
  or _63806_ (_12166_, _12165_, _12162_);
  and _63807_ (_12167_, _09087_, _07954_);
  or _63808_ (_12168_, _12110_, _09107_);
  or _63809_ (_12169_, _12168_, _12167_);
  and _63810_ (_12170_, _12169_, _09112_);
  and _63811_ (_12171_, _12170_, _12166_);
  nor _63812_ (_12172_, _09095_, _12109_);
  or _63813_ (_12173_, _12172_, _12110_);
  and _63814_ (_12174_, _12173_, _06602_);
  or _63815_ (_12175_, _12174_, _06639_);
  or _63816_ (_12176_, _12175_, _12171_);
  or _63817_ (_12177_, _12118_, _07048_);
  and _63818_ (_12178_, _12177_, _06651_);
  and _63819_ (_12179_, _12178_, _12176_);
  and _63820_ (_12180_, _08605_, _07954_);
  or _63821_ (_12181_, _12180_, _12110_);
  and _63822_ (_12182_, _12181_, _06646_);
  or _63823_ (_12183_, _12182_, _01446_);
  or _63824_ (_12184_, _12183_, _12179_);
  or _63825_ (_12185_, _01442_, \oc8051_golden_model_1.TH0 [7]);
  and _63826_ (_12186_, _12185_, _43634_);
  and _63827_ (_41508_, _12186_, _12184_);
  not _63828_ (_12187_, _06021_);
  not _63829_ (_12188_, _05685_);
  and _63830_ (_12189_, _08608_, _12188_);
  and _63831_ (_12190_, _12189_, \oc8051_golden_model_1.PC [7]);
  and _63832_ (_12191_, _12190_, \oc8051_golden_model_1.PC [8]);
  and _63833_ (_12192_, _12191_, \oc8051_golden_model_1.PC [9]);
  and _63834_ (_12193_, _12192_, \oc8051_golden_model_1.PC [10]);
  and _63835_ (_12194_, _12193_, \oc8051_golden_model_1.PC [11]);
  and _63836_ (_12195_, _12194_, \oc8051_golden_model_1.PC [12]);
  and _63837_ (_12196_, _12195_, \oc8051_golden_model_1.PC [13]);
  and _63838_ (_12197_, _12196_, \oc8051_golden_model_1.PC [14]);
  or _63839_ (_12198_, _12197_, \oc8051_golden_model_1.PC [15]);
  nand _63840_ (_12199_, _12197_, \oc8051_golden_model_1.PC [15]);
  and _63841_ (_12200_, _12199_, _12198_);
  and _63842_ (_12201_, _11292_, _11248_);
  or _63843_ (_12202_, _12201_, _12200_);
  nand _63844_ (_12203_, _08107_, _06621_);
  nor _63845_ (_12204_, _09540_, \oc8051_golden_model_1.PC [14]);
  nor _63846_ (_12205_, _12204_, _09541_);
  and _63847_ (_12206_, _12205_, _06238_);
  nor _63848_ (_12207_, _12205_, _06238_);
  nor _63849_ (_12208_, _12207_, _12206_);
  nor _63850_ (_12209_, _09539_, \oc8051_golden_model_1.PC [13]);
  nor _63851_ (_12210_, _12209_, _09540_);
  nor _63852_ (_12211_, _12210_, _06238_);
  and _63853_ (_12212_, _12210_, _06238_);
  not _63854_ (_12213_, _12212_);
  nor _63855_ (_12214_, _09538_, \oc8051_golden_model_1.PC [12]);
  nor _63856_ (_12215_, _12214_, _09539_);
  and _63857_ (_12216_, _12215_, _06238_);
  not _63858_ (_12217_, \oc8051_golden_model_1.PC [11]);
  nor _63859_ (_12218_, _09537_, _12217_);
  and _63860_ (_12219_, _09537_, _12217_);
  or _63861_ (_12220_, _12219_, _12218_);
  and _63862_ (_12221_, _12220_, _06238_);
  nor _63863_ (_12222_, _12220_, _06238_);
  nor _63864_ (_12223_, _09543_, \oc8051_golden_model_1.PC [10]);
  nor _63865_ (_12224_, _12223_, _09544_);
  and _63866_ (_12225_, _12224_, _06238_);
  nor _63867_ (_12226_, _12224_, _06238_);
  nor _63868_ (_12227_, _12226_, _12225_);
  and _63869_ (_12228_, _08618_, \oc8051_golden_model_1.PC [8]);
  nor _63870_ (_12229_, _12228_, \oc8051_golden_model_1.PC [9]);
  nor _63871_ (_12230_, _12229_, _09543_);
  and _63872_ (_12231_, _12230_, _06238_);
  nor _63873_ (_12232_, _12230_, _06238_);
  nor _63874_ (_12233_, _08618_, \oc8051_golden_model_1.PC [8]);
  nor _63875_ (_12234_, _12233_, _12228_);
  and _63876_ (_12235_, _12234_, _06238_);
  and _63877_ (_12236_, _08620_, _06238_);
  nor _63878_ (_12237_, _08620_, _06238_);
  and _63879_ (_12238_, _08607_, _06148_);
  nor _63880_ (_12239_, _12238_, \oc8051_golden_model_1.PC [6]);
  nor _63881_ (_12240_, _12239_, _08617_);
  not _63882_ (_12241_, _12240_);
  nor _63883_ (_12242_, _12241_, _06397_);
  and _63884_ (_12243_, _12241_, _06397_);
  nor _63885_ (_12244_, _12243_, _12242_);
  not _63886_ (_12245_, _12244_);
  and _63887_ (_12246_, _06148_, \oc8051_golden_model_1.PC [4]);
  nor _63888_ (_12247_, _12246_, \oc8051_golden_model_1.PC [5]);
  nor _63889_ (_12248_, _12247_, _12238_);
  not _63890_ (_12249_, _12248_);
  nor _63891_ (_12250_, _12249_, _06685_);
  and _63892_ (_12251_, _12249_, _06685_);
  nor _63893_ (_12252_, _06148_, \oc8051_golden_model_1.PC [4]);
  nor _63894_ (_12253_, _12252_, _12246_);
  not _63895_ (_12254_, _12253_);
  nor _63896_ (_12255_, _12254_, _07093_);
  nor _63897_ (_12256_, _06269_, _06521_);
  and _63898_ (_12257_, _06269_, _06521_);
  nor _63899_ (_12258_, _06727_, _06113_);
  nor _63900_ (_12259_, _07127_, \oc8051_golden_model_1.PC [1]);
  nor _63901_ (_12260_, _06310_, _05701_);
  and _63902_ (_12261_, _07127_, \oc8051_golden_model_1.PC [1]);
  nor _63903_ (_12262_, _12261_, _12259_);
  and _63904_ (_12263_, _12262_, _12260_);
  nor _63905_ (_12264_, _12263_, _12259_);
  and _63906_ (_12265_, _06727_, _06113_);
  nor _63907_ (_12266_, _12265_, _12258_);
  not _63908_ (_12267_, _12266_);
  nor _63909_ (_12268_, _12267_, _12264_);
  nor _63910_ (_12269_, _12268_, _12258_);
  nor _63911_ (_12270_, _12269_, _12257_);
  nor _63912_ (_12271_, _12270_, _12256_);
  and _63913_ (_12272_, _12254_, _07093_);
  nor _63914_ (_12273_, _12272_, _12255_);
  not _63915_ (_12274_, _12273_);
  nor _63916_ (_12275_, _12274_, _12271_);
  nor _63917_ (_12276_, _12275_, _12255_);
  nor _63918_ (_12277_, _12276_, _12251_);
  nor _63919_ (_12278_, _12277_, _12250_);
  nor _63920_ (_12279_, _12278_, _12245_);
  nor _63921_ (_12280_, _12279_, _12242_);
  nor _63922_ (_12281_, _12280_, _12237_);
  or _63923_ (_12282_, _12281_, _12236_);
  nor _63924_ (_12283_, _12234_, _06238_);
  nor _63925_ (_12284_, _12283_, _12235_);
  and _63926_ (_12285_, _12284_, _12282_);
  nor _63927_ (_12286_, _12285_, _12235_);
  nor _63928_ (_12287_, _12286_, _12232_);
  nor _63929_ (_12288_, _12287_, _12231_);
  not _63930_ (_12289_, _12288_);
  and _63931_ (_12290_, _12289_, _12227_);
  nor _63932_ (_12291_, _12290_, _12225_);
  nor _63933_ (_12292_, _12291_, _12222_);
  or _63934_ (_12293_, _12292_, _12221_);
  nor _63935_ (_12294_, _12215_, _06238_);
  nor _63936_ (_12295_, _12294_, _12216_);
  and _63937_ (_12296_, _12295_, _12293_);
  nor _63938_ (_12297_, _12296_, _12216_);
  and _63939_ (_12298_, _12297_, _12213_);
  or _63940_ (_12299_, _12298_, _12211_);
  not _63941_ (_12300_, _12299_);
  and _63942_ (_12301_, _12300_, _12208_);
  nor _63943_ (_12302_, _12301_, _12206_);
  nor _63944_ (_12303_, _09550_, _06238_);
  and _63945_ (_12304_, _09550_, _06238_);
  nor _63946_ (_12305_, _12304_, _12303_);
  and _63947_ (_12306_, _12305_, _12302_);
  nor _63948_ (_12307_, _12305_, _12302_);
  or _63949_ (_12308_, _12307_, _12306_);
  or _63950_ (_12309_, _12308_, _10967_);
  and _63951_ (_12310_, _06508_, _05988_);
  or _63952_ (_12311_, _09550_, \oc8051_golden_model_1.PSW [7]);
  and _63953_ (_12312_, _12311_, _12310_);
  and _63954_ (_12313_, _12312_, _12309_);
  nor _63955_ (_12314_, _11114_, _06604_);
  not _63956_ (_12315_, _12314_);
  nor _63957_ (_12316_, _10709_, _06022_);
  not _63958_ (_12317_, _12316_);
  nor _63959_ (_12318_, _06320_, _06022_);
  nor _63960_ (_12319_, _12318_, _06987_);
  and _63961_ (_12320_, _12319_, _12317_);
  or _63962_ (_12321_, _12320_, _12200_);
  nor _63963_ (_12322_, _11089_, _06608_);
  not _63964_ (_12323_, _12322_);
  nor _63965_ (_12324_, _10709_, _06017_);
  not _63966_ (_12325_, _12324_);
  nor _63967_ (_12326_, _06320_, _06017_);
  nor _63968_ (_12327_, _12326_, _06976_);
  and _63969_ (_12328_, _12327_, _12325_);
  or _63970_ (_12329_, _12328_, _12200_);
  nor _63971_ (_12330_, _11064_, _06613_);
  not _63972_ (_12331_, _12330_);
  nor _63973_ (_12332_, _11052_, _11036_);
  and _63974_ (_12333_, _12332_, _11049_);
  or _63975_ (_12334_, _12333_, _12200_);
  and _63976_ (_12335_, _09565_, _06037_);
  nor _63977_ (_12336_, _10623_, _06453_);
  not _63978_ (_12337_, _12336_);
  not _63979_ (_12338_, _10784_);
  nor _63980_ (_12339_, _10853_, _12338_);
  or _63981_ (_12340_, _12339_, _12200_);
  and _63982_ (_12341_, _06443_, _06036_);
  not _63983_ (_12342_, _12341_);
  nor _63984_ (_12343_, _11603_, _09606_);
  and _63985_ (_12344_, _12343_, _12342_);
  not _63986_ (_12345_, _12344_);
  and _63987_ (_12346_, _12345_, _12200_);
  and _63988_ (_12347_, _06344_, _06030_);
  not _63989_ (_12348_, _12347_);
  not _63990_ (_12349_, _06490_);
  or _63991_ (_12350_, _08778_, _06366_);
  and _63992_ (_12351_, _12350_, _08822_);
  or _63993_ (_12352_, _09172_, _06397_);
  nand _63994_ (_12353_, _09172_, _06397_);
  and _63995_ (_12354_, _12353_, _12352_);
  and _63996_ (_12355_, _12354_, _12351_);
  nand _63997_ (_12356_, _09218_, _06685_);
  or _63998_ (_12357_, _09218_, _06685_);
  and _63999_ (_12358_, _12357_, _12356_);
  or _64000_ (_12359_, _09264_, _07093_);
  nand _64001_ (_12360_, _09264_, _07093_);
  and _64002_ (_12361_, _12360_, _12359_);
  and _64003_ (_12362_, _12361_, _12358_);
  and _64004_ (_12363_, _12362_, _12355_);
  or _64005_ (_12364_, _09310_, _06269_);
  or _64006_ (_12365_, _09356_, _06727_);
  nand _64007_ (_12366_, _12365_, _12364_);
  nand _64008_ (_12367_, _09310_, _06269_);
  nand _64009_ (_12368_, _09356_, _06727_);
  nand _64010_ (_12369_, _12368_, _12367_);
  nor _64011_ (_12370_, _12369_, _12366_);
  or _64012_ (_12371_, _09447_, _06310_);
  nand _64013_ (_12372_, _09447_, _06310_);
  or _64014_ (_12373_, _11310_, _07383_);
  or _64015_ (_12374_, _09402_, _07127_);
  and _64016_ (_12375_, _12374_, _12373_);
  and _64017_ (_12376_, _12375_, _12372_);
  and _64018_ (_12377_, _12376_, _12371_);
  and _64019_ (_12378_, _12377_, _12370_);
  nand _64020_ (_12379_, _12378_, _12363_);
  nor _64021_ (_12380_, _09555_, \oc8051_golden_model_1.PC [14]);
  nor _64022_ (_12381_, _12380_, _09556_);
  and _64023_ (_12382_, _12381_, _08880_);
  nor _64024_ (_12383_, _12381_, _08880_);
  nor _64025_ (_12384_, _12383_, _12382_);
  nor _64026_ (_12385_, _09554_, \oc8051_golden_model_1.PC [13]);
  nor _64027_ (_12386_, _12385_, _09555_);
  nor _64028_ (_12387_, _12386_, _08880_);
  and _64029_ (_12388_, _12386_, _08880_);
  not _64030_ (_12389_, _12388_);
  nor _64031_ (_12390_, _09553_, \oc8051_golden_model_1.PC [12]);
  nor _64032_ (_12391_, _12390_, _09554_);
  and _64033_ (_12392_, _12391_, _08880_);
  nor _64034_ (_12393_, _09552_, _12217_);
  and _64035_ (_12394_, _09552_, _12217_);
  or _64036_ (_12395_, _12394_, _12393_);
  not _64037_ (_12396_, _12395_);
  nor _64038_ (_12397_, _12396_, _08879_);
  and _64039_ (_12398_, _12396_, _08879_);
  nor _64040_ (_12399_, _09558_, \oc8051_golden_model_1.PC [10]);
  nor _64041_ (_12400_, _12399_, _09559_);
  not _64042_ (_12401_, _12400_);
  nor _64043_ (_12402_, _12401_, _08879_);
  and _64044_ (_12403_, _12401_, _08879_);
  nor _64045_ (_12404_, _12403_, _12402_);
  and _64046_ (_12405_, _08612_, \oc8051_golden_model_1.PC [8]);
  nor _64047_ (_12406_, _12405_, \oc8051_golden_model_1.PC [9]);
  nor _64048_ (_12407_, _12406_, _09558_);
  not _64049_ (_12408_, _12407_);
  nor _64050_ (_12409_, _12408_, _08879_);
  and _64051_ (_12410_, _12408_, _08879_);
  nor _64052_ (_12411_, _08612_, \oc8051_golden_model_1.PC [8]);
  nor _64053_ (_12412_, _12411_, _12405_);
  not _64054_ (_12413_, _12412_);
  nor _64055_ (_12414_, _12413_, _08879_);
  nor _64056_ (_12415_, _08879_, _08615_);
  and _64057_ (_12416_, _08879_, _08615_);
  and _64058_ (_12417_, _08610_, _08607_);
  nor _64059_ (_12418_, _12417_, \oc8051_golden_model_1.PC [6]);
  nor _64060_ (_12419_, _12418_, _08611_);
  not _64061_ (_12420_, _12419_);
  nor _64062_ (_12421_, _12420_, _08918_);
  and _64063_ (_12422_, _12420_, _08918_);
  nor _64064_ (_12423_, _12422_, _12421_);
  not _64065_ (_12424_, _12423_);
  and _64066_ (_12425_, _08610_, \oc8051_golden_model_1.PC [4]);
  nor _64067_ (_12426_, _12425_, \oc8051_golden_model_1.PC [5]);
  nor _64068_ (_12427_, _12426_, _12417_);
  not _64069_ (_12428_, _12427_);
  nor _64070_ (_12429_, _12428_, _08953_);
  and _64071_ (_12430_, _12428_, _08953_);
  nor _64072_ (_12431_, _08610_, \oc8051_golden_model_1.PC [4]);
  nor _64073_ (_12432_, _12431_, _12425_);
  not _64074_ (_12433_, _12432_);
  nor _64075_ (_12434_, _12433_, _08986_);
  nor _64076_ (_12435_, _08609_, \oc8051_golden_model_1.PC [3]);
  nor _64077_ (_12436_, _12435_, _08610_);
  not _64078_ (_12437_, _12436_);
  nor _64079_ (_12438_, _12437_, _06595_);
  and _64080_ (_12439_, _12437_, _06595_);
  nor _64081_ (_12440_, _05705_, \oc8051_golden_model_1.PC [2]);
  nor _64082_ (_12441_, _12440_, _08609_);
  not _64083_ (_12442_, _12441_);
  nor _64084_ (_12443_, _12442_, _06769_);
  not _64085_ (_12444_, _06089_);
  nor _64086_ (_12445_, _07160_, _12444_);
  nor _64087_ (_12446_, _06950_, \oc8051_golden_model_1.PC [0]);
  and _64088_ (_12447_, _07160_, _12444_);
  nor _64089_ (_12448_, _12447_, _12445_);
  and _64090_ (_12449_, _12448_, _12446_);
  nor _64091_ (_12450_, _12449_, _12445_);
  and _64092_ (_12451_, _12442_, _06769_);
  nor _64093_ (_12452_, _12451_, _12443_);
  not _64094_ (_12453_, _12452_);
  nor _64095_ (_12454_, _12453_, _12450_);
  nor _64096_ (_12455_, _12454_, _12443_);
  nor _64097_ (_12456_, _12455_, _12439_);
  nor _64098_ (_12457_, _12456_, _12438_);
  and _64099_ (_12458_, _12433_, _08986_);
  nor _64100_ (_12459_, _12458_, _12434_);
  not _64101_ (_12460_, _12459_);
  nor _64102_ (_12461_, _12460_, _12457_);
  nor _64103_ (_12462_, _12461_, _12434_);
  nor _64104_ (_12463_, _12462_, _12430_);
  nor _64105_ (_12464_, _12463_, _12429_);
  nor _64106_ (_12465_, _12464_, _12424_);
  nor _64107_ (_12466_, _12465_, _12421_);
  nor _64108_ (_12467_, _12466_, _12416_);
  or _64109_ (_12468_, _12467_, _12415_);
  and _64110_ (_12469_, _12413_, _08879_);
  nor _64111_ (_12470_, _12469_, _12414_);
  and _64112_ (_12471_, _12470_, _12468_);
  nor _64113_ (_12472_, _12471_, _12414_);
  nor _64114_ (_12473_, _12472_, _12410_);
  nor _64115_ (_12474_, _12473_, _12409_);
  not _64116_ (_12475_, _12474_);
  and _64117_ (_12476_, _12475_, _12404_);
  nor _64118_ (_12477_, _12476_, _12402_);
  nor _64119_ (_12478_, _12477_, _12398_);
  or _64120_ (_12479_, _12478_, _12397_);
  nor _64121_ (_12480_, _12391_, _08880_);
  nor _64122_ (_12481_, _12480_, _12392_);
  and _64123_ (_12482_, _12481_, _12479_);
  nor _64124_ (_12483_, _12482_, _12392_);
  and _64125_ (_12484_, _12483_, _12389_);
  or _64126_ (_12485_, _12484_, _12387_);
  not _64127_ (_12486_, _12485_);
  and _64128_ (_12487_, _12486_, _12384_);
  nor _64129_ (_12488_, _12487_, _12382_);
  not _64130_ (_12489_, _09565_);
  and _64131_ (_12490_, _12489_, _08879_);
  nor _64132_ (_12491_, _12489_, _08879_);
  nor _64133_ (_12492_, _12491_, _12490_);
  and _64134_ (_12493_, _12492_, _12488_);
  nor _64135_ (_12494_, _12492_, _12488_);
  or _64136_ (_12495_, _12494_, _12493_);
  and _64137_ (_12496_, _12495_, _12379_);
  nor _64138_ (_12497_, _12379_, _12489_);
  or _64139_ (_12498_, _12497_, _12496_);
  or _64140_ (_12499_, _12498_, _06473_);
  and _64141_ (_12500_, _09550_, _06417_);
  and _64142_ (_12501_, _06355_, _06030_);
  nor _64143_ (_12502_, _12501_, _10729_);
  and _64144_ (_12503_, _12502_, _07270_);
  not _64145_ (_12504_, _12503_);
  and _64146_ (_12505_, _12504_, _12200_);
  and _64147_ (_12506_, _08453_, _08403_);
  and _64148_ (_12507_, _08785_, _12506_);
  and _64149_ (_12508_, _08211_, _08109_);
  and _64150_ (_12509_, _12508_, _08783_);
  nand _64151_ (_12510_, _12509_, _12507_);
  or _64152_ (_12511_, _12510_, _09565_);
  and _64153_ (_12512_, _12509_, _12507_);
  or _64154_ (_12513_, _12512_, _12495_);
  and _64155_ (_12514_, _12513_, _06474_);
  and _64156_ (_12515_, _12514_, _12511_);
  and _64157_ (_12516_, _10714_, _06062_);
  not _64158_ (_12517_, _06855_);
  nor _64159_ (_12518_, _07576_, _07560_);
  and _64160_ (_12519_, _12518_, _12517_);
  and _64161_ (_12520_, _12519_, _12516_);
  or _64162_ (_12521_, _12520_, _12200_);
  not _64163_ (_12522_, _09550_);
  or _64164_ (_12523_, _07259_, _06816_);
  and _64165_ (_12524_, _12523_, _12522_);
  nor _64166_ (_12525_, _06855_, _07259_);
  nor _64167_ (_12526_, _06816_, \oc8051_golden_model_1.PC [15]);
  and _64168_ (_12527_, _12526_, _12525_);
  and _64169_ (_12528_, _12527_, _12518_);
  or _64170_ (_12529_, _12528_, _12524_);
  nand _64171_ (_12530_, _12529_, _12516_);
  and _64172_ (_12531_, _12530_, _08685_);
  and _64173_ (_12532_, _12531_, _12521_);
  and _64174_ (_12533_, _08209_, _08107_);
  and _64175_ (_12534_, _12533_, _08675_);
  and _64176_ (_12535_, _07448_, _07250_);
  and _64177_ (_12536_, _12535_, _08676_);
  nand _64178_ (_12537_, _12536_, _12534_);
  and _64179_ (_12538_, _12537_, _12308_);
  and _64180_ (_12539_, _12536_, _12534_);
  and _64181_ (_12540_, _12539_, _09550_);
  or _64182_ (_12541_, _12540_, _12538_);
  and _64183_ (_12542_, _12541_, _08687_);
  or _64184_ (_12543_, _12542_, _12532_);
  nor _64185_ (_12544_, _07269_, _06474_);
  and _64186_ (_12545_, _12544_, _12543_);
  or _64187_ (_12546_, _12545_, _12515_);
  and _64188_ (_12547_, _12546_, _12502_);
  or _64189_ (_12548_, _12547_, _12505_);
  and _64190_ (_12549_, _06418_, _06052_);
  and _64191_ (_12550_, _12549_, _12548_);
  nor _64192_ (_12551_, _10696_, _07289_);
  not _64193_ (_12552_, _12551_);
  nor _64194_ (_12553_, _12549_, _12522_);
  or _64195_ (_12554_, _12553_, _12552_);
  or _64196_ (_12555_, _12554_, _12550_);
  or _64197_ (_12556_, _12551_, _12200_);
  and _64198_ (_12557_, _12556_, _06426_);
  and _64199_ (_12558_, _12557_, _12555_);
  or _64200_ (_12559_, _12558_, _12500_);
  and _64201_ (_12560_, _06350_, _06030_);
  nor _64202_ (_12561_, _12560_, _10694_);
  and _64203_ (_12562_, _12561_, _12559_);
  not _64204_ (_12563_, _12561_);
  and _64205_ (_12564_, _12563_, _12200_);
  not _64206_ (_12565_, _06057_);
  nor _64207_ (_12566_, _06351_, _12565_);
  and _64208_ (_12567_, _12566_, _06353_);
  not _64209_ (_12568_, _12567_);
  or _64210_ (_12569_, _12568_, _12564_);
  or _64211_ (_12570_, _12569_, _12562_);
  not _64212_ (_12571_, _06469_);
  nor _64213_ (_12572_, _06320_, _06048_);
  nor _64214_ (_12573_, _12572_, _06483_);
  and _64215_ (_12574_, _12573_, _12571_);
  or _64216_ (_12575_, _12567_, _09550_);
  and _64217_ (_12576_, _12575_, _12574_);
  and _64218_ (_12577_, _12576_, _12570_);
  not _64219_ (_12578_, _08108_);
  and _64220_ (_12579_, _08107_, _06238_);
  nor _64221_ (_12580_, _12579_, _12578_);
  and _64222_ (_12581_, _08209_, _07741_);
  nor _64223_ (_12582_, _08209_, _07741_);
  nor _64224_ (_12583_, _12582_, _12581_);
  and _64225_ (_12584_, _12583_, _12580_);
  or _64226_ (_12585_, _08305_, _07983_);
  and _64227_ (_12586_, _08305_, _07983_);
  not _64228_ (_12587_, _12586_);
  and _64229_ (_12588_, _12587_, _12585_);
  nor _64230_ (_12589_, _08596_, _07959_);
  and _64231_ (_12590_, _08596_, _07959_);
  nor _64232_ (_12591_, _12590_, _12589_);
  and _64233_ (_12592_, _12591_, _12588_);
  and _64234_ (_12593_, _12592_, _12584_);
  and _64235_ (_12594_, _07680_, _06622_);
  and _64236_ (_12595_, _07854_, _07799_);
  or _64237_ (_12596_, _12595_, _12594_);
  or _64238_ (_12597_, _07680_, _06622_);
  or _64239_ (_12598_, _07854_, _07799_);
  nand _64240_ (_12599_, _12598_, _12597_);
  nor _64241_ (_12600_, _12599_, _12596_);
  nand _64242_ (_12601_, _07250_, _06310_);
  nor _64243_ (_12602_, _07448_, _07383_);
  and _64244_ (_12603_, _07448_, _07383_);
  nor _64245_ (_12604_, _12603_, _12602_);
  and _64246_ (_12605_, _12604_, _12601_);
  and _64247_ (_12606_, _12605_, _12600_);
  or _64248_ (_12607_, _07250_, _06310_);
  and _64249_ (_12608_, _12607_, _12606_);
  and _64250_ (_12609_, _12608_, _12593_);
  nand _64251_ (_12610_, _12609_, _12489_);
  not _64252_ (_12611_, _12574_);
  or _64253_ (_12612_, _12609_, _12495_);
  and _64254_ (_12613_, _12612_, _12611_);
  and _64255_ (_12614_, _12613_, _12610_);
  or _64256_ (_12615_, _12614_, _06472_);
  or _64257_ (_12616_, _12615_, _12577_);
  and _64258_ (_12617_, _12616_, _06500_);
  and _64259_ (_12618_, _12617_, _12499_);
  nor _64260_ (_12619_, _10574_, _10573_);
  nor _64261_ (_12620_, _12619_, _10583_);
  not _64262_ (_12621_, _10579_);
  nor _64263_ (_12622_, _08453_, \oc8051_golden_model_1.ACC [0]);
  or _64264_ (_12623_, _12622_, _10577_);
  and _64265_ (_12624_, _12623_, _12621_);
  and _64266_ (_12625_, _12624_, _12620_);
  nor _64267_ (_12626_, _10569_, _10570_);
  nor _64268_ (_12627_, _12626_, _10590_);
  nor _64269_ (_12628_, _10596_, _09096_);
  and _64270_ (_12629_, _12628_, _12627_);
  and _64271_ (_12630_, _12629_, _12625_);
  and _64272_ (_12631_, _12630_, _09565_);
  not _64273_ (_12632_, _12630_);
  and _64274_ (_12633_, _12632_, _12495_);
  or _64275_ (_12634_, _12633_, _12631_);
  and _64276_ (_12635_, _12634_, _06431_);
  or _64277_ (_12636_, _12635_, _12618_);
  and _64278_ (_12637_, _12636_, _12349_);
  nor _64279_ (_12638_, _11345_, _11346_);
  nor _64280_ (_12639_, _12638_, _11349_);
  and _64281_ (_12640_, _06310_, _06071_);
  nor _64282_ (_12641_, _12640_, _11351_);
  nor _64283_ (_12642_, _11355_, _12641_);
  and _64284_ (_12643_, _12642_, _12639_);
  nor _64285_ (_12644_, _11339_, _11340_);
  nor _64286_ (_12645_, _12644_, _11344_);
  nor _64287_ (_12646_, _11338_, _11070_);
  and _64288_ (_12647_, _12646_, _12645_);
  and _64289_ (_12648_, _12647_, _12643_);
  or _64290_ (_12649_, _12648_, _12495_);
  nand _64291_ (_12650_, _12648_, _12489_);
  and _64292_ (_12651_, _12650_, _06490_);
  and _64293_ (_12652_, _12651_, _12649_);
  or _64294_ (_12653_, _12652_, _12637_);
  and _64295_ (_12654_, _12653_, _12348_);
  nand _64296_ (_12655_, _12347_, _12200_);
  nor _64297_ (_12656_, _07309_, _07596_);
  and _64298_ (_12657_, _12656_, _06346_);
  and _64299_ (_12658_, _06785_, _06443_);
  nor _64300_ (_12659_, _12658_, _06404_);
  nor _64301_ (_12660_, _07889_, _07487_);
  and _64302_ (_12661_, _12660_, _12659_);
  and _64303_ (_12662_, _12661_, _12657_);
  nand _64304_ (_12663_, _12662_, _12655_);
  or _64305_ (_12664_, _12663_, _12654_);
  or _64306_ (_12665_, _12662_, _09550_);
  and _64307_ (_12666_, _12665_, _12344_);
  and _64308_ (_12667_, _12666_, _12664_);
  or _64309_ (_12668_, _12667_, _12346_);
  and _64310_ (_12669_, _06446_, _06055_);
  and _64311_ (_12670_, _12669_, _12668_);
  not _64312_ (_12671_, _12339_);
  nor _64313_ (_12672_, _12669_, _12522_);
  or _64314_ (_12673_, _12672_, _12671_);
  or _64315_ (_12674_, _12673_, _12670_);
  and _64316_ (_12675_, _12674_, _12340_);
  or _64317_ (_12676_, _12675_, _12337_);
  or _64318_ (_12677_, _12336_, _09550_);
  and _64319_ (_12678_, _12677_, _06043_);
  and _64320_ (_12679_, _12678_, _12676_);
  nand _64321_ (_12680_, _12200_, _06042_);
  nor _64322_ (_12681_, _06339_, _06039_);
  nand _64323_ (_12682_, _12681_, _12680_);
  or _64324_ (_12683_, _12682_, _12679_);
  or _64325_ (_12684_, _12681_, _09550_);
  and _64326_ (_12685_, _12684_, _06487_);
  and _64327_ (_12686_, _12685_, _12683_);
  nand _64328_ (_12687_, _09565_, _06486_);
  nand _64329_ (_12688_, _12687_, _06334_);
  or _64330_ (_12689_, _12688_, _12686_);
  or _64331_ (_12690_, _09550_, _06334_);
  and _64332_ (_12691_, _12690_, _06313_);
  and _64333_ (_12692_, _12691_, _12689_);
  or _64334_ (_12693_, _12692_, _12335_);
  nor _64335_ (_12694_, _10166_, _06031_);
  and _64336_ (_12695_, _12694_, _12693_);
  not _64337_ (_12696_, _06004_);
  nor _64338_ (_12697_, _06401_, _12696_);
  not _64339_ (_12698_, _12697_);
  not _64340_ (_12700_, _12694_);
  and _64341_ (_12701_, _12700_, _12200_);
  or _64342_ (_12702_, _12701_, _12698_);
  or _64343_ (_12703_, _12702_, _12695_);
  and _64344_ (_12704_, _06002_, _05988_);
  not _64345_ (_12705_, _12704_);
  or _64346_ (_12706_, _12697_, _09550_);
  and _64347_ (_12707_, _12706_, _12705_);
  and _64348_ (_12708_, _12707_, _12703_);
  and _64349_ (_12709_, _12704_, _12308_);
  or _64350_ (_12710_, _12709_, _08848_);
  or _64351_ (_12711_, _12710_, _12708_);
  and _64352_ (_12712_, _09550_, _06278_);
  or _64353_ (_12713_, _12712_, _08627_);
  and _64354_ (_12714_, _12713_, _12711_);
  and _64355_ (_12715_, _09565_, _06277_);
  or _64356_ (_12716_, _12715_, _11028_);
  or _64357_ (_12717_, _12716_, _12714_);
  and _64358_ (_12718_, _06030_, _06276_);
  not _64359_ (_12719_, _12718_);
  or _64360_ (_12721_, _11029_, _09550_);
  and _64361_ (_12722_, _12721_, _12719_);
  and _64362_ (_12723_, _12722_, _12717_);
  nor _64363_ (_12724_, _06400_, _06275_);
  not _64364_ (_12725_, _12724_);
  not _64365_ (_12726_, \oc8051_golden_model_1.DPH [0]);
  and _64366_ (_12727_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _64367_ (_12728_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _64368_ (_12729_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _64369_ (_12730_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _64370_ (_12731_, _12730_, _12729_);
  not _64371_ (_12732_, _12731_);
  and _64372_ (_12733_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _64373_ (_12734_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _64374_ (_12735_, _12734_, _12733_);
  not _64375_ (_12736_, _12735_);
  and _64376_ (_12737_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _64377_ (_12738_, _06168_, _06164_);
  nor _64378_ (_12739_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _64379_ (_12740_, _12739_, _12737_);
  not _64380_ (_12741_, _12740_);
  nor _64381_ (_12742_, _12741_, _12738_);
  nor _64382_ (_12743_, _12742_, _12737_);
  nor _64383_ (_12744_, _12743_, _12736_);
  nor _64384_ (_12745_, _12744_, _12733_);
  nor _64385_ (_12746_, _12745_, _12732_);
  nor _64386_ (_12747_, _12746_, _12729_);
  nor _64387_ (_12748_, _12747_, _12728_);
  nor _64388_ (_12749_, _12748_, _12727_);
  nor _64389_ (_12750_, _12749_, _12726_);
  and _64390_ (_12751_, _12750_, \oc8051_golden_model_1.DPH [1]);
  and _64391_ (_12752_, _12751_, \oc8051_golden_model_1.DPH [2]);
  and _64392_ (_12753_, _12752_, \oc8051_golden_model_1.DPH [3]);
  and _64393_ (_12754_, _12753_, \oc8051_golden_model_1.DPH [4]);
  and _64394_ (_12755_, _12754_, \oc8051_golden_model_1.DPH [5]);
  and _64395_ (_12756_, _12755_, \oc8051_golden_model_1.DPH [6]);
  nand _64396_ (_12757_, _12756_, \oc8051_golden_model_1.DPH [7]);
  or _64397_ (_12758_, _12756_, \oc8051_golden_model_1.DPH [7]);
  and _64398_ (_12759_, _12758_, _12718_);
  and _64399_ (_12760_, _12759_, _12757_);
  or _64400_ (_12761_, _12760_, _12725_);
  or _64401_ (_12762_, _12761_, _12723_);
  and _64402_ (_12763_, _06276_, _05988_);
  not _64403_ (_12764_, _12763_);
  or _64404_ (_12765_, _12724_, _09550_);
  and _64405_ (_12766_, _12765_, _12764_);
  and _64406_ (_12767_, _12766_, _12762_);
  not _64407_ (_12768_, _12333_);
  or _64408_ (_12769_, _12308_, _11389_);
  not _64409_ (_12770_, _11389_);
  or _64410_ (_12771_, _12770_, _09550_);
  and _64411_ (_12772_, _12771_, _12763_);
  and _64412_ (_12773_, _12772_, _12769_);
  or _64413_ (_12774_, _12773_, _12768_);
  or _64414_ (_12775_, _12774_, _12767_);
  and _64415_ (_12776_, _12775_, _12334_);
  or _64416_ (_12777_, _12776_, _12331_);
  or _64417_ (_12778_, _12330_, _09550_);
  and _64418_ (_12779_, _12778_, _07334_);
  and _64419_ (_12780_, _12779_, _12777_);
  and _64420_ (_12781_, _09565_, _06502_);
  not _64421_ (_12782_, _06012_);
  nor _64422_ (_12783_, _06615_, _12782_);
  not _64423_ (_12784_, _12783_);
  or _64424_ (_12785_, _12784_, _12781_);
  or _64425_ (_12786_, _12785_, _12780_);
  and _64426_ (_12787_, _06501_, _05988_);
  not _64427_ (_12788_, _12787_);
  or _64428_ (_12789_, _12783_, _09550_);
  and _64429_ (_12790_, _12789_, _12788_);
  and _64430_ (_12791_, _12790_, _12786_);
  not _64431_ (_12792_, _12328_);
  or _64432_ (_12793_, _12308_, _12770_);
  or _64433_ (_12794_, _11389_, _09550_);
  and _64434_ (_12795_, _12794_, _12787_);
  and _64435_ (_12796_, _12795_, _12793_);
  or _64436_ (_12797_, _12796_, _12792_);
  or _64437_ (_12798_, _12797_, _12791_);
  and _64438_ (_12799_, _12798_, _12329_);
  or _64439_ (_12800_, _12799_, _12323_);
  or _64440_ (_12801_, _12322_, _09550_);
  and _64441_ (_12802_, _12801_, _07339_);
  and _64442_ (_12803_, _12802_, _12800_);
  and _64443_ (_12804_, _09565_, _06507_);
  nor _64444_ (_12805_, _06610_, _07330_);
  not _64445_ (_12806_, _12805_);
  or _64446_ (_12807_, _12806_, _12804_);
  or _64447_ (_12808_, _12807_, _12803_);
  and _64448_ (_12809_, _06506_, _05988_);
  not _64449_ (_12810_, _12809_);
  or _64450_ (_12811_, _12805_, _09550_);
  and _64451_ (_12812_, _12811_, _12810_);
  and _64452_ (_12813_, _12812_, _12808_);
  not _64453_ (_12814_, _12320_);
  or _64454_ (_12815_, _12308_, \oc8051_golden_model_1.PSW [7]);
  or _64455_ (_12816_, _09550_, _10967_);
  and _64456_ (_12817_, _12816_, _12809_);
  and _64457_ (_12818_, _12817_, _12815_);
  or _64458_ (_12819_, _12818_, _12814_);
  or _64459_ (_12820_, _12819_, _12813_);
  and _64460_ (_12821_, _12820_, _12321_);
  or _64461_ (_12822_, _12821_, _12315_);
  or _64462_ (_12823_, _12314_, _09550_);
  and _64463_ (_12824_, _12823_, _09107_);
  and _64464_ (_12825_, _12824_, _12822_);
  and _64465_ (_12826_, _09565_, _06509_);
  not _64466_ (_12827_, _06023_);
  nor _64467_ (_12828_, _06602_, _12827_);
  not _64468_ (_12829_, _12828_);
  or _64469_ (_12830_, _12829_, _12826_);
  or _64470_ (_12831_, _12830_, _12825_);
  not _64471_ (_12832_, _12310_);
  or _64472_ (_12833_, _12828_, _09550_);
  and _64473_ (_12834_, _12833_, _12832_);
  and _64474_ (_12835_, _12834_, _12831_);
  or _64475_ (_12836_, _12835_, _12313_);
  and _64476_ (_12837_, _11158_, _11127_);
  and _64477_ (_12838_, _12837_, _12836_);
  not _64478_ (_12839_, _12837_);
  and _64479_ (_12840_, _12839_, _12200_);
  or _64480_ (_12841_, _12840_, _11188_);
  or _64481_ (_12842_, _12841_, _12838_);
  or _64482_ (_12843_, _11187_, _09550_);
  and _64483_ (_12844_, _12843_, _11217_);
  and _64484_ (_12845_, _12844_, _12842_);
  and _64485_ (_12846_, _12200_, _11216_);
  or _64486_ (_12847_, _12846_, _06621_);
  or _64487_ (_12848_, _12847_, _12845_);
  and _64488_ (_12849_, _12848_, _12203_);
  or _64489_ (_12850_, _12849_, _07350_);
  or _64490_ (_12851_, _09550_, _06016_);
  and _64491_ (_12852_, _12851_, _06629_);
  and _64492_ (_12853_, _12852_, _12850_);
  not _64493_ (_12854_, _12201_);
  not _64494_ (_12855_, _08000_);
  and _64495_ (_12856_, _08633_, \oc8051_golden_model_1.TCON [2]);
  and _64496_ (_12857_, _08645_, \oc8051_golden_model_1.ACC [2]);
  nor _64497_ (_12858_, _12857_, _12856_);
  and _64498_ (_12859_, _08643_, \oc8051_golden_model_1.IP [2]);
  not _64499_ (_12860_, _12859_);
  and _64500_ (_12861_, _08640_, \oc8051_golden_model_1.PSW [2]);
  and _64501_ (_12862_, _08637_, \oc8051_golden_model_1.B [2]);
  nor _64502_ (_12863_, _12862_, _12861_);
  and _64503_ (_12864_, _12863_, _12860_);
  and _64504_ (_12865_, _12864_, _12858_);
  and _64505_ (_12866_, _08650_, \oc8051_golden_model_1.SCON [2]);
  and _64506_ (_12867_, _08652_, \oc8051_golden_model_1.IE [2]);
  nor _64507_ (_12868_, _12867_, _12866_);
  and _64508_ (_12869_, _08655_, \oc8051_golden_model_1.P2INREG [2]);
  and _64509_ (_12870_, _08657_, \oc8051_golden_model_1.P3INREG [2]);
  nor _64510_ (_12871_, _12870_, _12869_);
  and _64511_ (_12872_, _07993_, \oc8051_golden_model_1.P0INREG [2]);
  and _64512_ (_12873_, _08661_, \oc8051_golden_model_1.P1INREG [2]);
  nor _64513_ (_12874_, _12873_, _12872_);
  and _64514_ (_12875_, _12874_, _12871_);
  and _64515_ (_12876_, _12875_, _12868_);
  and _64516_ (_12877_, _12876_, _12865_);
  and _64517_ (_12878_, _12877_, _08501_);
  nor _64518_ (_12879_, _12878_, _12855_);
  not _64519_ (_12880_, _07957_);
  and _64520_ (_12881_, _07993_, \oc8051_golden_model_1.P0INREG [1]);
  and _64521_ (_12882_, _08661_, \oc8051_golden_model_1.P1INREG [1]);
  nor _64522_ (_12883_, _12882_, _12881_);
  and _64523_ (_12884_, _08650_, \oc8051_golden_model_1.SCON [1]);
  and _64524_ (_12885_, _08652_, \oc8051_golden_model_1.IE [1]);
  nor _64525_ (_12886_, _12885_, _12884_);
  and _64526_ (_12887_, _08643_, \oc8051_golden_model_1.IP [1]);
  and _64527_ (_12888_, _08637_, \oc8051_golden_model_1.B [1]);
  nor _64528_ (_12889_, _12888_, _12887_);
  and _64529_ (_12890_, _08640_, \oc8051_golden_model_1.PSW [1]);
  and _64530_ (_12891_, _08645_, \oc8051_golden_model_1.ACC [1]);
  nor _64531_ (_12892_, _12891_, _12890_);
  and _64532_ (_12893_, _12892_, _12889_);
  and _64533_ (_12894_, _08633_, \oc8051_golden_model_1.TCON [1]);
  and _64534_ (_12895_, _08657_, \oc8051_golden_model_1.P3INREG [1]);
  and _64535_ (_12896_, _08655_, \oc8051_golden_model_1.P2INREG [1]);
  or _64536_ (_12897_, _12896_, _12895_);
  nor _64537_ (_12898_, _12897_, _12894_);
  and _64538_ (_12899_, _12898_, _12893_);
  and _64539_ (_12900_, _12899_, _12886_);
  and _64540_ (_12901_, _12900_, _12883_);
  and _64541_ (_12902_, _12901_, _08402_);
  nor _64542_ (_12903_, _12902_, _12880_);
  nor _64543_ (_12904_, _12903_, _12879_);
  and _64544_ (_12905_, _08633_, \oc8051_golden_model_1.TCON [4]);
  and _64545_ (_12906_, _08645_, \oc8051_golden_model_1.ACC [4]);
  nor _64546_ (_12907_, _12906_, _12905_);
  and _64547_ (_12908_, _08640_, \oc8051_golden_model_1.PSW [4]);
  not _64548_ (_12909_, _12908_);
  and _64549_ (_12910_, _08643_, \oc8051_golden_model_1.IP [4]);
  and _64550_ (_12911_, _08637_, \oc8051_golden_model_1.B [4]);
  nor _64551_ (_12912_, _12911_, _12910_);
  and _64552_ (_12913_, _12912_, _12909_);
  and _64553_ (_12914_, _12913_, _12907_);
  and _64554_ (_12915_, _08650_, \oc8051_golden_model_1.SCON [4]);
  and _64555_ (_12916_, _08652_, \oc8051_golden_model_1.IE [4]);
  nor _64556_ (_12917_, _12916_, _12915_);
  and _64557_ (_12918_, _08655_, \oc8051_golden_model_1.P2INREG [4]);
  and _64558_ (_12919_, _08657_, \oc8051_golden_model_1.P3INREG [4]);
  nor _64559_ (_12920_, _12919_, _12918_);
  and _64560_ (_12921_, _07993_, \oc8051_golden_model_1.P0INREG [4]);
  and _64561_ (_12922_, _08661_, \oc8051_golden_model_1.P1INREG [4]);
  nor _64562_ (_12923_, _12922_, _12921_);
  and _64563_ (_12924_, _12923_, _12920_);
  and _64564_ (_12925_, _12924_, _12917_);
  and _64565_ (_12926_, _12925_, _12914_);
  and _64566_ (_12927_, _12926_, _08597_);
  and _64567_ (_12928_, _07950_, _07799_);
  not _64568_ (_12929_, _12928_);
  nor _64569_ (_12930_, _12929_, _12927_);
  nor _64570_ (_12931_, _12930_, _08808_);
  and _64571_ (_12932_, _12931_, _12904_);
  not _64572_ (_12933_, _07967_);
  and _64573_ (_12934_, _07993_, \oc8051_golden_model_1.P0INREG [0]);
  and _64574_ (_12935_, _08661_, \oc8051_golden_model_1.P1INREG [0]);
  nor _64575_ (_12936_, _12935_, _12934_);
  and _64576_ (_12937_, _08650_, \oc8051_golden_model_1.SCON [0]);
  and _64577_ (_12938_, _08652_, \oc8051_golden_model_1.IE [0]);
  nor _64578_ (_12939_, _12938_, _12937_);
  and _64579_ (_12940_, _08640_, \oc8051_golden_model_1.PSW [0]);
  and _64580_ (_12941_, _08645_, \oc8051_golden_model_1.ACC [0]);
  nor _64581_ (_12942_, _12941_, _12940_);
  and _64582_ (_12943_, _08643_, \oc8051_golden_model_1.IP [0]);
  and _64583_ (_12944_, _08637_, \oc8051_golden_model_1.B [0]);
  nor _64584_ (_12945_, _12944_, _12943_);
  and _64585_ (_12946_, _12945_, _12942_);
  and _64586_ (_12947_, _08633_, \oc8051_golden_model_1.TCON [0]);
  and _64587_ (_12948_, _08657_, \oc8051_golden_model_1.P3INREG [0]);
  and _64588_ (_12949_, _08655_, \oc8051_golden_model_1.P2INREG [0]);
  or _64589_ (_12950_, _12949_, _12948_);
  nor _64590_ (_12951_, _12950_, _12947_);
  and _64591_ (_12952_, _12951_, _12946_);
  and _64592_ (_12953_, _12952_, _12939_);
  and _64593_ (_12954_, _12953_, _12936_);
  and _64594_ (_12955_, _12954_, _08452_);
  nor _64595_ (_12956_, _12955_, _12933_);
  and _64596_ (_12957_, _08633_, \oc8051_golden_model_1.TCON [6]);
  and _64597_ (_12958_, _08637_, \oc8051_golden_model_1.B [6]);
  nor _64598_ (_12959_, _12958_, _12957_);
  and _64599_ (_12960_, _08643_, \oc8051_golden_model_1.IP [6]);
  not _64600_ (_12961_, _12960_);
  and _64601_ (_12962_, _08640_, \oc8051_golden_model_1.PSW [6]);
  and _64602_ (_12963_, _08645_, \oc8051_golden_model_1.ACC [6]);
  nor _64603_ (_12964_, _12963_, _12962_);
  and _64604_ (_12965_, _12964_, _12961_);
  and _64605_ (_12966_, _12965_, _12959_);
  and _64606_ (_12967_, _08650_, \oc8051_golden_model_1.SCON [6]);
  and _64607_ (_12968_, _08652_, \oc8051_golden_model_1.IE [6]);
  nor _64608_ (_12969_, _12968_, _12967_);
  and _64609_ (_12970_, _08655_, \oc8051_golden_model_1.P2INREG [6]);
  and _64610_ (_12971_, _08657_, \oc8051_golden_model_1.P3INREG [6]);
  nor _64611_ (_12972_, _12971_, _12970_);
  and _64612_ (_12973_, _07993_, \oc8051_golden_model_1.P0INREG [6]);
  and _64613_ (_12974_, _08661_, \oc8051_golden_model_1.P1INREG [6]);
  nor _64614_ (_12975_, _12974_, _12973_);
  and _64615_ (_12976_, _12975_, _12972_);
  and _64616_ (_12977_, _12976_, _12969_);
  and _64617_ (_12978_, _12977_, _12966_);
  and _64618_ (_12979_, _12978_, _08210_);
  and _64619_ (_12980_, _07973_, _07799_);
  not _64620_ (_12981_, _12980_);
  nor _64621_ (_12982_, _12981_, _12979_);
  nor _64622_ (_12983_, _12982_, _12956_);
  not _64623_ (_12984_, _07994_);
  and _64624_ (_12985_, _08633_, \oc8051_golden_model_1.TCON [3]);
  and _64625_ (_12986_, _08637_, \oc8051_golden_model_1.B [3]);
  nor _64626_ (_12987_, _12986_, _12985_);
  and _64627_ (_12988_, _08640_, \oc8051_golden_model_1.PSW [3]);
  not _64628_ (_12989_, _12988_);
  and _64629_ (_12990_, _08643_, \oc8051_golden_model_1.IP [3]);
  and _64630_ (_12991_, _08645_, \oc8051_golden_model_1.ACC [3]);
  nor _64631_ (_12992_, _12991_, _12990_);
  and _64632_ (_12993_, _12992_, _12989_);
  and _64633_ (_12994_, _12993_, _12987_);
  and _64634_ (_12995_, _08650_, \oc8051_golden_model_1.SCON [3]);
  and _64635_ (_12996_, _08652_, \oc8051_golden_model_1.IE [3]);
  nor _64636_ (_12997_, _12996_, _12995_);
  and _64637_ (_12998_, _08655_, \oc8051_golden_model_1.P2INREG [3]);
  and _64638_ (_12999_, _08657_, \oc8051_golden_model_1.P3INREG [3]);
  nor _64639_ (_13000_, _12999_, _12998_);
  and _64640_ (_13001_, _07993_, \oc8051_golden_model_1.P0INREG [3]);
  and _64641_ (_13002_, _08661_, \oc8051_golden_model_1.P1INREG [3]);
  nor _64642_ (_13003_, _13002_, _13001_);
  and _64643_ (_13004_, _13003_, _13000_);
  and _64644_ (_13005_, _13004_, _12997_);
  and _64645_ (_13006_, _13005_, _12994_);
  and _64646_ (_13007_, _13006_, _08357_);
  nor _64647_ (_13008_, _13007_, _12984_);
  and _64648_ (_13009_, _08633_, \oc8051_golden_model_1.TCON [5]);
  and _64649_ (_13010_, _08637_, \oc8051_golden_model_1.B [5]);
  nor _64650_ (_13011_, _13010_, _13009_);
  and _64651_ (_13012_, _08643_, \oc8051_golden_model_1.IP [5]);
  not _64652_ (_13013_, _13012_);
  and _64653_ (_13014_, _08640_, \oc8051_golden_model_1.PSW [5]);
  and _64654_ (_13015_, _08645_, \oc8051_golden_model_1.ACC [5]);
  nor _64655_ (_13016_, _13015_, _13014_);
  and _64656_ (_13017_, _13016_, _13013_);
  and _64657_ (_13018_, _13017_, _13011_);
  and _64658_ (_13019_, _08650_, \oc8051_golden_model_1.SCON [5]);
  and _64659_ (_13020_, _08652_, \oc8051_golden_model_1.IE [5]);
  nor _64660_ (_13021_, _13020_, _13019_);
  and _64661_ (_13022_, _08655_, \oc8051_golden_model_1.P2INREG [5]);
  and _64662_ (_13023_, _08657_, \oc8051_golden_model_1.P3INREG [5]);
  nor _64663_ (_13024_, _13023_, _13022_);
  and _64664_ (_13025_, _07993_, \oc8051_golden_model_1.P0INREG [5]);
  and _64665_ (_13026_, _08661_, \oc8051_golden_model_1.P1INREG [5]);
  nor _64666_ (_13027_, _13026_, _13025_);
  and _64667_ (_13028_, _13027_, _13024_);
  and _64668_ (_13029_, _13028_, _13021_);
  and _64669_ (_13030_, _13029_, _13018_);
  and _64670_ (_13031_, _13030_, _08306_);
  and _64671_ (_13032_, _07956_, _07799_);
  not _64672_ (_13033_, _13032_);
  nor _64673_ (_13034_, _13033_, _13031_);
  nor _64674_ (_13035_, _13034_, _13008_);
  and _64675_ (_13036_, _13035_, _12983_);
  and _64676_ (_13037_, _13036_, _12932_);
  not _64677_ (_13038_, _13037_);
  or _64678_ (_13039_, _12495_, _13038_);
  or _64679_ (_13040_, _09565_, _13037_);
  and _64680_ (_13041_, _13040_, _06512_);
  and _64681_ (_13042_, _13041_, _13039_);
  or _64682_ (_13043_, _13042_, _12854_);
  or _64683_ (_13044_, _13043_, _12853_);
  and _64684_ (_13045_, _13044_, _12202_);
  nor _64685_ (_13046_, _10566_, _06363_);
  not _64686_ (_13047_, _13046_);
  or _64687_ (_13048_, _13047_, _13045_);
  not _64688_ (_13049_, _10564_);
  or _64689_ (_13050_, _13046_, _09550_);
  and _64690_ (_13051_, _13050_, _13049_);
  and _64691_ (_13052_, _13051_, _13048_);
  and _64692_ (_13053_, _12200_, _10564_);
  or _64693_ (_13054_, _13053_, _06361_);
  or _64694_ (_13055_, _13054_, _13052_);
  nand _64695_ (_13056_, _08107_, _06361_);
  and _64696_ (_13057_, _13056_, _13055_);
  or _64697_ (_13058_, _13057_, _12187_);
  or _64698_ (_13059_, _09550_, _06021_);
  and _64699_ (_13060_, _13059_, _07035_);
  and _64700_ (_13061_, _13060_, _13058_);
  not _64701_ (_13062_, _09123_);
  or _64702_ (_13063_, _12495_, _13037_);
  nand _64703_ (_13064_, _12489_, _13037_);
  and _64704_ (_13065_, _13064_, _13063_);
  and _64705_ (_13066_, _13065_, _06496_);
  or _64706_ (_13067_, _13066_, _13062_);
  or _64707_ (_13068_, _13067_, _13061_);
  or _64708_ (_13069_, _12200_, _09123_);
  and _64709_ (_13070_, _13069_, _07048_);
  and _64710_ (_13071_, _13070_, _13068_);
  nor _64711_ (_13072_, _11382_, _11377_);
  nand _64712_ (_13073_, _09550_, _06639_);
  nand _64713_ (_13074_, _13073_, _13072_);
  or _64714_ (_13075_, _13074_, _13071_);
  or _64715_ (_13076_, _12200_, _13072_);
  and _64716_ (_13077_, _13076_, _09534_);
  and _64717_ (_13078_, _13077_, _13075_);
  and _64718_ (_13079_, _06503_, _06238_);
  or _64719_ (_13080_, _13079_, _05998_);
  or _64720_ (_13081_, _13080_, _13078_);
  not _64721_ (_13082_, _05998_);
  or _64722_ (_13083_, _09550_, _13082_);
  and _64723_ (_13084_, _13083_, _05990_);
  and _64724_ (_13085_, _13084_, _13081_);
  and _64725_ (_13086_, _13065_, _05989_);
  and _64726_ (_13087_, _09473_, _07375_);
  not _64727_ (_13088_, _13087_);
  or _64728_ (_13089_, _13088_, _13086_);
  or _64729_ (_13090_, _13089_, _13085_);
  or _64730_ (_13091_, _13087_, _12200_);
  and _64731_ (_13092_, _13091_, _06651_);
  and _64732_ (_13093_, _13092_, _13090_);
  nand _64733_ (_13094_, _09550_, _06646_);
  nor _64734_ (_13095_, _11407_, _11400_);
  nand _64735_ (_13096_, _13095_, _13094_);
  or _64736_ (_13097_, _13096_, _13093_);
  not _64737_ (_13098_, _06488_);
  or _64738_ (_13099_, _13095_, _12200_);
  and _64739_ (_13100_, _13099_, _13098_);
  and _64740_ (_13101_, _13100_, _13097_);
  and _64741_ (_13102_, _06488_, _06238_);
  or _64742_ (_13103_, _13102_, _05997_);
  or _64743_ (_13104_, _13103_, _13101_);
  and _64744_ (_13105_, _05996_, _05988_);
  not _64745_ (_13106_, _13105_);
  not _64746_ (_13107_, _05997_);
  or _64747_ (_13108_, _09550_, _13107_);
  and _64748_ (_13109_, _13108_, _13106_);
  and _64749_ (_13110_, _13109_, _13104_);
  and _64750_ (_13111_, _13105_, _12200_);
  or _64751_ (_13112_, _13111_, _13110_);
  or _64752_ (_13113_, _13112_, _01446_);
  or _64753_ (_13114_, _01442_, \oc8051_golden_model_1.PC [15]);
  and _64754_ (_13115_, _13114_, _43634_);
  and _64755_ (_41509_, _13115_, _13113_);
  nor _64756_ (_13116_, \oc8051_golden_model_1.P2 [7], rst);
  nor _64757_ (_13117_, _13116_, _00000_);
  not _64758_ (_13118_, \oc8051_golden_model_1.P2 [7]);
  nor _64759_ (_13119_, _08032_, _13118_);
  and _64760_ (_13120_, _08029_, \oc8051_golden_model_1.P1 [7]);
  not _64761_ (_13121_, _13120_);
  and _64762_ (_13122_, _08032_, \oc8051_golden_model_1.P2 [7]);
  and _64763_ (_13123_, _08034_, \oc8051_golden_model_1.P3 [7]);
  nor _64764_ (_13124_, _13123_, _13122_);
  and _64765_ (_13125_, _13124_, _13121_);
  and _64766_ (_13126_, _13125_, _08028_);
  and _64767_ (_13127_, _08039_, \oc8051_golden_model_1.P0 [7]);
  nor _64768_ (_13128_, _13127_, _08043_);
  and _64769_ (_13129_, _13128_, _13126_);
  and _64770_ (_13130_, _13129_, _08009_);
  and _64771_ (_13131_, _13130_, _07999_);
  and _64772_ (_13132_, _13131_, _08108_);
  nand _64773_ (_13133_, _13132_, _08688_);
  or _64774_ (_13134_, _13132_, _08688_);
  and _64775_ (_13135_, _13134_, _13133_);
  and _64776_ (_13136_, _13135_, _08032_);
  or _64777_ (_13137_, _13136_, _13119_);
  and _64778_ (_13138_, _13137_, _06615_);
  not _64779_ (_13139_, _08032_);
  nor _64780_ (_13140_, _08107_, _13139_);
  or _64781_ (_13141_, _13140_, _13119_);
  or _64782_ (_13142_, _13141_, _06327_);
  nor _64783_ (_13143_, _08655_, _13118_);
  and _64784_ (_13144_, _08661_, \oc8051_golden_model_1.P1 [7]);
  and _64785_ (_13145_, _08657_, \oc8051_golden_model_1.P3 [7]);
  nor _64786_ (_13146_, _13145_, _13144_);
  and _64787_ (_13147_, _07993_, \oc8051_golden_model_1.P0 [7]);
  and _64788_ (_13148_, _08655_, \oc8051_golden_model_1.P2 [7]);
  nor _64789_ (_13149_, _13148_, _13147_);
  and _64790_ (_13150_, _13149_, _13146_);
  and _64791_ (_13151_, _13150_, _08654_);
  and _64792_ (_13152_, _13151_, _08649_);
  and _64793_ (_13153_, _13152_, _08108_);
  nor _64794_ (_13154_, _13153_, _08041_);
  and _64795_ (_13155_, _13154_, _08655_);
  or _64796_ (_13156_, _13155_, _13143_);
  and _64797_ (_13157_, _13156_, _06352_);
  not _64798_ (_13158_, _13132_);
  not _64799_ (_13159_, _08120_);
  nor _64800_ (_13160_, _08121_, _08123_);
  and _64801_ (_13161_, _13160_, _08135_);
  and _64802_ (_13162_, _13161_, _13159_);
  and _64803_ (_13163_, _08032_, \oc8051_golden_model_1.P2 [6]);
  and _64804_ (_13164_, _08034_, \oc8051_golden_model_1.P3 [6]);
  nor _64805_ (_13165_, _13164_, _13163_);
  and _64806_ (_13166_, _08039_, \oc8051_golden_model_1.P0 [6]);
  and _64807_ (_13167_, _08029_, \oc8051_golden_model_1.P1 [6]);
  nor _64808_ (_13168_, _13167_, _13166_);
  and _64809_ (_13169_, _13168_, _13165_);
  and _64810_ (_13170_, _13169_, _08119_);
  and _64811_ (_13171_, _08129_, _08144_);
  and _64812_ (_13172_, _13171_, _13170_);
  and _64813_ (_13173_, _13172_, _08161_);
  and _64814_ (_13174_, _13173_, _13162_);
  and _64815_ (_13175_, _13174_, _08210_);
  and _64816_ (_13176_, _08032_, \oc8051_golden_model_1.P2 [5]);
  and _64817_ (_13177_, _08034_, \oc8051_golden_model_1.P3 [5]);
  nor _64818_ (_13178_, _13177_, _13176_);
  and _64819_ (_13179_, _08039_, \oc8051_golden_model_1.P0 [5]);
  and _64820_ (_13180_, _08029_, \oc8051_golden_model_1.P1 [5]);
  nor _64821_ (_13181_, _13180_, _13179_);
  and _64822_ (_13182_, _13181_, _13178_);
  and _64823_ (_13183_, _13182_, _08248_);
  and _64824_ (_13184_, _13183_, _08242_);
  and _64825_ (_13185_, _13184_, _08226_);
  and _64826_ (_13186_, _13185_, _08306_);
  and _64827_ (_13187_, _08032_, \oc8051_golden_model_1.P2 [4]);
  and _64828_ (_13188_, _08034_, \oc8051_golden_model_1.P3 [4]);
  nor _64829_ (_13189_, _13188_, _13187_);
  and _64830_ (_13190_, _08039_, \oc8051_golden_model_1.P0 [4]);
  and _64831_ (_13191_, _08029_, \oc8051_golden_model_1.P1 [4]);
  nor _64832_ (_13192_, _13191_, _13190_);
  and _64833_ (_13193_, _13192_, _13189_);
  and _64834_ (_13194_, _13193_, _08539_);
  and _64835_ (_13195_, _13194_, _08533_);
  and _64836_ (_13196_, _13195_, _08527_);
  and _64837_ (_13197_, _13196_, _08597_);
  and _64838_ (_13198_, _08032_, \oc8051_golden_model_1.P2 [3]);
  and _64839_ (_13199_, _08034_, \oc8051_golden_model_1.P3 [3]);
  nor _64840_ (_13200_, _13199_, _13198_);
  and _64841_ (_13201_, _08039_, \oc8051_golden_model_1.P0 [3]);
  and _64842_ (_13202_, _08029_, \oc8051_golden_model_1.P1 [3]);
  nor _64843_ (_13203_, _13202_, _13201_);
  and _64844_ (_13204_, _13203_, _13200_);
  and _64845_ (_13205_, _13204_, _08344_);
  and _64846_ (_13206_, _13205_, _08338_);
  and _64847_ (_13207_, _13206_, _08322_);
  and _64848_ (_13208_, _13207_, _08357_);
  and _64849_ (_13209_, _08032_, \oc8051_golden_model_1.P2 [2]);
  and _64850_ (_13210_, _08034_, \oc8051_golden_model_1.P3 [2]);
  nor _64851_ (_13211_, _13210_, _13209_);
  and _64852_ (_13212_, _08039_, \oc8051_golden_model_1.P0 [2]);
  and _64853_ (_13213_, _08029_, \oc8051_golden_model_1.P1 [2]);
  nor _64854_ (_13214_, _13213_, _13212_);
  and _64855_ (_13215_, _13214_, _13211_);
  and _64856_ (_13216_, _13215_, _08488_);
  and _64857_ (_13217_, _13216_, _08482_);
  and _64858_ (_13218_, _13217_, _08476_);
  and _64859_ (_13219_, _13218_, _08501_);
  and _64860_ (_13220_, _08032_, \oc8051_golden_model_1.P2 [1]);
  and _64861_ (_13221_, _08034_, \oc8051_golden_model_1.P3 [1]);
  nor _64862_ (_13222_, _13221_, _13220_);
  and _64863_ (_13223_, _08039_, \oc8051_golden_model_1.P0 [1]);
  and _64864_ (_13224_, _08029_, \oc8051_golden_model_1.P1 [1]);
  nor _64865_ (_13225_, _13224_, _13223_);
  and _64866_ (_13226_, _13225_, _13222_);
  and _64867_ (_13227_, _08390_, _08376_);
  not _64868_ (_13228_, _08368_);
  and _64869_ (_13229_, _08398_, _13228_);
  nor _64870_ (_13230_, _08384_, _08381_);
  nand _64871_ (_13231_, _13230_, _08393_);
  nor _64872_ (_13232_, _13231_, _08382_);
  and _64873_ (_13233_, _13232_, _13229_);
  and _64874_ (_13234_, _13233_, _13227_);
  and _64875_ (_13235_, _13234_, _13226_);
  and _64876_ (_13236_, _13235_, _08366_);
  and _64877_ (_13237_, _13236_, _08402_);
  and _64878_ (_13238_, _08032_, \oc8051_golden_model_1.P2 [0]);
  and _64879_ (_13239_, _08034_, \oc8051_golden_model_1.P3 [0]);
  nor _64880_ (_13240_, _13239_, _13238_);
  and _64881_ (_13241_, _08039_, \oc8051_golden_model_1.P0 [0]);
  and _64882_ (_13242_, _08029_, \oc8051_golden_model_1.P1 [0]);
  nor _64883_ (_13243_, _13242_, _13241_);
  and _64884_ (_13244_, _13243_, _13240_);
  and _64885_ (_13245_, _13244_, _08438_);
  and _64886_ (_13246_, _13245_, _08432_);
  and _64887_ (_13247_, _13246_, _08426_);
  and _64888_ (_13248_, _13247_, _08452_);
  and _64889_ (_13249_, _13248_, _13237_);
  and _64890_ (_13250_, _13249_, _13219_);
  and _64891_ (_13251_, _13250_, _13208_);
  and _64892_ (_13252_, _13251_, _13197_);
  and _64893_ (_13253_, _13252_, _13186_);
  and _64894_ (_13254_, _13253_, _13175_);
  or _64895_ (_13255_, _13254_, _13158_);
  nand _64896_ (_13256_, _13254_, _13158_);
  and _64897_ (_13257_, _13256_, _13255_);
  and _64898_ (_13258_, _13257_, _08032_);
  or _64899_ (_13259_, _13258_, _13119_);
  or _64900_ (_13260_, _13259_, _07275_);
  and _64901_ (_13261_, _08032_, \oc8051_golden_model_1.ACC [7]);
  or _64902_ (_13262_, _13261_, _13119_);
  and _64903_ (_13263_, _13262_, _07259_);
  nor _64904_ (_13264_, _07259_, _13118_);
  or _64905_ (_13265_, _13264_, _06474_);
  or _64906_ (_13266_, _13265_, _13263_);
  and _64907_ (_13267_, _13266_, _06357_);
  and _64908_ (_13268_, _13267_, _13260_);
  nand _64909_ (_13269_, _13153_, _08671_);
  and _64910_ (_13270_, _13269_, _08655_);
  or _64911_ (_13271_, _13270_, _13143_);
  and _64912_ (_13272_, _13271_, _06356_);
  or _64913_ (_13273_, _13272_, _06410_);
  or _64914_ (_13274_, _13273_, _13268_);
  or _64915_ (_13275_, _13141_, _06772_);
  and _64916_ (_13276_, _13275_, _13274_);
  or _64917_ (_13277_, _13276_, _06417_);
  or _64918_ (_13278_, _13262_, _06426_);
  and _64919_ (_13279_, _13278_, _06353_);
  and _64920_ (_13280_, _13279_, _13277_);
  or _64921_ (_13281_, _13280_, _13157_);
  and _64922_ (_13282_, _13281_, _06346_);
  or _64923_ (_13283_, _13153_, _08671_);
  or _64924_ (_13284_, _13283_, _13143_);
  and _64925_ (_13285_, _13271_, _06345_);
  and _64926_ (_13286_, _13285_, _13284_);
  or _64927_ (_13287_, _13286_, _13282_);
  and _64928_ (_13288_, _13287_, _06340_);
  or _64929_ (_13289_, _13154_, _08827_);
  and _64930_ (_13290_, _13289_, _08655_);
  or _64931_ (_13291_, _13290_, _13143_);
  and _64932_ (_13292_, _13291_, _06339_);
  or _64933_ (_13293_, _13292_, _10153_);
  or _64934_ (_13294_, _13293_, _13288_);
  and _64935_ (_13295_, _13294_, _13142_);
  or _64936_ (_13296_, _13295_, _09572_);
  and _64937_ (_13297_, _08778_, _08032_);
  or _64938_ (_13298_, _13119_, _06333_);
  or _64939_ (_13299_, _13298_, _13297_);
  and _64940_ (_13300_, _13299_, _06313_);
  and _64941_ (_13301_, _13300_, _13296_);
  and _64942_ (_13302_, _08993_, \oc8051_golden_model_1.P0 [7]);
  and _64943_ (_13303_, _08989_, \oc8051_golden_model_1.P2 [7]);
  and _64944_ (_13304_, _08998_, \oc8051_golden_model_1.P1 [7]);
  and _64945_ (_13305_, _09002_, \oc8051_golden_model_1.P3 [7]);
  or _64946_ (_13306_, _13305_, _13304_);
  or _64947_ (_13307_, _13306_, _13303_);
  or _64948_ (_13308_, _13307_, _13302_);
  or _64949_ (_13309_, _13308_, _09019_);
  or _64950_ (_13310_, _13309_, _09044_);
  or _64951_ (_13311_, _13310_, _09074_);
  or _64952_ (_13312_, _13311_, _08881_);
  and _64953_ (_13313_, _13312_, _08032_);
  or _64954_ (_13314_, _13313_, _13119_);
  and _64955_ (_13315_, _13314_, _06037_);
  or _64956_ (_13316_, _13315_, _06277_);
  or _64957_ (_13317_, _13316_, _13301_);
  and _64958_ (_13318_, _08880_, _08032_);
  or _64959_ (_13319_, _13318_, _13119_);
  or _64960_ (_13320_, _13319_, _06278_);
  and _64961_ (_13321_, _13320_, _13317_);
  or _64962_ (_13322_, _13321_, _06502_);
  nand _64963_ (_13323_, _13132_, _08879_);
  or _64964_ (_13324_, _13132_, _08879_);
  and _64965_ (_13325_, _13324_, _13323_);
  and _64966_ (_13326_, _13325_, _08032_);
  or _64967_ (_13327_, _13119_, _07334_);
  or _64968_ (_13328_, _13327_, _13326_);
  and _64969_ (_13329_, _13328_, _07337_);
  and _64970_ (_13330_, _13329_, _13322_);
  or _64971_ (_13331_, _13330_, _13138_);
  and _64972_ (_13332_, _13331_, _07339_);
  or _64973_ (_13333_, _13158_, _13119_);
  and _64974_ (_13334_, _13319_, _06507_);
  and _64975_ (_13335_, _13334_, _13333_);
  or _64976_ (_13336_, _13335_, _13332_);
  and _64977_ (_13337_, _13336_, _07331_);
  and _64978_ (_13338_, _13262_, _06610_);
  and _64979_ (_13339_, _13338_, _13333_);
  or _64980_ (_13340_, _13339_, _06509_);
  or _64981_ (_13341_, _13340_, _13337_);
  and _64982_ (_13342_, _13323_, _08032_);
  or _64983_ (_13343_, _13119_, _09107_);
  or _64984_ (_13344_, _13343_, _13342_);
  and _64985_ (_13345_, _13344_, _09112_);
  and _64986_ (_13346_, _13345_, _13341_);
  and _64987_ (_13347_, _13133_, _08032_);
  or _64988_ (_13348_, _13347_, _13119_);
  and _64989_ (_13349_, _13348_, _06602_);
  or _64990_ (_13350_, _13349_, _06639_);
  or _64991_ (_13351_, _13350_, _13346_);
  or _64992_ (_13352_, _13259_, _07048_);
  and _64993_ (_13353_, _13352_, _05990_);
  and _64994_ (_13354_, _13353_, _13351_);
  and _64995_ (_13355_, _13156_, _05989_);
  or _64996_ (_13356_, _13355_, _06646_);
  or _64997_ (_13357_, _13356_, _13354_);
  not _64998_ (_13358_, _13175_);
  not _64999_ (_13359_, _13186_);
  not _65000_ (_13360_, _13197_);
  not _65001_ (_13361_, _13208_);
  not _65002_ (_13362_, _13219_);
  nor _65003_ (_13363_, _13248_, _13237_);
  and _65004_ (_13364_, _13363_, _13362_);
  and _65005_ (_13365_, _13364_, _13361_);
  and _65006_ (_13366_, _13365_, _13360_);
  and _65007_ (_13367_, _13366_, _13359_);
  and _65008_ (_13368_, _13367_, _13358_);
  or _65009_ (_13369_, _13368_, _13158_);
  nand _65010_ (_13370_, _13368_, _13158_);
  and _65011_ (_13371_, _13370_, _13369_);
  and _65012_ (_13372_, _13371_, _08032_);
  or _65013_ (_13373_, _13119_, _06651_);
  or _65014_ (_13374_, _13373_, _13372_);
  and _65015_ (_13375_, _13374_, _01442_);
  and _65016_ (_13376_, _13375_, _13357_);
  or _65017_ (_41510_, _13376_, _13117_);
  nor _65018_ (_13377_, \oc8051_golden_model_1.P3 [7], rst);
  nor _65019_ (_13378_, _13377_, _00000_);
  not _65020_ (_13379_, _08034_);
  and _65021_ (_13380_, _13379_, \oc8051_golden_model_1.P3 [7]);
  and _65022_ (_13381_, _13135_, _08034_);
  or _65023_ (_13382_, _13381_, _13380_);
  and _65024_ (_13383_, _13382_, _06615_);
  nor _65025_ (_13384_, _08107_, _13379_);
  or _65026_ (_13385_, _13384_, _13380_);
  or _65027_ (_13386_, _13385_, _06327_);
  not _65028_ (_13387_, _08657_);
  and _65029_ (_13388_, _13387_, \oc8051_golden_model_1.P3 [7]);
  and _65030_ (_13389_, _13154_, _08657_);
  or _65031_ (_13390_, _13389_, _13388_);
  and _65032_ (_13391_, _13390_, _06352_);
  and _65033_ (_13392_, _13257_, _08034_);
  or _65034_ (_13393_, _13392_, _13380_);
  or _65035_ (_13394_, _13393_, _07275_);
  and _65036_ (_13395_, _08034_, \oc8051_golden_model_1.ACC [7]);
  or _65037_ (_13396_, _13395_, _13380_);
  and _65038_ (_13397_, _13396_, _07259_);
  and _65039_ (_13398_, _07260_, \oc8051_golden_model_1.P3 [7]);
  or _65040_ (_13399_, _13398_, _06474_);
  or _65041_ (_13400_, _13399_, _13397_);
  and _65042_ (_13401_, _13400_, _06357_);
  and _65043_ (_13402_, _13401_, _13394_);
  and _65044_ (_13403_, _13269_, _08657_);
  or _65045_ (_13404_, _13403_, _13388_);
  and _65046_ (_13405_, _13404_, _06356_);
  or _65047_ (_13406_, _13405_, _06410_);
  or _65048_ (_13407_, _13406_, _13402_);
  or _65049_ (_13408_, _13385_, _06772_);
  and _65050_ (_13409_, _13408_, _13407_);
  or _65051_ (_13410_, _13409_, _06417_);
  or _65052_ (_13411_, _13396_, _06426_);
  and _65053_ (_13412_, _13411_, _06353_);
  and _65054_ (_13413_, _13412_, _13410_);
  or _65055_ (_13414_, _13413_, _13391_);
  and _65056_ (_13415_, _13414_, _06346_);
  or _65057_ (_13416_, _13388_, _13283_);
  and _65058_ (_13417_, _13404_, _06345_);
  and _65059_ (_13418_, _13417_, _13416_);
  or _65060_ (_13419_, _13418_, _13415_);
  and _65061_ (_13420_, _13419_, _06340_);
  and _65062_ (_13421_, _13289_, _08657_);
  or _65063_ (_13422_, _13421_, _13388_);
  and _65064_ (_13423_, _13422_, _06339_);
  or _65065_ (_13424_, _13423_, _10153_);
  or _65066_ (_13425_, _13424_, _13420_);
  and _65067_ (_13426_, _13425_, _13386_);
  or _65068_ (_13427_, _13426_, _09572_);
  and _65069_ (_13428_, _08778_, _08034_);
  or _65070_ (_13429_, _13380_, _06333_);
  or _65071_ (_13430_, _13429_, _13428_);
  and _65072_ (_13431_, _13430_, _06313_);
  and _65073_ (_13432_, _13431_, _13427_);
  and _65074_ (_13433_, _13312_, _08034_);
  or _65075_ (_13434_, _13433_, _13380_);
  and _65076_ (_13435_, _13434_, _06037_);
  or _65077_ (_13436_, _13435_, _06277_);
  or _65078_ (_13437_, _13436_, _13432_);
  and _65079_ (_13438_, _08880_, _08034_);
  or _65080_ (_13439_, _13438_, _13380_);
  or _65081_ (_13440_, _13439_, _06278_);
  and _65082_ (_13441_, _13440_, _13437_);
  or _65083_ (_13442_, _13441_, _06502_);
  and _65084_ (_13443_, _13325_, _08034_);
  or _65085_ (_13444_, _13380_, _07334_);
  or _65086_ (_13445_, _13444_, _13443_);
  and _65087_ (_13446_, _13445_, _07337_);
  and _65088_ (_13447_, _13446_, _13442_);
  or _65089_ (_13448_, _13447_, _13383_);
  and _65090_ (_13449_, _13448_, _07339_);
  or _65091_ (_13450_, _13380_, _13158_);
  and _65092_ (_13451_, _13439_, _06507_);
  and _65093_ (_13452_, _13451_, _13450_);
  or _65094_ (_13453_, _13452_, _13449_);
  and _65095_ (_13454_, _13453_, _07331_);
  and _65096_ (_13455_, _13396_, _06610_);
  and _65097_ (_13456_, _13455_, _13450_);
  or _65098_ (_13457_, _13456_, _06509_);
  or _65099_ (_13458_, _13457_, _13454_);
  and _65100_ (_13459_, _13323_, _08034_);
  or _65101_ (_13460_, _13380_, _09107_);
  or _65102_ (_13461_, _13460_, _13459_);
  and _65103_ (_13462_, _13461_, _09112_);
  and _65104_ (_13463_, _13462_, _13458_);
  and _65105_ (_13464_, _13133_, _08034_);
  or _65106_ (_13465_, _13464_, _13380_);
  and _65107_ (_13466_, _13465_, _06602_);
  or _65108_ (_13467_, _13466_, _06639_);
  or _65109_ (_13468_, _13467_, _13463_);
  or _65110_ (_13469_, _13393_, _07048_);
  and _65111_ (_13470_, _13469_, _05990_);
  and _65112_ (_13471_, _13470_, _13468_);
  and _65113_ (_13472_, _13390_, _05989_);
  or _65114_ (_13473_, _13472_, _06646_);
  or _65115_ (_13474_, _13473_, _13471_);
  and _65116_ (_13475_, _13371_, _08034_);
  or _65117_ (_13476_, _13380_, _06651_);
  or _65118_ (_13477_, _13476_, _13475_);
  and _65119_ (_13478_, _13477_, _01442_);
  and _65120_ (_13479_, _13478_, _13474_);
  or _65121_ (_41511_, _13479_, _13378_);
  nor _65122_ (_13480_, \oc8051_golden_model_1.P0 [7], rst);
  nor _65123_ (_13481_, _13480_, _00000_);
  not _65124_ (_13482_, _08039_);
  and _65125_ (_13483_, _13482_, \oc8051_golden_model_1.P0 [7]);
  and _65126_ (_13484_, _13135_, _08039_);
  or _65127_ (_13485_, _13484_, _13483_);
  and _65128_ (_13486_, _13485_, _06615_);
  nor _65129_ (_13487_, _08107_, _13482_);
  or _65130_ (_13488_, _13487_, _13483_);
  or _65131_ (_13489_, _13488_, _06327_);
  not _65132_ (_13490_, _07993_);
  and _65133_ (_13491_, _13490_, \oc8051_golden_model_1.P0 [7]);
  and _65134_ (_13492_, _13154_, _07993_);
  or _65135_ (_13493_, _13492_, _13491_);
  and _65136_ (_13494_, _13493_, _06352_);
  and _65137_ (_13495_, _13257_, _08039_);
  or _65138_ (_13496_, _13495_, _13483_);
  or _65139_ (_13497_, _13496_, _07275_);
  and _65140_ (_13498_, _08039_, \oc8051_golden_model_1.ACC [7]);
  or _65141_ (_13499_, _13498_, _13483_);
  and _65142_ (_13500_, _13499_, _07259_);
  and _65143_ (_13501_, _07260_, \oc8051_golden_model_1.P0 [7]);
  or _65144_ (_13502_, _13501_, _06474_);
  or _65145_ (_13503_, _13502_, _13500_);
  and _65146_ (_13504_, _13503_, _06357_);
  and _65147_ (_13505_, _13504_, _13497_);
  and _65148_ (_13506_, _13269_, _07993_);
  or _65149_ (_13507_, _13506_, _13491_);
  and _65150_ (_13508_, _13507_, _06356_);
  or _65151_ (_13509_, _13508_, _06410_);
  or _65152_ (_13510_, _13509_, _13505_);
  or _65153_ (_13511_, _13488_, _06772_);
  and _65154_ (_13512_, _13511_, _13510_);
  or _65155_ (_13513_, _13512_, _06417_);
  or _65156_ (_13514_, _13499_, _06426_);
  and _65157_ (_13515_, _13514_, _06353_);
  and _65158_ (_13516_, _13515_, _13513_);
  or _65159_ (_13517_, _13516_, _13494_);
  and _65160_ (_13518_, _13517_, _06346_);
  or _65161_ (_13519_, _13491_, _13283_);
  and _65162_ (_13520_, _13507_, _06345_);
  and _65163_ (_13521_, _13520_, _13519_);
  or _65164_ (_13522_, _13521_, _13518_);
  and _65165_ (_13523_, _13522_, _06340_);
  and _65166_ (_13524_, _13289_, _07993_);
  or _65167_ (_13525_, _13524_, _13491_);
  and _65168_ (_13526_, _13525_, _06339_);
  or _65169_ (_13527_, _13526_, _10153_);
  or _65170_ (_13528_, _13527_, _13523_);
  and _65171_ (_13529_, _13528_, _13489_);
  or _65172_ (_13530_, _13529_, _09572_);
  and _65173_ (_13531_, _08778_, _08039_);
  or _65174_ (_13532_, _13483_, _06333_);
  or _65175_ (_13533_, _13532_, _13531_);
  and _65176_ (_13534_, _13533_, _06313_);
  and _65177_ (_13535_, _13534_, _13530_);
  and _65178_ (_13536_, _13312_, _08039_);
  or _65179_ (_13537_, _13536_, _13483_);
  and _65180_ (_13538_, _13537_, _06037_);
  or _65181_ (_13539_, _13538_, _06277_);
  or _65182_ (_13540_, _13539_, _13535_);
  and _65183_ (_13541_, _08880_, _08039_);
  or _65184_ (_13542_, _13541_, _13483_);
  or _65185_ (_13543_, _13542_, _06278_);
  and _65186_ (_13544_, _13543_, _13540_);
  or _65187_ (_13545_, _13544_, _06502_);
  and _65188_ (_13546_, _13325_, _08039_);
  or _65189_ (_13547_, _13483_, _07334_);
  or _65190_ (_13548_, _13547_, _13546_);
  and _65191_ (_13549_, _13548_, _07337_);
  and _65192_ (_13550_, _13549_, _13545_);
  or _65193_ (_13551_, _13550_, _13486_);
  and _65194_ (_13552_, _13551_, _07339_);
  or _65195_ (_13553_, _13483_, _13158_);
  and _65196_ (_13554_, _13542_, _06507_);
  and _65197_ (_13555_, _13554_, _13553_);
  or _65198_ (_13556_, _13555_, _13552_);
  and _65199_ (_13557_, _13556_, _07331_);
  and _65200_ (_13558_, _13499_, _06610_);
  and _65201_ (_13559_, _13558_, _13553_);
  or _65202_ (_13560_, _13559_, _06509_);
  or _65203_ (_13561_, _13560_, _13557_);
  and _65204_ (_13562_, _13323_, _08039_);
  or _65205_ (_13563_, _13483_, _09107_);
  or _65206_ (_13564_, _13563_, _13562_);
  and _65207_ (_13565_, _13564_, _09112_);
  and _65208_ (_13566_, _13565_, _13561_);
  and _65209_ (_13567_, _13133_, _08039_);
  or _65210_ (_13568_, _13567_, _13483_);
  and _65211_ (_13569_, _13568_, _06602_);
  or _65212_ (_13570_, _13569_, _06639_);
  or _65213_ (_13571_, _13570_, _13566_);
  or _65214_ (_13572_, _13496_, _07048_);
  and _65215_ (_13573_, _13572_, _05990_);
  and _65216_ (_13574_, _13573_, _13571_);
  and _65217_ (_13575_, _13493_, _05989_);
  or _65218_ (_13576_, _13575_, _06646_);
  or _65219_ (_13577_, _13576_, _13574_);
  and _65220_ (_13578_, _13371_, _08039_);
  or _65221_ (_13579_, _13483_, _06651_);
  or _65222_ (_13580_, _13579_, _13578_);
  and _65223_ (_13581_, _13580_, _01442_);
  and _65224_ (_13582_, _13581_, _13577_);
  or _65225_ (_41513_, _13582_, _13481_);
  nor _65226_ (_13583_, \oc8051_golden_model_1.P1 [7], rst);
  nor _65227_ (_13584_, _13583_, _00000_);
  not _65228_ (_13585_, _08029_);
  and _65229_ (_13586_, _13585_, \oc8051_golden_model_1.P1 [7]);
  and _65230_ (_13587_, _13135_, _08029_);
  or _65231_ (_13588_, _13587_, _13586_);
  and _65232_ (_13589_, _13588_, _06615_);
  nor _65233_ (_13590_, _08107_, _13585_);
  or _65234_ (_13591_, _13590_, _13586_);
  or _65235_ (_13592_, _13591_, _06327_);
  not _65236_ (_13593_, _08661_);
  and _65237_ (_13594_, _13593_, \oc8051_golden_model_1.P1 [7]);
  and _65238_ (_13595_, _13154_, _08661_);
  or _65239_ (_13596_, _13595_, _13594_);
  and _65240_ (_13597_, _13596_, _06352_);
  and _65241_ (_13598_, _13257_, _08029_);
  or _65242_ (_13599_, _13598_, _13586_);
  or _65243_ (_13600_, _13599_, _07275_);
  and _65244_ (_13601_, _08029_, \oc8051_golden_model_1.ACC [7]);
  or _65245_ (_13602_, _13601_, _13586_);
  and _65246_ (_13603_, _13602_, _07259_);
  and _65247_ (_13604_, _07260_, \oc8051_golden_model_1.P1 [7]);
  or _65248_ (_13605_, _13604_, _06474_);
  or _65249_ (_13606_, _13605_, _13603_);
  and _65250_ (_13607_, _13606_, _06357_);
  and _65251_ (_13608_, _13607_, _13600_);
  and _65252_ (_13609_, _13269_, _08661_);
  or _65253_ (_13610_, _13609_, _13594_);
  and _65254_ (_13611_, _13610_, _06356_);
  or _65255_ (_13612_, _13611_, _06410_);
  or _65256_ (_13613_, _13612_, _13608_);
  or _65257_ (_13614_, _13591_, _06772_);
  and _65258_ (_13615_, _13614_, _13613_);
  or _65259_ (_13616_, _13615_, _06417_);
  or _65260_ (_13617_, _13602_, _06426_);
  and _65261_ (_13618_, _13617_, _06353_);
  and _65262_ (_13619_, _13618_, _13616_);
  or _65263_ (_13620_, _13619_, _13597_);
  and _65264_ (_13621_, _13620_, _06346_);
  or _65265_ (_13622_, _13594_, _13283_);
  and _65266_ (_13623_, _13610_, _06345_);
  and _65267_ (_13624_, _13623_, _13622_);
  or _65268_ (_13625_, _13624_, _13621_);
  and _65269_ (_13626_, _13625_, _06340_);
  and _65270_ (_13627_, _13289_, _08661_);
  or _65271_ (_13628_, _13627_, _13594_);
  and _65272_ (_13629_, _13628_, _06339_);
  or _65273_ (_13630_, _13629_, _10153_);
  or _65274_ (_13631_, _13630_, _13626_);
  and _65275_ (_13632_, _13631_, _13592_);
  or _65276_ (_13633_, _13632_, _09572_);
  and _65277_ (_13634_, _08778_, _08029_);
  or _65278_ (_13635_, _13586_, _06333_);
  or _65279_ (_13636_, _13635_, _13634_);
  and _65280_ (_13638_, _13636_, _06313_);
  and _65281_ (_13639_, _13638_, _13633_);
  and _65282_ (_13640_, _13312_, _08029_);
  or _65283_ (_13641_, _13640_, _13586_);
  and _65284_ (_13642_, _13641_, _06037_);
  or _65285_ (_13643_, _13642_, _06277_);
  or _65286_ (_13644_, _13643_, _13639_);
  and _65287_ (_13645_, _08880_, _08029_);
  or _65288_ (_13646_, _13645_, _13586_);
  or _65289_ (_13647_, _13646_, _06278_);
  and _65290_ (_13649_, _13647_, _13644_);
  or _65291_ (_13650_, _13649_, _06502_);
  and _65292_ (_13651_, _13325_, _08029_);
  or _65293_ (_13652_, _13586_, _07334_);
  or _65294_ (_13653_, _13652_, _13651_);
  and _65295_ (_13654_, _13653_, _07337_);
  and _65296_ (_13655_, _13654_, _13650_);
  or _65297_ (_13656_, _13655_, _13589_);
  and _65298_ (_13657_, _13656_, _07339_);
  or _65299_ (_13658_, _13586_, _13158_);
  and _65300_ (_13660_, _13646_, _06507_);
  and _65301_ (_13661_, _13660_, _13658_);
  or _65302_ (_13662_, _13661_, _13657_);
  and _65303_ (_13663_, _13662_, _07331_);
  and _65304_ (_13664_, _13602_, _06610_);
  and _65305_ (_13665_, _13664_, _13658_);
  or _65306_ (_13666_, _13665_, _06509_);
  or _65307_ (_13667_, _13666_, _13663_);
  and _65308_ (_13668_, _13323_, _08029_);
  or _65309_ (_13669_, _13586_, _09107_);
  or _65310_ (_13671_, _13669_, _13668_);
  and _65311_ (_13672_, _13671_, _09112_);
  and _65312_ (_13673_, _13672_, _13667_);
  and _65313_ (_13674_, _13133_, _08029_);
  or _65314_ (_13675_, _13674_, _13586_);
  and _65315_ (_13676_, _13675_, _06602_);
  or _65316_ (_13677_, _13676_, _06639_);
  or _65317_ (_13678_, _13677_, _13673_);
  or _65318_ (_13679_, _13599_, _07048_);
  and _65319_ (_13680_, _13679_, _05990_);
  and _65320_ (_13682_, _13680_, _13678_);
  and _65321_ (_13683_, _13596_, _05989_);
  or _65322_ (_13684_, _13683_, _06646_);
  or _65323_ (_13685_, _13684_, _13682_);
  and _65324_ (_13686_, _13371_, _08029_);
  or _65325_ (_13687_, _13586_, _06651_);
  or _65326_ (_13688_, _13687_, _13686_);
  and _65327_ (_13689_, _13688_, _01442_);
  and _65328_ (_13690_, _13689_, _13685_);
  or _65329_ (_41514_, _13690_, _13584_);
  and _65330_ (_13692_, _01446_, \oc8051_golden_model_1.IP [7]);
  not _65331_ (_13693_, _08022_);
  and _65332_ (_13694_, _13693_, \oc8051_golden_model_1.IP [7]);
  and _65333_ (_13695_, _09096_, _08022_);
  or _65334_ (_13696_, _13695_, _13694_);
  and _65335_ (_13697_, _13696_, _06615_);
  nor _65336_ (_13698_, _08107_, _13693_);
  or _65337_ (_13699_, _13698_, _13694_);
  or _65338_ (_13700_, _13699_, _06327_);
  not _65339_ (_13701_, _08643_);
  and _65340_ (_13703_, _13701_, \oc8051_golden_model_1.IP [7]);
  and _65341_ (_13704_, _08668_, _08643_);
  or _65342_ (_13705_, _13704_, _13703_);
  and _65343_ (_13706_, _13705_, _06352_);
  and _65344_ (_13707_, _08791_, _08022_);
  or _65345_ (_13708_, _13707_, _13694_);
  or _65346_ (_13709_, _13708_, _07275_);
  and _65347_ (_13710_, _08022_, \oc8051_golden_model_1.ACC [7]);
  or _65348_ (_13711_, _13710_, _13694_);
  and _65349_ (_13712_, _13711_, _07259_);
  and _65350_ (_13714_, _07260_, \oc8051_golden_model_1.IP [7]);
  or _65351_ (_13715_, _13714_, _06474_);
  or _65352_ (_13716_, _13715_, _13712_);
  and _65353_ (_13717_, _13716_, _06357_);
  and _65354_ (_13718_, _13717_, _13709_);
  and _65355_ (_13719_, _08672_, _08643_);
  or _65356_ (_13720_, _13719_, _13703_);
  and _65357_ (_13721_, _13720_, _06356_);
  or _65358_ (_13722_, _13721_, _06410_);
  or _65359_ (_13723_, _13722_, _13718_);
  or _65360_ (_13725_, _13699_, _06772_);
  and _65361_ (_13726_, _13725_, _13723_);
  or _65362_ (_13727_, _13726_, _06417_);
  or _65363_ (_13728_, _13711_, _06426_);
  and _65364_ (_13729_, _13728_, _06353_);
  and _65365_ (_13730_, _13729_, _13727_);
  or _65366_ (_13731_, _13730_, _13706_);
  and _65367_ (_13732_, _13731_, _06346_);
  and _65368_ (_13733_, _08810_, _08643_);
  or _65369_ (_13734_, _13733_, _13703_);
  and _65370_ (_13736_, _13734_, _06345_);
  or _65371_ (_13737_, _13736_, _13732_);
  and _65372_ (_13738_, _13737_, _06340_);
  and _65373_ (_13739_, _08828_, _08643_);
  or _65374_ (_13740_, _13739_, _13703_);
  and _65375_ (_13741_, _13740_, _06339_);
  or _65376_ (_13742_, _13741_, _10153_);
  or _65377_ (_13743_, _13742_, _13738_);
  and _65378_ (_13744_, _13743_, _13700_);
  or _65379_ (_13745_, _13744_, _09572_);
  and _65380_ (_13747_, _08778_, _08022_);
  or _65381_ (_13748_, _13694_, _06333_);
  or _65382_ (_13749_, _13748_, _13747_);
  and _65383_ (_13750_, _13749_, _06313_);
  and _65384_ (_13751_, _13750_, _13745_);
  and _65385_ (_13752_, _09076_, _08022_);
  or _65386_ (_13753_, _13752_, _13694_);
  and _65387_ (_13754_, _13753_, _06037_);
  or _65388_ (_13755_, _13754_, _06277_);
  or _65389_ (_13756_, _13755_, _13751_);
  and _65390_ (_13758_, _08880_, _08022_);
  or _65391_ (_13759_, _13758_, _13694_);
  or _65392_ (_13760_, _13759_, _06278_);
  and _65393_ (_13761_, _13760_, _13756_);
  or _65394_ (_13762_, _13761_, _06502_);
  and _65395_ (_13763_, _09090_, _08022_);
  or _65396_ (_13764_, _13694_, _07334_);
  or _65397_ (_13765_, _13764_, _13763_);
  and _65398_ (_13766_, _13765_, _07337_);
  and _65399_ (_13767_, _13766_, _13762_);
  or _65400_ (_13769_, _13767_, _13697_);
  and _65401_ (_13770_, _13769_, _07339_);
  or _65402_ (_13771_, _13694_, _08110_);
  and _65403_ (_13772_, _13759_, _06507_);
  and _65404_ (_13773_, _13772_, _13771_);
  or _65405_ (_13774_, _13773_, _13770_);
  and _65406_ (_13775_, _13774_, _07331_);
  and _65407_ (_13776_, _13711_, _06610_);
  and _65408_ (_13777_, _13776_, _13771_);
  or _65409_ (_13778_, _13777_, _06509_);
  or _65410_ (_13780_, _13778_, _13775_);
  and _65411_ (_13781_, _09087_, _08022_);
  or _65412_ (_13782_, _13694_, _09107_);
  or _65413_ (_13783_, _13782_, _13781_);
  and _65414_ (_13784_, _13783_, _09112_);
  and _65415_ (_13785_, _13784_, _13780_);
  nor _65416_ (_13786_, _09095_, _13693_);
  or _65417_ (_13787_, _13786_, _13694_);
  and _65418_ (_13788_, _13787_, _06602_);
  or _65419_ (_13789_, _13788_, _06639_);
  or _65420_ (_13790_, _13789_, _13785_);
  or _65421_ (_13791_, _13708_, _07048_);
  and _65422_ (_13792_, _13791_, _05990_);
  and _65423_ (_13793_, _13792_, _13790_);
  and _65424_ (_13794_, _13705_, _05989_);
  or _65425_ (_13795_, _13794_, _06646_);
  or _65426_ (_13796_, _13795_, _13793_);
  and _65427_ (_13797_, _08605_, _08022_);
  or _65428_ (_13798_, _13694_, _06651_);
  or _65429_ (_13799_, _13798_, _13797_);
  and _65430_ (_13800_, _13799_, _01442_);
  and _65431_ (_13801_, _13800_, _13796_);
  or _65432_ (_13802_, _13801_, _13692_);
  and _65433_ (_41515_, _13802_, _43634_);
  and _65434_ (_13803_, _01446_, \oc8051_golden_model_1.IE [7]);
  not _65435_ (_13804_, _07986_);
  and _65436_ (_13805_, _13804_, \oc8051_golden_model_1.IE [7]);
  and _65437_ (_13806_, _09096_, _07986_);
  or _65438_ (_13807_, _13806_, _13805_);
  and _65439_ (_13808_, _13807_, _06615_);
  nor _65440_ (_13809_, _08107_, _13804_);
  or _65441_ (_13810_, _13809_, _13805_);
  or _65442_ (_13811_, _13810_, _06327_);
  not _65443_ (_13812_, _08652_);
  and _65444_ (_13813_, _13812_, \oc8051_golden_model_1.IE [7]);
  and _65445_ (_13814_, _08668_, _08652_);
  or _65446_ (_13815_, _13814_, _13813_);
  and _65447_ (_13816_, _13815_, _06352_);
  and _65448_ (_13817_, _08791_, _07986_);
  or _65449_ (_13818_, _13817_, _13805_);
  or _65450_ (_13819_, _13818_, _07275_);
  and _65451_ (_13820_, _07986_, \oc8051_golden_model_1.ACC [7]);
  or _65452_ (_13821_, _13820_, _13805_);
  and _65453_ (_13822_, _13821_, _07259_);
  and _65454_ (_13823_, _07260_, \oc8051_golden_model_1.IE [7]);
  or _65455_ (_13824_, _13823_, _06474_);
  or _65456_ (_13825_, _13824_, _13822_);
  and _65457_ (_13826_, _13825_, _06357_);
  and _65458_ (_13827_, _13826_, _13819_);
  and _65459_ (_13828_, _08672_, _08652_);
  or _65460_ (_13829_, _13828_, _13813_);
  and _65461_ (_13830_, _13829_, _06356_);
  or _65462_ (_13831_, _13830_, _06410_);
  or _65463_ (_13832_, _13831_, _13827_);
  or _65464_ (_13833_, _13810_, _06772_);
  and _65465_ (_13834_, _13833_, _13832_);
  or _65466_ (_13835_, _13834_, _06417_);
  or _65467_ (_13836_, _13821_, _06426_);
  and _65468_ (_13837_, _13836_, _06353_);
  and _65469_ (_13838_, _13837_, _13835_);
  or _65470_ (_13839_, _13838_, _13816_);
  and _65471_ (_13840_, _13839_, _06346_);
  and _65472_ (_13841_, _08810_, _08652_);
  or _65473_ (_13842_, _13841_, _13813_);
  and _65474_ (_13843_, _13842_, _06345_);
  or _65475_ (_13844_, _13843_, _13840_);
  and _65476_ (_13845_, _13844_, _06340_);
  and _65477_ (_13846_, _08828_, _08652_);
  or _65478_ (_13847_, _13846_, _13813_);
  and _65479_ (_13848_, _13847_, _06339_);
  or _65480_ (_13849_, _13848_, _10153_);
  or _65481_ (_13850_, _13849_, _13845_);
  and _65482_ (_13851_, _13850_, _13811_);
  or _65483_ (_13852_, _13851_, _09572_);
  and _65484_ (_13853_, _08778_, _07986_);
  or _65485_ (_13854_, _13805_, _06333_);
  or _65486_ (_13855_, _13854_, _13853_);
  and _65487_ (_13856_, _13855_, _06313_);
  and _65488_ (_13857_, _13856_, _13852_);
  and _65489_ (_13858_, _09076_, _07986_);
  or _65490_ (_13859_, _13858_, _13805_);
  and _65491_ (_13860_, _13859_, _06037_);
  or _65492_ (_13861_, _13860_, _06277_);
  or _65493_ (_13862_, _13861_, _13857_);
  and _65494_ (_13863_, _08880_, _07986_);
  or _65495_ (_13864_, _13863_, _13805_);
  or _65496_ (_13865_, _13864_, _06278_);
  and _65497_ (_13866_, _13865_, _13862_);
  or _65498_ (_13867_, _13866_, _06502_);
  and _65499_ (_13868_, _09090_, _07986_);
  or _65500_ (_13869_, _13805_, _07334_);
  or _65501_ (_13870_, _13869_, _13868_);
  and _65502_ (_13871_, _13870_, _07337_);
  and _65503_ (_13872_, _13871_, _13867_);
  or _65504_ (_13873_, _13872_, _13808_);
  and _65505_ (_13874_, _13873_, _07339_);
  or _65506_ (_13875_, _13805_, _08110_);
  and _65507_ (_13876_, _13864_, _06507_);
  and _65508_ (_13877_, _13876_, _13875_);
  or _65509_ (_13878_, _13877_, _13874_);
  and _65510_ (_13879_, _13878_, _07331_);
  and _65511_ (_13880_, _13821_, _06610_);
  and _65512_ (_13881_, _13880_, _13875_);
  or _65513_ (_13882_, _13881_, _06509_);
  or _65514_ (_13883_, _13882_, _13879_);
  and _65515_ (_13884_, _09087_, _07986_);
  or _65516_ (_13885_, _13805_, _09107_);
  or _65517_ (_13886_, _13885_, _13884_);
  and _65518_ (_13887_, _13886_, _09112_);
  and _65519_ (_13888_, _13887_, _13883_);
  nor _65520_ (_13889_, _09095_, _13804_);
  or _65521_ (_13890_, _13889_, _13805_);
  and _65522_ (_13891_, _13890_, _06602_);
  or _65523_ (_13892_, _13891_, _06639_);
  or _65524_ (_13893_, _13892_, _13888_);
  or _65525_ (_13894_, _13818_, _07048_);
  and _65526_ (_13895_, _13894_, _05990_);
  and _65527_ (_13896_, _13895_, _13893_);
  and _65528_ (_13897_, _13815_, _05989_);
  or _65529_ (_13898_, _13897_, _06646_);
  or _65530_ (_13899_, _13898_, _13896_);
  and _65531_ (_13900_, _08605_, _07986_);
  or _65532_ (_13901_, _13805_, _06651_);
  or _65533_ (_13902_, _13901_, _13900_);
  and _65534_ (_13903_, _13902_, _01442_);
  and _65535_ (_13904_, _13903_, _13899_);
  or _65536_ (_13905_, _13904_, _13803_);
  and _65537_ (_41516_, _13905_, _43634_);
  and _65538_ (_13906_, _01446_, \oc8051_golden_model_1.SCON [7]);
  not _65539_ (_13907_, _07969_);
  and _65540_ (_13908_, _13907_, \oc8051_golden_model_1.SCON [7]);
  and _65541_ (_13909_, _09096_, _07969_);
  or _65542_ (_13910_, _13909_, _13908_);
  and _65543_ (_13911_, _13910_, _06615_);
  nor _65544_ (_13912_, _08107_, _13907_);
  or _65545_ (_13913_, _13912_, _13908_);
  or _65546_ (_13914_, _13913_, _06327_);
  not _65547_ (_13915_, _08650_);
  and _65548_ (_13916_, _13915_, \oc8051_golden_model_1.SCON [7]);
  and _65549_ (_13917_, _08668_, _08650_);
  or _65550_ (_13918_, _13917_, _13916_);
  and _65551_ (_13919_, _13918_, _06352_);
  and _65552_ (_13920_, _08791_, _07969_);
  or _65553_ (_13921_, _13920_, _13908_);
  or _65554_ (_13922_, _13921_, _07275_);
  and _65555_ (_13923_, _07969_, \oc8051_golden_model_1.ACC [7]);
  or _65556_ (_13924_, _13923_, _13908_);
  and _65557_ (_13925_, _13924_, _07259_);
  and _65558_ (_13926_, _07260_, \oc8051_golden_model_1.SCON [7]);
  or _65559_ (_13927_, _13926_, _06474_);
  or _65560_ (_13928_, _13927_, _13925_);
  and _65561_ (_13929_, _13928_, _06357_);
  and _65562_ (_13930_, _13929_, _13922_);
  and _65563_ (_13931_, _08672_, _08650_);
  or _65564_ (_13932_, _13931_, _13916_);
  and _65565_ (_13933_, _13932_, _06356_);
  or _65566_ (_13934_, _13933_, _06410_);
  or _65567_ (_13935_, _13934_, _13930_);
  or _65568_ (_13936_, _13913_, _06772_);
  and _65569_ (_13937_, _13936_, _13935_);
  or _65570_ (_13938_, _13937_, _06417_);
  or _65571_ (_13939_, _13924_, _06426_);
  and _65572_ (_13940_, _13939_, _06353_);
  and _65573_ (_13941_, _13940_, _13938_);
  or _65574_ (_13942_, _13941_, _13919_);
  and _65575_ (_13943_, _13942_, _06346_);
  and _65576_ (_13944_, _08810_, _08650_);
  or _65577_ (_13945_, _13944_, _13916_);
  and _65578_ (_13946_, _13945_, _06345_);
  or _65579_ (_13947_, _13946_, _13943_);
  and _65580_ (_13948_, _13947_, _06340_);
  and _65581_ (_13949_, _08828_, _08650_);
  or _65582_ (_13950_, _13949_, _13916_);
  and _65583_ (_13951_, _13950_, _06339_);
  or _65584_ (_13952_, _13951_, _10153_);
  or _65585_ (_13953_, _13952_, _13948_);
  and _65586_ (_13954_, _13953_, _13914_);
  or _65587_ (_13955_, _13954_, _09572_);
  and _65588_ (_13956_, _08778_, _07969_);
  or _65589_ (_13957_, _13908_, _06333_);
  or _65590_ (_13958_, _13957_, _13956_);
  and _65591_ (_13959_, _13958_, _06313_);
  and _65592_ (_13960_, _13959_, _13955_);
  and _65593_ (_13961_, _09076_, _07969_);
  or _65594_ (_13962_, _13961_, _13908_);
  and _65595_ (_13963_, _13962_, _06037_);
  or _65596_ (_13964_, _13963_, _06277_);
  or _65597_ (_13965_, _13964_, _13960_);
  and _65598_ (_13966_, _08880_, _07969_);
  or _65599_ (_13967_, _13966_, _13908_);
  or _65600_ (_13968_, _13967_, _06278_);
  and _65601_ (_13969_, _13968_, _13965_);
  or _65602_ (_13970_, _13969_, _06502_);
  and _65603_ (_13971_, _09090_, _07969_);
  or _65604_ (_13972_, _13908_, _07334_);
  or _65605_ (_13973_, _13972_, _13971_);
  and _65606_ (_13974_, _13973_, _07337_);
  and _65607_ (_13975_, _13974_, _13970_);
  or _65608_ (_13976_, _13975_, _13911_);
  and _65609_ (_13977_, _13976_, _07339_);
  or _65610_ (_13978_, _13908_, _08110_);
  and _65611_ (_13979_, _13967_, _06507_);
  and _65612_ (_13980_, _13979_, _13978_);
  or _65613_ (_13981_, _13980_, _13977_);
  and _65614_ (_13982_, _13981_, _07331_);
  and _65615_ (_13983_, _13924_, _06610_);
  and _65616_ (_13984_, _13983_, _13978_);
  or _65617_ (_13985_, _13984_, _06509_);
  or _65618_ (_13986_, _13985_, _13982_);
  and _65619_ (_13987_, _09087_, _07969_);
  or _65620_ (_13988_, _13908_, _09107_);
  or _65621_ (_13989_, _13988_, _13987_);
  and _65622_ (_13990_, _13989_, _09112_);
  and _65623_ (_13991_, _13990_, _13986_);
  nor _65624_ (_13992_, _09095_, _13907_);
  or _65625_ (_13993_, _13992_, _13908_);
  and _65626_ (_13994_, _13993_, _06602_);
  or _65627_ (_13995_, _13994_, _06639_);
  or _65628_ (_13996_, _13995_, _13991_);
  or _65629_ (_13997_, _13921_, _07048_);
  and _65630_ (_13998_, _13997_, _05990_);
  and _65631_ (_13999_, _13998_, _13996_);
  and _65632_ (_14000_, _13918_, _05989_);
  or _65633_ (_14001_, _14000_, _06646_);
  or _65634_ (_14002_, _14001_, _13999_);
  and _65635_ (_14003_, _08605_, _07969_);
  or _65636_ (_14004_, _13908_, _06651_);
  or _65637_ (_14005_, _14004_, _14003_);
  and _65638_ (_14006_, _14005_, _01442_);
  and _65639_ (_14007_, _14006_, _14002_);
  or _65640_ (_14008_, _14007_, _13906_);
  and _65641_ (_41517_, _14008_, _43634_);
  not _65642_ (_14009_, \oc8051_golden_model_1.SP [7]);
  nor _65643_ (_14010_, _01442_, _14009_);
  and _65644_ (_14011_, _07688_, \oc8051_golden_model_1.SP [4]);
  and _65645_ (_14012_, _14011_, \oc8051_golden_model_1.SP [5]);
  and _65646_ (_14013_, _14012_, \oc8051_golden_model_1.SP [6]);
  or _65647_ (_14014_, _14013_, \oc8051_golden_model_1.SP [7]);
  nand _65648_ (_14015_, _14013_, \oc8051_golden_model_1.SP [7]);
  and _65649_ (_14016_, _14015_, _14014_);
  or _65650_ (_14017_, _14016_, _07367_);
  nor _65651_ (_14018_, _08004_, _14009_);
  and _65652_ (_14019_, _09096_, _08004_);
  or _65653_ (_14020_, _14019_, _14018_);
  and _65654_ (_14021_, _14020_, _06615_);
  not _65655_ (_14022_, _06334_);
  not _65656_ (_14023_, _08004_);
  nor _65657_ (_14024_, _08107_, _14023_);
  and _65658_ (_14025_, _06471_, _06002_);
  or _65659_ (_14026_, _14018_, _14025_);
  or _65660_ (_14027_, _14026_, _14024_);
  and _65661_ (_14028_, _14027_, _14022_);
  and _65662_ (_14029_, _08791_, _08004_);
  or _65663_ (_14030_, _14029_, _14018_);
  or _65664_ (_14031_, _14030_, _07275_);
  and _65665_ (_14032_, _08004_, \oc8051_golden_model_1.ACC [7]);
  or _65666_ (_14033_, _14032_, _14018_);
  or _65667_ (_14034_, _14033_, _07260_);
  or _65668_ (_14035_, _07259_, \oc8051_golden_model_1.SP [7]);
  and _65669_ (_14036_, _14035_, _07564_);
  and _65670_ (_14037_, _14036_, _14034_);
  and _65671_ (_14038_, _14016_, _06816_);
  or _65672_ (_14039_, _14038_, _06474_);
  or _65673_ (_14040_, _14039_, _14037_);
  and _65674_ (_14041_, _14040_, _06052_);
  and _65675_ (_14042_, _14041_, _14031_);
  and _65676_ (_14043_, _14016_, _07692_);
  or _65677_ (_14044_, _14043_, _06410_);
  or _65678_ (_14045_, _14044_, _14042_);
  not _65679_ (_14046_, \oc8051_golden_model_1.SP [6]);
  not _65680_ (_14047_, \oc8051_golden_model_1.SP [5]);
  not _65681_ (_14048_, \oc8051_golden_model_1.SP [4]);
  and _65682_ (_14049_, _08699_, _14048_);
  and _65683_ (_14050_, _14049_, _14047_);
  and _65684_ (_14051_, _14050_, _14046_);
  and _65685_ (_14052_, _14051_, _06342_);
  nor _65686_ (_14053_, _14052_, _14009_);
  and _65687_ (_14054_, _14052_, _14009_);
  nor _65688_ (_14055_, _14054_, _14053_);
  nand _65689_ (_14056_, _14055_, _06410_);
  and _65690_ (_14057_, _14056_, _14045_);
  or _65691_ (_14058_, _14057_, _06417_);
  or _65692_ (_14059_, _14033_, _06426_);
  and _65693_ (_14060_, _14059_, _07394_);
  and _65694_ (_14061_, _14060_, _14058_);
  nor _65695_ (_14062_, _06806_, _05992_);
  and _65696_ (_14063_, _14012_, \oc8051_golden_model_1.SP [0]);
  and _65697_ (_14064_, _14063_, \oc8051_golden_model_1.SP [6]);
  nor _65698_ (_14065_, _14064_, _14009_);
  and _65699_ (_14066_, _14064_, _14009_);
  or _65700_ (_14067_, _14066_, _14065_);
  and _65701_ (_14068_, _14067_, _06351_);
  or _65702_ (_14069_, _14068_, _14062_);
  or _65703_ (_14070_, _14069_, _14061_);
  or _65704_ (_14071_, _14016_, _07597_);
  and _65705_ (_14072_, _14071_, _14070_);
  and _65706_ (_14073_, _14072_, _06327_);
  or _65707_ (_14074_, _14073_, _14028_);
  and _65708_ (_14075_, _08778_, _08004_);
  or _65709_ (_14076_, _14018_, _06333_);
  or _65710_ (_14077_, _14076_, _14075_);
  and _65711_ (_14078_, _14077_, _06313_);
  and _65712_ (_14079_, _14078_, _14074_);
  and _65713_ (_14080_, _09076_, _08004_);
  or _65714_ (_14081_, _14080_, _14018_);
  and _65715_ (_14082_, _14081_, _06037_);
  or _65716_ (_14083_, _14082_, _06277_);
  or _65717_ (_14084_, _14083_, _14079_);
  and _65718_ (_14085_, _08880_, _08004_);
  or _65719_ (_14086_, _14085_, _14018_);
  or _65720_ (_14087_, _14086_, _06278_);
  and _65721_ (_14088_, _14087_, _14084_);
  or _65722_ (_14089_, _14088_, _06275_);
  or _65723_ (_14090_, _14016_, _06009_);
  and _65724_ (_14091_, _14090_, _14089_);
  or _65725_ (_14092_, _14091_, _06502_);
  and _65726_ (_14093_, _09090_, _08004_);
  or _65727_ (_14094_, _14018_, _07334_);
  or _65728_ (_14095_, _14094_, _14093_);
  and _65729_ (_14096_, _14095_, _07337_);
  and _65730_ (_14097_, _14096_, _14092_);
  or _65731_ (_14098_, _14097_, _14021_);
  and _65732_ (_14099_, _14098_, _07339_);
  or _65733_ (_14100_, _14018_, _08110_);
  and _65734_ (_14101_, _14086_, _06507_);
  and _65735_ (_14102_, _14101_, _14100_);
  or _65736_ (_14103_, _14102_, _14099_);
  and _65737_ (_14104_, _14103_, _12805_);
  and _65738_ (_14105_, _14033_, _06610_);
  and _65739_ (_14106_, _14105_, _14100_);
  and _65740_ (_14107_, _14016_, _07330_);
  or _65741_ (_14108_, _14107_, _06509_);
  or _65742_ (_14109_, _14108_, _14106_);
  or _65743_ (_14110_, _14109_, _14104_);
  and _65744_ (_14111_, _09087_, _08004_);
  or _65745_ (_14112_, _14111_, _14018_);
  or _65746_ (_14113_, _14112_, _09107_);
  and _65747_ (_14114_, _14113_, _14110_);
  or _65748_ (_14115_, _14114_, _06602_);
  not _65749_ (_14116_, _06621_);
  nor _65750_ (_14117_, _09095_, _14023_);
  or _65751_ (_14118_, _14018_, _09112_);
  or _65752_ (_14119_, _14118_, _14117_);
  and _65753_ (_14120_, _14119_, _14116_);
  and _65754_ (_14121_, _14120_, _14115_);
  or _65755_ (_14122_, _14051_, \oc8051_golden_model_1.SP [7]);
  nand _65756_ (_14123_, _14051_, \oc8051_golden_model_1.SP [7]);
  and _65757_ (_14124_, _14123_, _14122_);
  and _65758_ (_14125_, _14124_, _06621_);
  or _65759_ (_14126_, _14125_, _07350_);
  or _65760_ (_14127_, _14126_, _14121_);
  or _65761_ (_14128_, _14016_, _06016_);
  and _65762_ (_14129_, _14128_, _14127_);
  or _65763_ (_14130_, _14129_, _06361_);
  or _65764_ (_14131_, _14124_, _06362_);
  and _65765_ (_14132_, _14131_, _07048_);
  and _65766_ (_14133_, _14132_, _14130_);
  and _65767_ (_14134_, _14030_, _06639_);
  or _65768_ (_14135_, _14134_, _07783_);
  or _65769_ (_14136_, _14135_, _14133_);
  and _65770_ (_14137_, _14136_, _14017_);
  or _65771_ (_14138_, _14137_, _06646_);
  and _65772_ (_14139_, _08605_, _08004_);
  or _65773_ (_14140_, _14018_, _06651_);
  or _65774_ (_14141_, _14140_, _14139_);
  and _65775_ (_14142_, _14141_, _01442_);
  and _65776_ (_14143_, _14142_, _14138_);
  or _65777_ (_14144_, _14143_, _14010_);
  and _65778_ (_41519_, _14144_, _43634_);
  not _65779_ (_14145_, _07962_);
  and _65780_ (_14146_, _14145_, \oc8051_golden_model_1.SBUF [7]);
  and _65781_ (_14147_, _09096_, _07962_);
  or _65782_ (_14148_, _14147_, _14146_);
  and _65783_ (_14149_, _14148_, _06615_);
  nor _65784_ (_14150_, _08107_, _14145_);
  or _65785_ (_14151_, _14150_, _14146_);
  or _65786_ (_14152_, _14151_, _06327_);
  and _65787_ (_14153_, _08791_, _07962_);
  or _65788_ (_14154_, _14153_, _14146_);
  or _65789_ (_14155_, _14154_, _07275_);
  and _65790_ (_14156_, _07962_, \oc8051_golden_model_1.ACC [7]);
  or _65791_ (_14157_, _14156_, _14146_);
  and _65792_ (_14158_, _14157_, _07259_);
  and _65793_ (_14159_, _07260_, \oc8051_golden_model_1.SBUF [7]);
  or _65794_ (_14160_, _14159_, _06474_);
  or _65795_ (_14161_, _14160_, _14158_);
  and _65796_ (_14162_, _14161_, _06772_);
  and _65797_ (_14163_, _14162_, _14155_);
  and _65798_ (_14164_, _14151_, _06410_);
  or _65799_ (_14165_, _14164_, _14163_);
  and _65800_ (_14166_, _14165_, _06426_);
  and _65801_ (_14167_, _14157_, _06417_);
  or _65802_ (_14168_, _14167_, _10153_);
  or _65803_ (_14169_, _14168_, _14166_);
  and _65804_ (_14170_, _14169_, _14152_);
  or _65805_ (_14171_, _14170_, _09572_);
  and _65806_ (_14172_, _08778_, _07962_);
  or _65807_ (_14173_, _14146_, _06333_);
  or _65808_ (_14174_, _14173_, _14172_);
  and _65809_ (_14175_, _14174_, _06313_);
  and _65810_ (_14176_, _14175_, _14171_);
  and _65811_ (_14177_, _09076_, _07962_);
  or _65812_ (_14178_, _14177_, _14146_);
  and _65813_ (_14179_, _14178_, _06037_);
  or _65814_ (_14180_, _14179_, _06277_);
  or _65815_ (_14181_, _14180_, _14176_);
  and _65816_ (_14182_, _08880_, _07962_);
  or _65817_ (_14183_, _14182_, _14146_);
  or _65818_ (_14184_, _14183_, _06278_);
  and _65819_ (_14185_, _14184_, _14181_);
  or _65820_ (_14186_, _14185_, _06502_);
  and _65821_ (_14187_, _09090_, _07962_);
  or _65822_ (_14188_, _14146_, _07334_);
  or _65823_ (_14189_, _14188_, _14187_);
  and _65824_ (_14190_, _14189_, _07337_);
  and _65825_ (_14191_, _14190_, _14186_);
  or _65826_ (_14192_, _14191_, _14149_);
  and _65827_ (_14193_, _14192_, _07339_);
  or _65828_ (_14194_, _14146_, _08110_);
  and _65829_ (_14195_, _14183_, _06507_);
  and _65830_ (_14196_, _14195_, _14194_);
  or _65831_ (_14197_, _14196_, _14193_);
  and _65832_ (_14198_, _14197_, _07331_);
  and _65833_ (_14199_, _14157_, _06610_);
  and _65834_ (_14200_, _14199_, _14194_);
  or _65835_ (_14201_, _14200_, _06509_);
  or _65836_ (_14202_, _14201_, _14198_);
  and _65837_ (_14203_, _09087_, _07962_);
  or _65838_ (_14204_, _14146_, _09107_);
  or _65839_ (_14205_, _14204_, _14203_);
  and _65840_ (_14206_, _14205_, _09112_);
  and _65841_ (_14207_, _14206_, _14202_);
  nor _65842_ (_14208_, _09095_, _14145_);
  or _65843_ (_14209_, _14208_, _14146_);
  and _65844_ (_14210_, _14209_, _06602_);
  or _65845_ (_14211_, _14210_, _06639_);
  or _65846_ (_14212_, _14211_, _14207_);
  or _65847_ (_14213_, _14154_, _07048_);
  and _65848_ (_14214_, _14213_, _06651_);
  and _65849_ (_14215_, _14214_, _14212_);
  and _65850_ (_14216_, _08605_, _07962_);
  or _65851_ (_14217_, _14216_, _14146_);
  and _65852_ (_14218_, _14217_, _06646_);
  or _65853_ (_14219_, _14218_, _01446_);
  or _65854_ (_14220_, _14219_, _14215_);
  or _65855_ (_14221_, _01442_, \oc8051_golden_model_1.SBUF [7]);
  and _65856_ (_14222_, _14221_, _43634_);
  and _65857_ (_41520_, _14222_, _14220_);
  nor _65858_ (_14223_, _01442_, _10967_);
  nor _65859_ (_14224_, _08640_, _10967_);
  and _65860_ (_14225_, _08668_, _08640_);
  or _65861_ (_14226_, _14225_, _14224_);
  or _65862_ (_14227_, _14226_, _05990_);
  nor _65863_ (_14228_, _10796_, _08688_);
  or _65864_ (_14229_, _14228_, _11152_);
  or _65865_ (_14230_, _14229_, _10794_);
  or _65866_ (_14231_, _14230_, _11127_);
  nor _65867_ (_14232_, _08014_, _10967_);
  and _65868_ (_14233_, _09096_, _08014_);
  or _65869_ (_14234_, _14233_, _14232_);
  and _65870_ (_14235_, _14234_, _06615_);
  and _65871_ (_14236_, _09076_, _08014_);
  or _65872_ (_14237_, _14236_, _14232_);
  and _65873_ (_14238_, _14237_, _06037_);
  not _65874_ (_14239_, _08014_);
  nor _65875_ (_14240_, _08107_, _14239_);
  or _65876_ (_14241_, _14240_, _14232_);
  or _65877_ (_14242_, _14241_, _06327_);
  and _65878_ (_14243_, _10868_, _10863_);
  nor _65879_ (_14244_, _14243_, _10861_);
  nand _65880_ (_14245_, _10916_, _10863_);
  or _65881_ (_14246_, _14245_, _10914_);
  and _65882_ (_14247_, _14246_, _14244_);
  and _65883_ (_14248_, _10857_, _08778_);
  or _65884_ (_14249_, _14248_, _10854_);
  or _65885_ (_14250_, _14249_, _14247_);
  not _65886_ (_14251_, _06444_);
  not _65887_ (_14252_, _06445_);
  nor _65888_ (_14253_, _13037_, _14252_);
  and _65889_ (_14254_, _12367_, _12366_);
  not _65890_ (_14255_, _12374_);
  or _65891_ (_14256_, _12376_, _14255_);
  and _65892_ (_14257_, _14256_, _12370_);
  or _65893_ (_14258_, _14257_, _14254_);
  and _65894_ (_14259_, _14258_, _12363_);
  and _65895_ (_14260_, _12352_, _12350_);
  and _65896_ (_14261_, _12356_, _12353_);
  nand _65897_ (_14262_, _14261_, _14260_);
  and _65898_ (_14263_, _12359_, _12357_);
  or _65899_ (_14264_, _14263_, _14262_);
  nand _65900_ (_14265_, _14264_, _14260_);
  and _65901_ (_14266_, _14265_, _08822_);
  or _65902_ (_14267_, _14266_, _14259_);
  and _65903_ (_14268_, _14267_, _12379_);
  or _65904_ (_14269_, _14268_, _06473_);
  not _65905_ (_14270_, _12609_);
  and _65906_ (_14271_, _12603_, _12600_);
  and _65907_ (_14272_, _12597_, _12596_);
  or _65908_ (_14273_, _14272_, _12606_);
  or _65909_ (_14274_, _14273_, _14271_);
  and _65910_ (_14275_, _14274_, _12593_);
  or _65911_ (_14276_, _12590_, _12586_);
  and _65912_ (_14277_, _12584_, _14276_);
  and _65913_ (_14278_, _14277_, _12585_);
  or _65914_ (_14279_, _12579_, _12581_);
  and _65915_ (_14280_, _14279_, _08108_);
  or _65916_ (_14281_, _14280_, _14278_);
  or _65917_ (_14282_, _14281_, _14275_);
  and _65918_ (_14283_, _14282_, _14270_);
  or _65919_ (_14284_, _14283_, _12574_);
  and _65920_ (_14285_, _08791_, _08014_);
  or _65921_ (_14286_, _14285_, _14232_);
  or _65922_ (_14287_, _14286_, _07275_);
  and _65923_ (_14288_, _08014_, \oc8051_golden_model_1.ACC [7]);
  or _65924_ (_14289_, _14288_, _14232_);
  and _65925_ (_14290_, _14289_, _07259_);
  nor _65926_ (_14291_, _07259_, _10967_);
  or _65927_ (_14292_, _14291_, _06474_);
  or _65928_ (_14293_, _14292_, _14290_);
  and _65929_ (_14294_, _14293_, _10730_);
  and _65930_ (_14295_, _14294_, _14287_);
  nor _65931_ (_14296_, _10750_, _10730_);
  not _65932_ (_14297_, _06418_);
  or _65933_ (_14298_, _12501_, _14297_);
  or _65934_ (_14299_, _14298_, _14296_);
  or _65935_ (_14300_, _14299_, _14295_);
  and _65936_ (_14301_, _08672_, _08640_);
  or _65937_ (_14302_, _14301_, _14224_);
  or _65938_ (_14303_, _14302_, _06357_);
  or _65939_ (_14304_, _14241_, _06772_);
  and _65940_ (_14305_, _14304_, _14303_);
  and _65941_ (_14306_, _14305_, _14300_);
  or _65942_ (_14307_, _14306_, _06417_);
  or _65943_ (_14308_, _14289_, _06426_);
  nor _65944_ (_14309_, _12560_, _06352_);
  and _65945_ (_14310_, _14309_, _14308_);
  and _65946_ (_14311_, _14310_, _14307_);
  and _65947_ (_14312_, _14226_, _06352_);
  or _65948_ (_14313_, _14312_, _12611_);
  or _65949_ (_14314_, _14313_, _14311_);
  and _65950_ (_14315_, _14314_, _14284_);
  or _65951_ (_14316_, _14315_, _06472_);
  and _65952_ (_14317_, _14316_, _06500_);
  and _65953_ (_14318_, _14317_, _14269_);
  nand _65954_ (_14319_, _08358_, \oc8051_golden_model_1.ACC [3]);
  nor _65955_ (_14320_, _08502_, \oc8051_golden_model_1.ACC [2]);
  nor _65956_ (_14321_, _08358_, \oc8051_golden_model_1.ACC [3]);
  or _65957_ (_14322_, _14321_, _14320_);
  and _65958_ (_14323_, _14322_, _14319_);
  nor _65959_ (_14324_, _08403_, \oc8051_golden_model_1.ACC [1]);
  nor _65960_ (_14325_, _08453_, _06071_);
  nor _65961_ (_14326_, _14325_, _10579_);
  or _65962_ (_14327_, _14326_, _14324_);
  and _65963_ (_14328_, _14327_, _12620_);
  or _65964_ (_14329_, _14328_, _14323_);
  and _65965_ (_14330_, _14329_, _12629_);
  nand _65966_ (_14331_, _08307_, \oc8051_golden_model_1.ACC [5]);
  nor _65967_ (_14332_, _08598_, \oc8051_golden_model_1.ACC [4]);
  nor _65968_ (_14333_, _08307_, \oc8051_golden_model_1.ACC [5]);
  or _65969_ (_14334_, _14333_, _14332_);
  and _65970_ (_14335_, _14334_, _14331_);
  and _65971_ (_14336_, _14335_, _12628_);
  nor _65972_ (_14337_, _08109_, \oc8051_golden_model_1.ACC [7]);
  or _65973_ (_14338_, _08211_, \oc8051_golden_model_1.ACC [6]);
  nor _65974_ (_14339_, _14338_, _09096_);
  or _65975_ (_14340_, _14339_, _14337_);
  or _65976_ (_14341_, _14340_, _14336_);
  or _65977_ (_14342_, _14341_, _14330_);
  nor _65978_ (_14343_, _12630_, _06500_);
  and _65979_ (_14344_, _14343_, _14342_);
  or _65980_ (_14345_, _14344_, _14318_);
  and _65981_ (_14346_, _14345_, _12349_);
  and _65982_ (_14347_, _06238_, _08688_);
  or _65983_ (_14348_, _06397_, \oc8051_golden_model_1.ACC [6]);
  nor _65984_ (_14349_, _14348_, _11070_);
  or _65985_ (_14350_, _14349_, _14347_);
  nand _65986_ (_14351_, _06685_, \oc8051_golden_model_1.ACC [5]);
  nor _65987_ (_14352_, _06685_, \oc8051_golden_model_1.ACC [5]);
  nor _65988_ (_14353_, _07093_, \oc8051_golden_model_1.ACC [4]);
  or _65989_ (_14354_, _14353_, _14352_);
  and _65990_ (_14355_, _14354_, _14351_);
  and _65991_ (_14356_, _14355_, _12646_);
  or _65992_ (_14357_, _14356_, _14350_);
  and _65993_ (_14358_, _06310_, \oc8051_golden_model_1.ACC [0]);
  nor _65994_ (_14359_, _14358_, _11352_);
  or _65995_ (_14360_, _14359_, _11353_);
  and _65996_ (_14361_, _14360_, _12639_);
  nand _65997_ (_14362_, _06269_, \oc8051_golden_model_1.ACC [3]);
  nor _65998_ (_14363_, _06269_, \oc8051_golden_model_1.ACC [3]);
  nor _65999_ (_14364_, _06727_, \oc8051_golden_model_1.ACC [2]);
  or _66000_ (_14365_, _14364_, _14363_);
  and _66001_ (_14366_, _14365_, _14362_);
  or _66002_ (_14367_, _14366_, _14361_);
  and _66003_ (_14368_, _14367_, _12647_);
  or _66004_ (_14369_, _14368_, _14357_);
  nor _66005_ (_14370_, _12648_, _12349_);
  and _66006_ (_14371_, _14370_, _14369_);
  or _66007_ (_14372_, _14371_, _12347_);
  or _66008_ (_14373_, _14372_, _14346_);
  nand _66009_ (_14374_, _12347_, \oc8051_golden_model_1.PSW [7]);
  and _66010_ (_14375_, _14374_, _06346_);
  and _66011_ (_14376_, _14375_, _14373_);
  or _66012_ (_14377_, _14224_, _08809_);
  and _66013_ (_14378_, _14302_, _06345_);
  and _66014_ (_14379_, _14378_, _14377_);
  nor _66015_ (_14380_, _14379_, _14376_);
  nor _66016_ (_14381_, _14380_, _06404_);
  and _66017_ (_14382_, _06404_, \oc8051_golden_model_1.PSW [7]);
  and _66018_ (_14383_, _14382_, _13037_);
  or _66019_ (_14384_, _14383_, _14381_);
  nor _66020_ (_14385_, _09606_, _06445_);
  and _66021_ (_14386_, _14385_, _14384_);
  or _66022_ (_14387_, _14386_, _14253_);
  and _66023_ (_14388_, _14387_, _14251_);
  and _66024_ (_14389_, _07577_, _06038_);
  and _66025_ (_14390_, _06480_, _06038_);
  or _66026_ (_14391_, _14390_, _14389_);
  or _66027_ (_14392_, _13037_, \oc8051_golden_model_1.PSW [7]);
  and _66028_ (_14393_, _14392_, _06444_);
  or _66029_ (_14394_, _14393_, _14391_);
  or _66030_ (_14395_, _14394_, _14388_);
  not _66031_ (_14396_, _06910_);
  and _66032_ (_14397_, _10803_, _10799_);
  nor _66033_ (_14398_, _14397_, _10797_);
  nand _66034_ (_14399_, _10845_, _10799_);
  or _66035_ (_14400_, _14399_, _10843_);
  and _66036_ (_14401_, _14400_, _14398_);
  or _66037_ (_14402_, _14401_, _10794_);
  and _66038_ (_14403_, _14402_, _14396_);
  or _66039_ (_14404_, _14403_, _10784_);
  and _66040_ (_14405_, _14404_, _14395_);
  and _66041_ (_14406_, _14402_, _06910_);
  or _66042_ (_14407_, _14406_, _10853_);
  or _66043_ (_14408_, _14407_, _14405_);
  and _66044_ (_14409_, _14408_, _14250_);
  or _66045_ (_14410_, _14409_, _06453_);
  and _66046_ (_14411_, _10635_, _08212_);
  and _66047_ (_14412_, _14411_, _08110_);
  and _66048_ (_14413_, _10638_, _10631_);
  nor _66049_ (_14414_, _14413_, _10629_);
  nand _66050_ (_14415_, _10684_, _10631_);
  or _66051_ (_14416_, _14415_, _10681_);
  and _66052_ (_14417_, _14416_, _14414_);
  or _66053_ (_14418_, _14417_, _14412_);
  or _66054_ (_14419_, _14418_, _06458_);
  and _66055_ (_14420_, _14419_, _10624_);
  and _66056_ (_14421_, _14420_, _14410_);
  and _66057_ (_14422_, _10927_, _08024_);
  and _66058_ (_14423_, _10939_, _10935_);
  nor _66059_ (_14424_, _14423_, _10933_);
  and _66060_ (_14425_, _10990_, _10935_);
  not _66061_ (_14426_, _14425_);
  or _66062_ (_14427_, _14426_, _10988_);
  and _66063_ (_14428_, _14427_, _14424_);
  or _66064_ (_14429_, _14428_, _14422_);
  and _66065_ (_14430_, _14429_, _10623_);
  or _66066_ (_14431_, _14430_, _10153_);
  or _66067_ (_14432_, _14431_, _14421_);
  and _66068_ (_14433_, _14432_, _14242_);
  or _66069_ (_14434_, _14433_, _09572_);
  and _66070_ (_14435_, _08778_, _08014_);
  or _66071_ (_14436_, _14232_, _06333_);
  or _66072_ (_14437_, _14436_, _14435_);
  and _66073_ (_14438_, _14437_, _06313_);
  and _66074_ (_14439_, _14438_, _14434_);
  or _66075_ (_14440_, _14439_, _14238_);
  nor _66076_ (_14441_, _10166_, _06401_);
  and _66077_ (_14442_, _14441_, _14440_);
  nor _66078_ (_14443_, _13037_, _10967_);
  and _66079_ (_14444_, _14443_, _06401_);
  or _66080_ (_14445_, _14444_, _06277_);
  or _66081_ (_14446_, _14445_, _14442_);
  and _66082_ (_14447_, _08880_, _08014_);
  or _66083_ (_14448_, _14447_, _14232_);
  or _66084_ (_14449_, _14448_, _06278_);
  and _66085_ (_14450_, _14449_, _14446_);
  or _66086_ (_14451_, _14450_, _06400_);
  nand _66087_ (_14452_, _13037_, _10967_);
  or _66088_ (_14453_, _14452_, _06958_);
  and _66089_ (_14454_, _14453_, _14451_);
  or _66090_ (_14455_, _14454_, _06502_);
  and _66091_ (_14456_, _09090_, _08014_);
  or _66092_ (_14457_, _14232_, _07334_);
  or _66093_ (_14458_, _14457_, _14456_);
  and _66094_ (_14459_, _14458_, _07337_);
  and _66095_ (_14460_, _14459_, _14455_);
  or _66096_ (_14461_, _14460_, _14235_);
  and _66097_ (_14462_, _14461_, _07339_);
  or _66098_ (_14463_, _14232_, _08110_);
  and _66099_ (_14464_, _14448_, _06507_);
  and _66100_ (_14465_, _14464_, _14463_);
  or _66101_ (_14466_, _14465_, _14462_);
  and _66102_ (_14467_, _14466_, _07331_);
  and _66103_ (_14468_, _14289_, _06610_);
  and _66104_ (_14469_, _14468_, _14463_);
  or _66105_ (_14470_, _14469_, _06509_);
  or _66106_ (_14471_, _14470_, _14467_);
  and _66107_ (_14472_, _09087_, _08014_);
  or _66108_ (_14473_, _14232_, _09107_);
  or _66109_ (_14474_, _14473_, _14472_);
  and _66110_ (_14475_, _14474_, _09112_);
  and _66111_ (_14476_, _14475_, _14471_);
  nor _66112_ (_14477_, _09095_, _14239_);
  or _66113_ (_14478_, _14477_, _14232_);
  and _66114_ (_14479_, _14478_, _06602_);
  or _66115_ (_14480_, _14479_, _11130_);
  or _66116_ (_14481_, _14480_, _14476_);
  and _66117_ (_14482_, _14481_, _14231_);
  or _66118_ (_14483_, _14482_, _11129_);
  nor _66119_ (_14484_, _10860_, _08688_);
  or _66120_ (_14485_, _14484_, _11180_);
  or _66121_ (_14486_, _11158_, _14248_);
  or _66122_ (_14487_, _14486_, _14485_);
  and _66123_ (_14488_, _14487_, _06601_);
  and _66124_ (_14489_, _14488_, _14483_);
  nor _66125_ (_14490_, _10628_, _08688_);
  or _66126_ (_14491_, _14490_, _11210_);
  or _66127_ (_14492_, _14491_, _14412_);
  and _66128_ (_14493_, _14492_, _06600_);
  or _66129_ (_14494_, _14493_, _11186_);
  or _66130_ (_14495_, _14494_, _14489_);
  nor _66131_ (_14496_, _10932_, _08688_);
  or _66132_ (_14497_, _14496_, _11239_);
  or _66133_ (_14498_, _14422_, _11218_);
  or _66134_ (_14499_, _14498_, _14497_);
  and _66135_ (_14500_, _14499_, _11217_);
  and _66136_ (_14501_, _14500_, _14495_);
  nand _66137_ (_14502_, _11216_, \oc8051_golden_model_1.ACC [7]);
  nand _66138_ (_14503_, _14502_, _11248_);
  or _66139_ (_14504_, _14503_, _14501_);
  and _66140_ (_14505_, _11283_, _11039_);
  nor _66141_ (_14506_, _11251_, _10612_);
  nor _66142_ (_14507_, _14506_, _10607_);
  or _66143_ (_14508_, _14507_, _11248_);
  or _66144_ (_14509_, _14508_, _14505_);
  and _66145_ (_14510_, _14509_, _14504_);
  or _66146_ (_14511_, _14510_, _11290_);
  and _66147_ (_14512_, _11325_, _11059_);
  nor _66148_ (_14513_, _11293_, _11058_);
  nor _66149_ (_14514_, _14513_, _11057_);
  or _66150_ (_14515_, _14514_, _11292_);
  or _66151_ (_14516_, _14515_, _14512_);
  and _66152_ (_14517_, _14516_, _06364_);
  and _66153_ (_14518_, _14517_, _14511_);
  not _66154_ (_14519_, _09095_);
  not _66155_ (_14520_, _09094_);
  nand _66156_ (_14521_, _10598_, _14520_);
  and _66157_ (_14522_, _14521_, _06363_);
  and _66158_ (_14523_, _14522_, _14519_);
  or _66159_ (_14524_, _14523_, _10566_);
  or _66160_ (_14525_, _14524_, _14518_);
  not _66161_ (_14526_, _11069_);
  nor _66162_ (_14527_, _11368_, _11068_);
  nor _66163_ (_14528_, _14527_, _10567_);
  nand _66164_ (_14529_, _14528_, _14526_);
  and _66165_ (_14530_, _14529_, _14525_);
  or _66166_ (_14531_, _14530_, _06639_);
  nor _66167_ (_14532_, _14286_, _07048_);
  nor _66168_ (_14533_, _14532_, _11382_);
  and _66169_ (_14534_, _14533_, _14531_);
  and _66170_ (_14535_, _11382_, \oc8051_golden_model_1.ACC [0]);
  or _66171_ (_14536_, _14535_, _05989_);
  or _66172_ (_14537_, _14536_, _14534_);
  and _66173_ (_14538_, _14537_, _14227_);
  or _66174_ (_14539_, _14538_, _06646_);
  and _66175_ (_14540_, _08605_, _08014_);
  or _66176_ (_14541_, _14232_, _06651_);
  or _66177_ (_14542_, _14541_, _14540_);
  and _66178_ (_14543_, _14542_, _01442_);
  and _66179_ (_14544_, _14543_, _14539_);
  or _66180_ (_14545_, _14544_, _14223_);
  and _66181_ (_41521_, _14545_, _43634_);
  or _66182_ (_14546_, _00000_, \oc8051_golden_model_1.P0INREG [7]);
  or _66183_ (_14547_, _07543_, p0_in[7]);
  and _66184_ (_41522_, _14547_, _14546_);
  or _66185_ (_14548_, _00000_, \oc8051_golden_model_1.P1INREG [7]);
  or _66186_ (_14549_, _07543_, p1_in[7]);
  and _66187_ (_41523_, _14549_, _14548_);
  or _66188_ (_14550_, _00000_, \oc8051_golden_model_1.P2INREG [7]);
  or _66189_ (_14551_, _07543_, p2_in[7]);
  and _66190_ (_41525_, _14551_, _14550_);
  or _66191_ (_14552_, _00000_, \oc8051_golden_model_1.P3INREG [7]);
  or _66192_ (_14553_, _07543_, p3_in[7]);
  and _66193_ (_41526_, _14553_, _14552_);
  and _66194_ (_14554_, _07631_, _07382_);
  nor _66195_ (_14555_, _14554_, _07633_);
  nor _66196_ (_14556_, _07798_, _07632_);
  nor _66197_ (_14557_, _14556_, _07941_);
  and _66198_ (_14558_, _14557_, _07631_);
  and _66199_ (_14559_, _14558_, _14555_);
  not _66200_ (_14560_, _14559_);
  nand _66201_ (_14561_, _05998_, _05701_);
  nand _66202_ (_14562_, _12622_, _09113_);
  or _66203_ (_14563_, _08453_, _09008_);
  and _66204_ (_14564_, _08453_, _09008_);
  not _66205_ (_14565_, _14564_);
  and _66206_ (_14566_, _14565_, _14563_);
  and _66207_ (_14567_, _14566_, _07335_);
  and _66208_ (_14568_, _06039_, \oc8051_golden_model_1.PC [0]);
  nor _66209_ (_14569_, _12955_, _07967_);
  or _66210_ (_14570_, _14569_, _08629_);
  nor _66211_ (_14571_, _08453_, _08782_);
  nand _66212_ (_14572_, _08687_, _07250_);
  nand _66213_ (_14573_, _06816_, _05701_);
  or _66214_ (_14574_, _06816_, \oc8051_golden_model_1.ACC [0]);
  and _66215_ (_14575_, _14574_, _14573_);
  nor _66216_ (_14576_, _14575_, _08687_);
  nor _66217_ (_14577_, _14576_, _07276_);
  and _66218_ (_14578_, _14577_, _14572_);
  or _66219_ (_14579_, _14578_, _14571_);
  and _66220_ (_14580_, _14579_, _08670_);
  nand _66221_ (_14581_, _12955_, _12933_);
  and _66222_ (_14582_, _14581_, _07274_);
  or _66223_ (_14583_, _14582_, _07692_);
  or _66224_ (_14584_, _14583_, _14580_);
  nor _66225_ (_14585_, _06052_, \oc8051_golden_model_1.PC [0]);
  nor _66226_ (_14586_, _14585_, _07284_);
  and _66227_ (_14587_, _14586_, _14584_);
  and _66228_ (_14588_, _07284_, _07250_);
  or _66229_ (_14589_, _14588_, _07294_);
  or _66230_ (_14590_, _14589_, _14587_);
  and _66231_ (_14591_, _14590_, _14570_);
  or _66232_ (_14592_, _14591_, _06351_);
  or _66233_ (_14593_, _08453_, _07394_);
  and _66234_ (_14594_, _14593_, _06349_);
  and _66235_ (_14595_, _14594_, _14592_);
  nor _66236_ (_14596_, _12956_, _06349_);
  and _66237_ (_14597_, _14596_, _14581_);
  or _66238_ (_14598_, _14597_, _14595_);
  and _66239_ (_14599_, _14598_, _06049_);
  nor _66240_ (_14600_, _06049_, _05701_);
  or _66241_ (_14601_, _06441_, _14600_);
  or _66242_ (_14602_, _14601_, _14599_);
  or _66243_ (_14603_, _08453_, _06448_);
  and _66244_ (_14604_, _14603_, _14602_);
  or _66245_ (_14605_, _14604_, _07309_);
  and _66246_ (_14606_, _09447_, _06366_);
  nand _66247_ (_14607_, _08450_, _07309_);
  or _66248_ (_14608_, _14607_, _14606_);
  and _66249_ (_14609_, _14608_, _08821_);
  and _66250_ (_14610_, _14609_, _14605_);
  and _66251_ (_14611_, _07967_, \oc8051_golden_model_1.PSW [7]);
  or _66252_ (_14612_, _14611_, _14569_);
  and _66253_ (_14613_, _14612_, _07308_);
  or _66254_ (_14614_, _14613_, _14610_);
  and _66255_ (_14615_, _14614_, _07745_);
  or _66256_ (_14616_, _14615_, _14568_);
  and _66257_ (_14617_, _14616_, _08836_);
  and _66258_ (_14618_, _08832_, _07250_);
  or _66259_ (_14619_, _14618_, _08838_);
  or _66260_ (_14620_, _14619_, _14617_);
  or _66261_ (_14621_, _09447_, _08844_);
  and _66262_ (_14622_, _14621_, _08842_);
  and _66263_ (_14623_, _14622_, _14620_);
  and _66264_ (_14624_, _08879_, _07250_);
  and _66265_ (_14625_, _09023_, \oc8051_golden_model_1.PSW [0]);
  and _66266_ (_14626_, _09026_, \oc8051_golden_model_1.IP [0]);
  and _66267_ (_14627_, _09028_, \oc8051_golden_model_1.ACC [0]);
  and _66268_ (_14628_, _09030_, \oc8051_golden_model_1.B [0]);
  or _66269_ (_14629_, _14628_, _14627_);
  or _66270_ (_14630_, _14629_, _14626_);
  or _66271_ (_14631_, _14630_, _14625_);
  and _66272_ (_14632_, _09070_, \oc8051_golden_model_1.TH1 [0]);
  and _66273_ (_14633_, _09010_, \oc8051_golden_model_1.SP [0]);
  and _66274_ (_14634_, _09017_, \oc8051_golden_model_1.TL0 [0]);
  or _66275_ (_14635_, _14634_, _14633_);
  or _66276_ (_14636_, _14635_, _14632_);
  or _66277_ (_14637_, _14636_, _14631_);
  and _66278_ (_14638_, _09048_, \oc8051_golden_model_1.TH0 [0]);
  and _66279_ (_14639_, _09052_, \oc8051_golden_model_1.TL1 [0]);
  or _66280_ (_14640_, _14639_, _14638_);
  and _66281_ (_14641_, _09055_, \oc8051_golden_model_1.TCON [0]);
  and _66282_ (_14642_, _09059_, \oc8051_golden_model_1.PCON [0]);
  or _66283_ (_14643_, _14642_, _14641_);
  or _66284_ (_14644_, _14643_, _14640_);
  and _66285_ (_14645_, _09068_, \oc8051_golden_model_1.DPL [0]);
  and _66286_ (_14646_, _08993_, \oc8051_golden_model_1.P0INREG [0]);
  and _66287_ (_14647_, _08989_, \oc8051_golden_model_1.P2INREG [0]);
  and _66288_ (_14648_, _08998_, \oc8051_golden_model_1.P1INREG [0]);
  and _66289_ (_14649_, _09002_, \oc8051_golden_model_1.P3INREG [0]);
  or _66290_ (_14650_, _14649_, _14648_);
  or _66291_ (_14651_, _14650_, _14647_);
  or _66292_ (_14652_, _14651_, _14646_);
  or _66293_ (_14653_, _14652_, _14645_);
  and _66294_ (_14654_, _09035_, \oc8051_golden_model_1.SCON [0]);
  and _66295_ (_14655_, _09038_, \oc8051_golden_model_1.SBUF [0]);
  or _66296_ (_14656_, _14655_, _14654_);
  and _66297_ (_14657_, _09041_, \oc8051_golden_model_1.IE [0]);
  or _66298_ (_14658_, _14657_, _14656_);
  and _66299_ (_14659_, _09063_, \oc8051_golden_model_1.TMOD [0]);
  and _66300_ (_14660_, _09065_, \oc8051_golden_model_1.DPH [0]);
  or _66301_ (_14661_, _14660_, _14659_);
  or _66302_ (_14662_, _14661_, _14658_);
  or _66303_ (_14663_, _14662_, _14653_);
  or _66304_ (_14664_, _14663_, _14644_);
  or _66305_ (_14665_, _14664_, _14637_);
  or _66306_ (_14666_, _14665_, _14624_);
  and _66307_ (_14667_, _14666_, _08841_);
  or _66308_ (_14668_, _14667_, _08848_);
  or _66309_ (_14669_, _14668_, _14623_);
  and _66310_ (_14670_, _08848_, _06310_);
  nor _66311_ (_14671_, _14670_, _06279_);
  and _66312_ (_14672_, _14671_, _14669_);
  and _66313_ (_14673_, _09008_, _06279_);
  or _66314_ (_14674_, _14673_, _06275_);
  or _66315_ (_14675_, _14674_, _14672_);
  nor _66316_ (_14676_, _06009_, \oc8051_golden_model_1.PC [0]);
  nor _66317_ (_14677_, _14676_, _07335_);
  and _66318_ (_14678_, _14677_, _14675_);
  or _66319_ (_14679_, _14678_, _14567_);
  and _66320_ (_14680_, _14679_, _09086_);
  nor _66321_ (_14681_, _12623_, _09086_);
  or _66322_ (_14682_, _14681_, _14680_);
  and _66323_ (_14683_, _14682_, _09100_);
  and _66324_ (_14684_, _14564_, _07340_);
  or _66325_ (_14685_, _14684_, _14683_);
  and _66326_ (_14686_, _14685_, _07333_);
  and _66327_ (_14687_, _10577_, _07332_);
  or _66328_ (_14688_, _14687_, _07330_);
  or _66329_ (_14689_, _14688_, _14686_);
  nor _66330_ (_14690_, _06018_, \oc8051_golden_model_1.PC [0]);
  nor _66331_ (_14691_, _14690_, _09108_);
  and _66332_ (_14692_, _14691_, _14689_);
  and _66333_ (_14693_, _14563_, _09108_);
  or _66334_ (_14694_, _14693_, _09113_);
  or _66335_ (_14695_, _14694_, _14692_);
  and _66336_ (_14696_, _14695_, _14562_);
  or _66337_ (_14697_, _14696_, _07350_);
  or _66338_ (_14698_, _06016_, \oc8051_golden_model_1.PC [0]);
  and _66339_ (_14699_, _14698_, _09459_);
  and _66340_ (_14700_, _14699_, _14697_);
  nor _66341_ (_14701_, _09459_, _07250_);
  or _66342_ (_14702_, _14701_, _07360_);
  or _66343_ (_14703_, _14702_, _14700_);
  nand _66344_ (_14704_, _09447_, _07360_);
  and _66345_ (_14705_, _14704_, _14703_);
  or _66346_ (_14706_, _14705_, _07359_);
  nand _66347_ (_14707_, _08453_, _07359_);
  and _66348_ (_14708_, _14707_, _09534_);
  and _66349_ (_14709_, _14708_, _14706_);
  and _66350_ (_14710_, _06503_, _05701_);
  or _66351_ (_14711_, _14710_, _05998_);
  or _66352_ (_14712_, _14711_, _14709_);
  and _66353_ (_14713_, _14712_, _14561_);
  or _66354_ (_14714_, _14713_, _06272_);
  or _66355_ (_14715_, _14569_, _06273_);
  and _66356_ (_14716_, _14715_, _09473_);
  and _66357_ (_14717_, _14716_, _14714_);
  nor _66358_ (_14718_, _09473_, _07250_);
  nor _66359_ (_14719_, _14718_, _14717_);
  or _66360_ (_14720_, _14719_, _07055_);
  or _66361_ (_14721_, _09447_, _07375_);
  and _66362_ (_14722_, _14721_, _09495_);
  and _66363_ (_14723_, _14722_, _14720_);
  not _66364_ (_14724_, _14723_);
  and _66365_ (_14725_, _08453_, _07379_);
  nor _66366_ (_14726_, _14725_, _07632_);
  and _66367_ (_14727_, _14726_, _14724_);
  or _66368_ (_14728_, _14727_, _14560_);
  or _66369_ (_14729_, _14559_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _66370_ (_14730_, _09531_, _09526_);
  and _66371_ (_14731_, _14730_, _07387_);
  and _66372_ (_14732_, _14731_, _09525_);
  not _66373_ (_14733_, _14732_);
  and _66374_ (_14734_, _14733_, _14729_);
  and _66375_ (_14735_, _14734_, _14728_);
  and _66376_ (_14736_, _12412_, _06503_);
  not _66377_ (_14737_, _12234_);
  nor _66378_ (_14738_, _14737_, _06503_);
  or _66379_ (_14739_, _14738_, _14736_);
  and _66380_ (_14740_, _14739_, _09525_);
  and _66381_ (_14741_, _14740_, _14731_);
  or _66382_ (_41541_, _14741_, _14735_);
  nor _66383_ (_14742_, _09497_, _09448_);
  or _66384_ (_14743_, _14742_, _07375_);
  nor _66385_ (_14744_, _08784_, _08454_);
  nand _66386_ (_14745_, _14744_, _07359_);
  nand _66387_ (_14746_, _08403_, _07160_);
  nor _66388_ (_14747_, _08403_, _07160_);
  not _66389_ (_14748_, _14747_);
  and _66390_ (_14749_, _14748_, _14746_);
  and _66391_ (_14750_, _14749_, _07335_);
  or _66392_ (_14751_, _11310_, _06238_);
  nand _66393_ (_14752_, _14751_, _08401_);
  and _66394_ (_14753_, _14752_, _07309_);
  nor _66395_ (_14754_, _12902_, _07957_);
  or _66396_ (_14755_, _14754_, _08629_);
  nor _66397_ (_14756_, _14744_, _08782_);
  nor _66398_ (_14757_, _09483_, _08677_);
  nand _66399_ (_14758_, _14757_, _08687_);
  and _66400_ (_14759_, _06816_, _05667_);
  nor _66401_ (_14760_, _06816_, _06097_);
  or _66402_ (_14761_, _14760_, _14759_);
  nor _66403_ (_14762_, _14761_, _08687_);
  nor _66404_ (_14763_, _14762_, _07276_);
  and _66405_ (_14764_, _14763_, _14758_);
  or _66406_ (_14765_, _14764_, _07274_);
  or _66407_ (_14766_, _14765_, _14756_);
  nand _66408_ (_14767_, _12902_, _12880_);
  or _66409_ (_14768_, _14767_, _08670_);
  and _66410_ (_14769_, _14768_, _14766_);
  or _66411_ (_14770_, _14769_, _07692_);
  nor _66412_ (_14771_, _06052_, _05667_);
  nor _66413_ (_14772_, _14771_, _07284_);
  and _66414_ (_14773_, _14772_, _14770_);
  and _66415_ (_14774_, _09482_, _07284_);
  or _66416_ (_14775_, _14774_, _07294_);
  or _66417_ (_14776_, _14775_, _14773_);
  and _66418_ (_14777_, _14776_, _14755_);
  or _66419_ (_14778_, _14777_, _06351_);
  nand _66420_ (_14779_, _08403_, _06351_);
  and _66421_ (_14780_, _14779_, _06349_);
  and _66422_ (_14781_, _14780_, _14778_);
  not _66423_ (_14782_, _12903_);
  and _66424_ (_14783_, _14767_, _14782_);
  and _66425_ (_14784_, _14783_, _06348_);
  or _66426_ (_14785_, _14784_, _14781_);
  and _66427_ (_14786_, _14785_, _06049_);
  nor _66428_ (_14787_, _06049_, \oc8051_golden_model_1.PC [1]);
  or _66429_ (_14788_, _06441_, _14787_);
  or _66430_ (_14789_, _14788_, _14786_);
  nand _66431_ (_14790_, _08403_, _06441_);
  and _66432_ (_14791_, _14790_, _07310_);
  and _66433_ (_14792_, _14791_, _14789_);
  or _66434_ (_14793_, _14792_, _14753_);
  and _66435_ (_14794_, _14793_, _08821_);
  and _66436_ (_14795_, _07957_, \oc8051_golden_model_1.PSW [7]);
  or _66437_ (_14796_, _14795_, _14754_);
  and _66438_ (_14797_, _14796_, _07308_);
  or _66439_ (_14798_, _14797_, _06039_);
  or _66440_ (_14799_, _14798_, _14794_);
  and _66441_ (_14800_, _06039_, \oc8051_golden_model_1.PC [1]);
  nor _66442_ (_14801_, _14800_, _08832_);
  and _66443_ (_14802_, _14801_, _14799_);
  nor _66444_ (_14803_, _08836_, _07448_);
  or _66445_ (_14804_, _14803_, _08838_);
  or _66446_ (_14805_, _14804_, _14802_);
  or _66447_ (_14806_, _09402_, _08844_);
  and _66448_ (_14807_, _14806_, _08842_);
  and _66449_ (_14808_, _14807_, _14805_);
  nor _66450_ (_14809_, _08880_, _07448_);
  and _66451_ (_14810_, _09035_, \oc8051_golden_model_1.SCON [1]);
  and _66452_ (_14811_, _09038_, \oc8051_golden_model_1.SBUF [1]);
  or _66453_ (_14812_, _14811_, _14810_);
  and _66454_ (_14813_, _09041_, \oc8051_golden_model_1.IE [1]);
  or _66455_ (_14814_, _14813_, _14812_);
  and _66456_ (_14815_, _09023_, \oc8051_golden_model_1.PSW [1]);
  and _66457_ (_14816_, _09026_, \oc8051_golden_model_1.IP [1]);
  and _66458_ (_14817_, _09028_, \oc8051_golden_model_1.ACC [1]);
  and _66459_ (_14818_, _09030_, \oc8051_golden_model_1.B [1]);
  or _66460_ (_14819_, _14818_, _14817_);
  or _66461_ (_14820_, _14819_, _14816_);
  or _66462_ (_14821_, _14820_, _14815_);
  and _66463_ (_14822_, _09063_, \oc8051_golden_model_1.TMOD [1]);
  and _66464_ (_14823_, _09065_, \oc8051_golden_model_1.DPH [1]);
  or _66465_ (_14824_, _14823_, _14822_);
  or _66466_ (_14825_, _14824_, _14821_);
  or _66467_ (_14826_, _14825_, _14814_);
  and _66468_ (_14827_, _09070_, \oc8051_golden_model_1.TH1 [1]);
  and _66469_ (_14828_, _09010_, \oc8051_golden_model_1.SP [1]);
  and _66470_ (_14829_, _09017_, \oc8051_golden_model_1.TL0 [1]);
  or _66471_ (_14830_, _14829_, _14828_);
  or _66472_ (_14831_, _14830_, _14827_);
  and _66473_ (_14832_, _09048_, \oc8051_golden_model_1.TH0 [1]);
  and _66474_ (_14833_, _09052_, \oc8051_golden_model_1.TL1 [1]);
  or _66475_ (_14834_, _14833_, _14832_);
  and _66476_ (_14835_, _09055_, \oc8051_golden_model_1.TCON [1]);
  and _66477_ (_14836_, _09059_, \oc8051_golden_model_1.PCON [1]);
  or _66478_ (_14837_, _14836_, _14835_);
  or _66479_ (_14838_, _14837_, _14834_);
  and _66480_ (_14839_, _09068_, \oc8051_golden_model_1.DPL [1]);
  and _66481_ (_14840_, _08989_, \oc8051_golden_model_1.P2INREG [1]);
  and _66482_ (_14841_, _08993_, \oc8051_golden_model_1.P0INREG [1]);
  and _66483_ (_14842_, _08998_, \oc8051_golden_model_1.P1INREG [1]);
  and _66484_ (_14843_, _09002_, \oc8051_golden_model_1.P3INREG [1]);
  or _66485_ (_14844_, _14843_, _14842_);
  or _66486_ (_14845_, _14844_, _14841_);
  or _66487_ (_14846_, _14845_, _14840_);
  or _66488_ (_14847_, _14846_, _14839_);
  or _66489_ (_14848_, _14847_, _14838_);
  or _66490_ (_14849_, _14848_, _14831_);
  or _66491_ (_14850_, _14849_, _14826_);
  or _66492_ (_14851_, _14850_, _14809_);
  and _66493_ (_14852_, _14851_, _08841_);
  or _66494_ (_14853_, _14852_, _08848_);
  or _66495_ (_14854_, _14853_, _14808_);
  and _66496_ (_14855_, _08848_, _07127_);
  nor _66497_ (_14856_, _14855_, _06279_);
  and _66498_ (_14857_, _14856_, _14854_);
  and _66499_ (_14858_, _09012_, _06279_);
  or _66500_ (_14859_, _14858_, _06275_);
  or _66501_ (_14860_, _14859_, _14857_);
  nor _66502_ (_14861_, _06009_, _05667_);
  nor _66503_ (_14862_, _14861_, _07335_);
  and _66504_ (_14863_, _14862_, _14860_);
  or _66505_ (_14864_, _14863_, _14750_);
  and _66506_ (_14865_, _14864_, _09086_);
  and _66507_ (_14866_, _10579_, _07338_);
  or _66508_ (_14867_, _14866_, _14865_);
  and _66509_ (_14868_, _14867_, _09100_);
  and _66510_ (_14869_, _14747_, _07340_);
  or _66511_ (_14870_, _14869_, _14868_);
  and _66512_ (_14871_, _14870_, _07333_);
  and _66513_ (_14872_, _10576_, _07332_);
  or _66514_ (_14873_, _14872_, _07330_);
  or _66515_ (_14874_, _14873_, _14871_);
  nor _66516_ (_14875_, _06018_, _05667_);
  nor _66517_ (_14876_, _14875_, _09108_);
  and _66518_ (_14877_, _14876_, _14874_);
  and _66519_ (_14878_, _14746_, _09108_);
  or _66520_ (_14879_, _14878_, _09113_);
  or _66521_ (_14880_, _14879_, _14877_);
  nand _66522_ (_14881_, _10578_, _09113_);
  and _66523_ (_14882_, _14881_, _06016_);
  and _66524_ (_14883_, _14882_, _14880_);
  nor _66525_ (_14884_, _06016_, \oc8051_golden_model_1.PC [1]);
  or _66526_ (_14885_, _07588_, _14884_);
  or _66527_ (_14886_, _14885_, _14883_);
  and _66528_ (_14887_, _14757_, _07588_);
  nor _66529_ (_14888_, _14887_, _07177_);
  and _66530_ (_14889_, _14888_, _14886_);
  not _66531_ (_14890_, _07924_);
  and _66532_ (_14891_, _14757_, _05921_);
  nor _66533_ (_14892_, _14891_, _14890_);
  or _66534_ (_14893_, _14892_, _14889_);
  nand _66535_ (_14894_, _14757_, _07521_);
  and _66536_ (_14895_, _14894_, _07361_);
  and _66537_ (_14896_, _14895_, _14893_);
  nor _66538_ (_14897_, _14742_, _07361_);
  or _66539_ (_14898_, _14897_, _07359_);
  or _66540_ (_14899_, _14898_, _14896_);
  and _66541_ (_14900_, _14899_, _14745_);
  or _66542_ (_14901_, _14900_, _06503_);
  nand _66543_ (_14902_, _06503_, _12444_);
  and _66544_ (_14903_, _14902_, _13082_);
  and _66545_ (_14904_, _14903_, _14901_);
  and _66546_ (_14905_, _05998_, _05667_);
  or _66547_ (_14906_, _06272_, _14905_);
  or _66548_ (_14907_, _14906_, _14904_);
  and _66549_ (_14908_, _06785_, _05996_);
  nor _66550_ (_14909_, _14754_, _06273_);
  nor _66551_ (_14910_, _14909_, _14908_);
  and _66552_ (_14911_, _14910_, _14907_);
  and _66553_ (_14912_, _14757_, _07581_);
  nor _66554_ (_14913_, _14912_, _14911_);
  nor _66555_ (_14914_, _14913_, _07534_);
  and _66556_ (_14915_, _06323_, _05996_);
  and _66557_ (_14916_, _14757_, _07534_);
  or _66558_ (_14917_, _14916_, _14915_);
  or _66559_ (_14918_, _14917_, _14914_);
  not _66560_ (_14919_, _07591_);
  or _66561_ (_14920_, _14891_, _14919_);
  and _66562_ (_14921_, _14920_, _14918_);
  and _66563_ (_14922_, _14757_, _07535_);
  or _66564_ (_14923_, _14922_, _07055_);
  or _66565_ (_14924_, _14923_, _14921_);
  and _66566_ (_14925_, _14924_, _14743_);
  or _66567_ (_14926_, _14925_, _07379_);
  or _66568_ (_14927_, _14744_, _09495_);
  and _66569_ (_14928_, _14927_, _07631_);
  and _66570_ (_14929_, _14928_, _14926_);
  or _66571_ (_14930_, _14929_, _14560_);
  or _66572_ (_14931_, _14559_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _66573_ (_14932_, _14931_, _14733_);
  and _66574_ (_14933_, _14932_, _14930_);
  not _66575_ (_14934_, _12230_);
  nor _66576_ (_14935_, _14934_, _06503_);
  and _66577_ (_14936_, _12407_, _06503_);
  or _66578_ (_14937_, _14936_, _14935_);
  and _66579_ (_14938_, _14937_, _09525_);
  and _66580_ (_14939_, _14938_, _14731_);
  or _66581_ (_41542_, _14939_, _14933_);
  or _66582_ (_14940_, _09483_, _09481_);
  nor _66583_ (_14941_, _09484_, _09473_);
  and _66584_ (_14942_, _14941_, _14940_);
  nand _66585_ (_14943_, _06329_, _05848_);
  nor _66586_ (_14944_, _06113_, _06016_);
  nand _66587_ (_14945_, _08502_, _06769_);
  nor _66588_ (_14946_, _08502_, _06769_);
  not _66589_ (_14947_, _14946_);
  and _66590_ (_14948_, _14947_, _14945_);
  and _66591_ (_14949_, _14948_, _07335_);
  nand _66592_ (_14950_, _09356_, _06366_);
  nand _66593_ (_14951_, _14950_, _08500_);
  and _66594_ (_14952_, _14951_, _07309_);
  nor _66595_ (_14953_, _12878_, _08000_);
  or _66596_ (_14954_, _14953_, _08629_);
  nand _66597_ (_14955_, _12878_, _12855_);
  or _66598_ (_14956_, _14955_, _08670_);
  and _66599_ (_14957_, _08784_, _08502_);
  nor _66600_ (_14958_, _08784_, _08502_);
  or _66601_ (_14959_, _14958_, _14957_);
  and _66602_ (_14960_, _14959_, _07276_);
  and _66603_ (_14961_, _08677_, _07854_);
  nor _66604_ (_14962_, _08677_, _07854_);
  or _66605_ (_14963_, _14962_, _14961_);
  or _66606_ (_14964_, _14963_, _08685_);
  and _66607_ (_14965_, _06816_, _06111_);
  nor _66608_ (_14966_, _06816_, _10280_);
  or _66609_ (_14967_, _14966_, _14965_);
  nor _66610_ (_14968_, _14967_, _08687_);
  nor _66611_ (_14969_, _14968_, _07276_);
  and _66612_ (_14970_, _14969_, _14964_);
  or _66613_ (_14971_, _14970_, _07274_);
  or _66614_ (_14972_, _14971_, _14960_);
  and _66615_ (_14973_, _14972_, _14956_);
  or _66616_ (_14974_, _14973_, _07692_);
  nor _66617_ (_14975_, _06111_, _06052_);
  nor _66618_ (_14976_, _14975_, _07284_);
  and _66619_ (_14977_, _14976_, _14974_);
  and _66620_ (_14978_, _09481_, _07284_);
  or _66621_ (_14979_, _14978_, _07294_);
  or _66622_ (_14980_, _14979_, _14977_);
  and _66623_ (_14981_, _14980_, _14954_);
  or _66624_ (_14982_, _14981_, _06351_);
  nand _66625_ (_14983_, _08502_, _06351_);
  and _66626_ (_14984_, _14983_, _06349_);
  and _66627_ (_14985_, _14984_, _14982_);
  not _66628_ (_14986_, _12879_);
  and _66629_ (_14987_, _14955_, _14986_);
  and _66630_ (_14988_, _14987_, _06348_);
  or _66631_ (_14989_, _14988_, _14985_);
  and _66632_ (_14990_, _14989_, _06049_);
  nor _66633_ (_14991_, _06113_, _06049_);
  or _66634_ (_14992_, _06441_, _14991_);
  or _66635_ (_14993_, _14992_, _14990_);
  nand _66636_ (_14994_, _08502_, _06441_);
  and _66637_ (_14995_, _14994_, _07310_);
  and _66638_ (_14996_, _14995_, _14993_);
  or _66639_ (_14997_, _14996_, _14952_);
  and _66640_ (_14998_, _14997_, _08821_);
  and _66641_ (_14999_, _08000_, \oc8051_golden_model_1.PSW [7]);
  or _66642_ (_15000_, _14999_, _14953_);
  and _66643_ (_15001_, _15000_, _07308_);
  or _66644_ (_15002_, _15001_, _06039_);
  or _66645_ (_15003_, _15002_, _14998_);
  and _66646_ (_15004_, _06113_, _06039_);
  nor _66647_ (_15005_, _15004_, _08832_);
  and _66648_ (_15006_, _15005_, _15003_);
  nor _66649_ (_15007_, _08836_, _07854_);
  or _66650_ (_15008_, _15007_, _08838_);
  or _66651_ (_15009_, _15008_, _15006_);
  not _66652_ (_15010_, _08838_);
  or _66653_ (_15011_, _09356_, _15010_);
  and _66654_ (_15012_, _15011_, _08842_);
  and _66655_ (_15013_, _15012_, _15009_);
  nor _66656_ (_15014_, _08880_, _07854_);
  and _66657_ (_15015_, _08989_, \oc8051_golden_model_1.P2INREG [2]);
  and _66658_ (_15016_, _08993_, \oc8051_golden_model_1.P0INREG [2]);
  and _66659_ (_15017_, _08998_, \oc8051_golden_model_1.P1INREG [2]);
  and _66660_ (_15018_, _09002_, \oc8051_golden_model_1.P3INREG [2]);
  or _66661_ (_15019_, _15018_, _15017_);
  or _66662_ (_15020_, _15019_, _15016_);
  or _66663_ (_15021_, _15020_, _15015_);
  and _66664_ (_15022_, _09010_, \oc8051_golden_model_1.SP [2]);
  and _66665_ (_15023_, _09017_, \oc8051_golden_model_1.TL0 [2]);
  or _66666_ (_15024_, _15023_, _15022_);
  or _66667_ (_15025_, _15024_, _15021_);
  and _66668_ (_15026_, _09023_, \oc8051_golden_model_1.PSW [2]);
  and _66669_ (_15027_, _09026_, \oc8051_golden_model_1.IP [2]);
  and _66670_ (_15028_, _09028_, \oc8051_golden_model_1.ACC [2]);
  and _66671_ (_15029_, _09030_, \oc8051_golden_model_1.B [2]);
  or _66672_ (_15030_, _15029_, _15028_);
  or _66673_ (_15031_, _15030_, _15027_);
  or _66674_ (_15032_, _15031_, _15026_);
  and _66675_ (_15033_, _09035_, \oc8051_golden_model_1.SCON [2]);
  and _66676_ (_15034_, _09038_, \oc8051_golden_model_1.SBUF [2]);
  or _66677_ (_15035_, _15034_, _15033_);
  and _66678_ (_15036_, _09041_, \oc8051_golden_model_1.IE [2]);
  or _66679_ (_15037_, _15036_, _15035_);
  or _66680_ (_15038_, _15037_, _15032_);
  or _66681_ (_15039_, _15038_, _15025_);
  and _66682_ (_15040_, _09048_, \oc8051_golden_model_1.TH0 [2]);
  and _66683_ (_15041_, _09052_, \oc8051_golden_model_1.TL1 [2]);
  or _66684_ (_15042_, _15041_, _15040_);
  and _66685_ (_15043_, _09055_, \oc8051_golden_model_1.TCON [2]);
  and _66686_ (_15044_, _09059_, \oc8051_golden_model_1.PCON [2]);
  or _66687_ (_15045_, _15044_, _15043_);
  or _66688_ (_15046_, _15045_, _15042_);
  and _66689_ (_15047_, _09063_, \oc8051_golden_model_1.TMOD [2]);
  and _66690_ (_15048_, _09065_, \oc8051_golden_model_1.DPH [2]);
  or _66691_ (_15049_, _15048_, _15047_);
  and _66692_ (_15050_, _09068_, \oc8051_golden_model_1.DPL [2]);
  and _66693_ (_15051_, _09070_, \oc8051_golden_model_1.TH1 [2]);
  or _66694_ (_15052_, _15051_, _15050_);
  or _66695_ (_15053_, _15052_, _15049_);
  or _66696_ (_15054_, _15053_, _15046_);
  or _66697_ (_15055_, _15054_, _15039_);
  or _66698_ (_15056_, _15055_, _15014_);
  and _66699_ (_15057_, _15056_, _08841_);
  or _66700_ (_15058_, _15057_, _08848_);
  or _66701_ (_15059_, _15058_, _15013_);
  and _66702_ (_15060_, _08848_, _06727_);
  nor _66703_ (_15061_, _15060_, _06279_);
  and _66704_ (_15062_, _15061_, _15059_);
  and _66705_ (_15063_, _09057_, _06279_);
  or _66706_ (_15064_, _15063_, _06275_);
  or _66707_ (_15065_, _15064_, _15062_);
  nor _66708_ (_15066_, _06111_, _06009_);
  nor _66709_ (_15067_, _15066_, _07335_);
  and _66710_ (_15068_, _15067_, _15065_);
  or _66711_ (_15069_, _15068_, _14949_);
  and _66712_ (_15070_, _15069_, _09086_);
  and _66713_ (_15071_, _10583_, _07338_);
  or _66714_ (_15072_, _15071_, _15070_);
  and _66715_ (_15073_, _15072_, _09100_);
  and _66716_ (_15074_, _14946_, _07340_);
  or _66717_ (_15075_, _15074_, _15073_);
  and _66718_ (_15076_, _15075_, _07333_);
  and _66719_ (_15077_, _10575_, _07332_);
  or _66720_ (_15078_, _15077_, _07330_);
  or _66721_ (_15079_, _15078_, _15076_);
  nor _66722_ (_15080_, _06111_, _06018_);
  nor _66723_ (_15081_, _15080_, _09108_);
  and _66724_ (_15082_, _15081_, _15079_);
  and _66725_ (_15083_, _14945_, _09108_);
  or _66726_ (_15084_, _15083_, _09113_);
  or _66727_ (_15085_, _15084_, _15082_);
  nand _66728_ (_15086_, _10582_, _09113_);
  and _66729_ (_15087_, _15086_, _06016_);
  and _66730_ (_15088_, _15087_, _15085_);
  or _66731_ (_15089_, _15088_, _14944_);
  and _66732_ (_15090_, _15089_, _09122_);
  not _66733_ (_15091_, _09122_);
  and _66734_ (_15092_, _14963_, _15091_);
  or _66735_ (_15093_, _15092_, _07521_);
  or _66736_ (_15094_, _15093_, _15090_);
  and _66737_ (_15095_, _06331_, _05848_);
  not _66738_ (_15096_, _15095_);
  not _66739_ (_15097_, _07521_);
  or _66740_ (_15098_, _14963_, _15097_);
  and _66741_ (_15099_, _15098_, _15096_);
  nand _66742_ (_15100_, _15099_, _15094_);
  nor _66743_ (_15101_, _09448_, _09357_);
  nor _66744_ (_15102_, _15101_, _09449_);
  or _66745_ (_15103_, _15102_, _15096_);
  nand _66746_ (_15104_, _15103_, _15100_);
  and _66747_ (_15105_, _15104_, _14943_);
  nor _66748_ (_15106_, _15102_, _14943_);
  or _66749_ (_15107_, _15106_, _15105_);
  and _66750_ (_15108_, _15107_, _09458_);
  and _66751_ (_15109_, _14959_, _07359_);
  or _66752_ (_15110_, _15109_, _06503_);
  or _66753_ (_15111_, _15110_, _15108_);
  nand _66754_ (_15112_, _12442_, _06503_);
  and _66755_ (_15113_, _15112_, _13082_);
  and _66756_ (_15114_, _15113_, _15111_);
  and _66757_ (_15115_, _06111_, _05998_);
  or _66758_ (_15116_, _06272_, _15115_);
  or _66759_ (_15117_, _15116_, _15114_);
  or _66760_ (_15118_, _14953_, _06273_);
  and _66761_ (_15119_, _15118_, _09473_);
  and _66762_ (_15120_, _15119_, _15117_);
  or _66763_ (_15121_, _15120_, _14942_);
  and _66764_ (_15122_, _15121_, _07375_);
  or _66765_ (_15123_, _09497_, _09356_);
  nor _66766_ (_15124_, _09498_, _07375_);
  and _66767_ (_15125_, _15124_, _15123_);
  or _66768_ (_15126_, _15125_, _07379_);
  or _66769_ (_15127_, _15126_, _15122_);
  nor _66770_ (_15128_, _08503_, _08454_);
  nor _66771_ (_15129_, _15128_, _08504_);
  or _66772_ (_15130_, _15129_, _09495_);
  and _66773_ (_15131_, _15130_, _07631_);
  and _66774_ (_15132_, _15131_, _15127_);
  or _66775_ (_15133_, _15132_, _14560_);
  or _66776_ (_15134_, _14559_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _66777_ (_15135_, _15134_, _14733_);
  and _66778_ (_15136_, _15135_, _15133_);
  and _66779_ (_15137_, _12400_, _06503_);
  and _66780_ (_15138_, _12224_, _09534_);
  or _66781_ (_15139_, _15138_, _15137_);
  and _66782_ (_15140_, _15139_, _09525_);
  and _66783_ (_15141_, _15140_, _14731_);
  or _66784_ (_41543_, _15141_, _15136_);
  nor _66785_ (_15142_, _09449_, _09311_);
  or _66786_ (_15143_, _15142_, _09450_);
  and _66787_ (_15144_, _15143_, _07360_);
  nor _66788_ (_15145_, _06521_, _06016_);
  or _66789_ (_15146_, _06150_, _06009_);
  nand _66790_ (_15147_, _08832_, _07680_);
  nor _66791_ (_15148_, _13007_, _07994_);
  or _66792_ (_15149_, _15148_, _08629_);
  nand _66793_ (_15150_, _13007_, _12984_);
  or _66794_ (_15151_, _15150_, _08670_);
  nor _66795_ (_15152_, _14957_, _08358_);
  or _66796_ (_15153_, _15152_, _08786_);
  and _66797_ (_15154_, _15153_, _07276_);
  nor _66798_ (_15155_, _14961_, _07680_);
  or _66799_ (_15156_, _15155_, _08678_);
  or _66800_ (_15157_, _15156_, _08685_);
  and _66801_ (_15158_, _06816_, _06150_);
  nor _66802_ (_15159_, _06816_, _10334_);
  or _66803_ (_15160_, _15159_, _15158_);
  nor _66804_ (_15161_, _15160_, _08687_);
  nor _66805_ (_15162_, _15161_, _07276_);
  and _66806_ (_15163_, _15162_, _15157_);
  or _66807_ (_15164_, _15163_, _07274_);
  or _66808_ (_15165_, _15164_, _15154_);
  and _66809_ (_15166_, _15165_, _15151_);
  or _66810_ (_15167_, _15166_, _07692_);
  nor _66811_ (_15168_, _06150_, _06052_);
  nor _66812_ (_15169_, _15168_, _07284_);
  and _66813_ (_15170_, _15169_, _15167_);
  and _66814_ (_15171_, _09480_, _07284_);
  or _66815_ (_15172_, _15171_, _07294_);
  or _66816_ (_15173_, _15172_, _15170_);
  and _66817_ (_15174_, _15173_, _15149_);
  or _66818_ (_15175_, _15174_, _06351_);
  nand _66819_ (_15176_, _08358_, _06351_);
  and _66820_ (_15178_, _15176_, _06349_);
  and _66821_ (_15179_, _15178_, _15175_);
  not _66822_ (_15180_, _13008_);
  and _66823_ (_15181_, _15150_, _15180_);
  and _66824_ (_15182_, _15181_, _06348_);
  or _66825_ (_15183_, _15182_, _15179_);
  and _66826_ (_15184_, _15183_, _06049_);
  nor _66827_ (_15185_, _06521_, _06049_);
  or _66828_ (_15186_, _06441_, _15185_);
  or _66829_ (_15187_, _15186_, _15184_);
  nand _66830_ (_15188_, _08358_, _06441_);
  and _66831_ (_15189_, _15188_, _15187_);
  or _66832_ (_15190_, _15189_, _07309_);
  and _66833_ (_15191_, _09310_, _06366_);
  nand _66834_ (_15192_, _08356_, _07309_);
  or _66835_ (_15193_, _15192_, _15191_);
  and _66836_ (_15194_, _15193_, _15190_);
  or _66837_ (_15195_, _15194_, _07308_);
  and _66838_ (_15196_, _07994_, \oc8051_golden_model_1.PSW [7]);
  or _66839_ (_15197_, _15148_, _15196_);
  or _66840_ (_15198_, _15197_, _08821_);
  and _66841_ (_15199_, _15198_, _07745_);
  and _66842_ (_15200_, _15199_, _15195_);
  and _66843_ (_15201_, _06150_, _06039_);
  or _66844_ (_15202_, _08832_, _15201_);
  or _66845_ (_15203_, _15202_, _15200_);
  and _66846_ (_15204_, _15203_, _15147_);
  or _66847_ (_15205_, _15204_, _08838_);
  or _66848_ (_15206_, _09310_, _15010_);
  and _66849_ (_15207_, _15206_, _08842_);
  and _66850_ (_15208_, _15207_, _15205_);
  nor _66851_ (_15209_, _08880_, _07680_);
  and _66852_ (_15210_, _08989_, \oc8051_golden_model_1.P2INREG [3]);
  and _66853_ (_15211_, _08993_, \oc8051_golden_model_1.P0INREG [3]);
  and _66854_ (_15212_, _08998_, \oc8051_golden_model_1.P1INREG [3]);
  and _66855_ (_15213_, _09002_, \oc8051_golden_model_1.P3INREG [3]);
  or _66856_ (_15214_, _15213_, _15212_);
  or _66857_ (_15215_, _15214_, _15211_);
  or _66858_ (_15216_, _15215_, _15210_);
  and _66859_ (_15217_, _09010_, \oc8051_golden_model_1.SP [3]);
  and _66860_ (_15218_, _09017_, \oc8051_golden_model_1.TL0 [3]);
  or _66861_ (_15219_, _15218_, _15217_);
  or _66862_ (_15220_, _15219_, _15216_);
  and _66863_ (_15221_, _09023_, \oc8051_golden_model_1.PSW [3]);
  and _66864_ (_15222_, _09026_, \oc8051_golden_model_1.IP [3]);
  and _66865_ (_15223_, _09028_, \oc8051_golden_model_1.ACC [3]);
  and _66866_ (_15224_, _09030_, \oc8051_golden_model_1.B [3]);
  or _66867_ (_15225_, _15224_, _15223_);
  or _66868_ (_15226_, _15225_, _15222_);
  or _66869_ (_15227_, _15226_, _15221_);
  and _66870_ (_15228_, _09035_, \oc8051_golden_model_1.SCON [3]);
  and _66871_ (_15229_, _09038_, \oc8051_golden_model_1.SBUF [3]);
  or _66872_ (_15230_, _15229_, _15228_);
  and _66873_ (_15231_, _09041_, \oc8051_golden_model_1.IE [3]);
  or _66874_ (_15232_, _15231_, _15230_);
  or _66875_ (_15233_, _15232_, _15227_);
  or _66876_ (_15234_, _15233_, _15220_);
  and _66877_ (_15235_, _09048_, \oc8051_golden_model_1.TH0 [3]);
  and _66878_ (_15236_, _09052_, \oc8051_golden_model_1.TL1 [3]);
  or _66879_ (_15237_, _15236_, _15235_);
  and _66880_ (_15238_, _09055_, \oc8051_golden_model_1.TCON [3]);
  and _66881_ (_15239_, _09059_, \oc8051_golden_model_1.PCON [3]);
  or _66882_ (_15240_, _15239_, _15238_);
  or _66883_ (_15241_, _15240_, _15237_);
  and _66884_ (_15242_, _09063_, \oc8051_golden_model_1.TMOD [3]);
  and _66885_ (_15243_, _09065_, \oc8051_golden_model_1.DPH [3]);
  or _66886_ (_15244_, _15243_, _15242_);
  and _66887_ (_15245_, _09068_, \oc8051_golden_model_1.DPL [3]);
  and _66888_ (_15246_, _09070_, \oc8051_golden_model_1.TH1 [3]);
  or _66889_ (_15247_, _15246_, _15245_);
  or _66890_ (_15248_, _15247_, _15244_);
  or _66891_ (_15249_, _15248_, _15241_);
  or _66892_ (_15250_, _15249_, _15234_);
  or _66893_ (_15251_, _15250_, _15209_);
  and _66894_ (_15252_, _15251_, _08841_);
  or _66895_ (_15253_, _15252_, _08848_);
  or _66896_ (_15254_, _15253_, _15208_);
  and _66897_ (_15255_, _08848_, _06269_);
  nor _66898_ (_15256_, _15255_, _06279_);
  and _66899_ (_15257_, _15256_, _15254_);
  and _66900_ (_15258_, _09014_, _06279_);
  or _66901_ (_15259_, _15258_, _06275_);
  or _66902_ (_15260_, _15259_, _15257_);
  and _66903_ (_15261_, _15260_, _15146_);
  or _66904_ (_15262_, _15261_, _07335_);
  nand _66905_ (_15263_, _08358_, _06595_);
  nor _66906_ (_15264_, _08358_, _06595_);
  not _66907_ (_15265_, _15264_);
  and _66908_ (_15266_, _15265_, _15263_);
  or _66909_ (_15267_, _15266_, _07336_);
  and _66910_ (_15268_, _15267_, _09086_);
  and _66911_ (_15269_, _15268_, _15262_);
  nor _66912_ (_15270_, _12619_, _07340_);
  nor _66913_ (_15271_, _15270_, _07341_);
  or _66914_ (_15272_, _15271_, _15269_);
  or _66915_ (_15273_, _15264_, _09100_);
  and _66916_ (_15274_, _15273_, _07333_);
  and _66917_ (_15275_, _15274_, _15272_);
  and _66918_ (_15276_, _10573_, _07332_);
  or _66919_ (_15277_, _15276_, _07330_);
  or _66920_ (_15278_, _15277_, _15275_);
  nor _66921_ (_15279_, _06150_, _06018_);
  nor _66922_ (_15280_, _15279_, _09108_);
  and _66923_ (_15281_, _15280_, _15278_);
  and _66924_ (_15282_, _15263_, _09108_);
  or _66925_ (_15283_, _15282_, _09113_);
  or _66926_ (_15284_, _15283_, _15281_);
  nand _66927_ (_15285_, _10574_, _09113_);
  and _66928_ (_15286_, _15285_, _06016_);
  and _66929_ (_15287_, _15286_, _15284_);
  or _66930_ (_15288_, _15287_, _15145_);
  and _66931_ (_15289_, _15288_, _09122_);
  and _66932_ (_15290_, _15156_, _15091_);
  or _66933_ (_15291_, _15290_, _07521_);
  or _66934_ (_15292_, _15291_, _15289_);
  or _66935_ (_15293_, _15156_, _15097_);
  and _66936_ (_15294_, _15293_, _07361_);
  and _66937_ (_15295_, _15294_, _15292_);
  or _66938_ (_15296_, _15295_, _15144_);
  and _66939_ (_15297_, _15296_, _09458_);
  and _66940_ (_15298_, _15153_, _07359_);
  or _66941_ (_15299_, _15298_, _06503_);
  or _66942_ (_15300_, _15299_, _15297_);
  nand _66943_ (_15301_, _12437_, _06503_);
  and _66944_ (_15302_, _15301_, _13082_);
  and _66945_ (_15303_, _15302_, _15300_);
  and _66946_ (_15304_, _06150_, _05998_);
  or _66947_ (_15305_, _06272_, _15304_);
  or _66948_ (_15306_, _15305_, _15303_);
  or _66949_ (_15307_, _15148_, _06273_);
  and _66950_ (_15308_, _15307_, _09473_);
  and _66951_ (_15309_, _15308_, _15306_);
  nor _66952_ (_15310_, _09484_, _09480_);
  nor _66953_ (_15311_, _15310_, _09485_);
  and _66954_ (_15312_, _15311_, _09474_);
  or _66955_ (_15313_, _15312_, _07055_);
  or _66956_ (_15314_, _15313_, _15309_);
  nor _66957_ (_15315_, _09498_, _09310_);
  nor _66958_ (_15316_, _15315_, _09499_);
  or _66959_ (_15317_, _15316_, _07375_);
  and _66960_ (_15318_, _15317_, _15314_);
  or _66961_ (_15319_, _15318_, _07379_);
  nor _66962_ (_15320_, _08504_, _08359_);
  nor _66963_ (_15321_, _15320_, _08505_);
  or _66964_ (_15322_, _15321_, _09495_);
  and _66965_ (_15323_, _15322_, _07631_);
  and _66966_ (_15324_, _15323_, _15319_);
  or _66967_ (_15325_, _15324_, _14560_);
  or _66968_ (_15326_, _14559_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _66969_ (_15327_, _15326_, _14733_);
  and _66970_ (_15328_, _15327_, _15325_);
  not _66971_ (_15329_, _12220_);
  nor _66972_ (_15330_, _15329_, _06503_);
  and _66973_ (_15331_, _12395_, _06503_);
  or _66974_ (_15332_, _15331_, _15330_);
  and _66975_ (_15333_, _15332_, _09525_);
  and _66976_ (_15334_, _15333_, _14731_);
  or _66977_ (_41545_, _15334_, _15328_);
  nor _66978_ (_15335_, _09499_, _09264_);
  nor _66979_ (_15336_, _15335_, _09500_);
  or _66980_ (_15337_, _15336_, _07375_);
  and _66981_ (_15338_, _08678_, _08596_);
  nor _66982_ (_15339_, _08678_, _08596_);
  nor _66983_ (_15340_, _15339_, _15338_);
  nand _66984_ (_15341_, _15340_, _15091_);
  nand _66985_ (_15342_, _08986_, _08598_);
  nor _66986_ (_15343_, _08986_, _08598_);
  not _66987_ (_15344_, _15343_);
  and _66988_ (_15345_, _15344_, _15342_);
  and _66989_ (_15346_, _15345_, _07335_);
  nand _66990_ (_15347_, _08832_, _08596_);
  nor _66991_ (_15348_, _12928_, _12927_);
  and _66992_ (_15349_, _12928_, \oc8051_golden_model_1.PSW [7]);
  or _66993_ (_15350_, _15349_, _15348_);
  and _66994_ (_15351_, _15350_, _07308_);
  or _66995_ (_15352_, _15348_, _08629_);
  nand _66996_ (_15353_, _12929_, _12927_);
  or _66997_ (_15354_, _15353_, _08670_);
  nand _66998_ (_15355_, _15340_, _08687_);
  and _66999_ (_15356_, _12253_, _06816_);
  or _67000_ (_15357_, _06816_, _10204_);
  nand _67001_ (_15358_, _15357_, _08685_);
  or _67002_ (_15359_, _15358_, _15356_);
  and _67003_ (_15360_, _15359_, _15355_);
  or _67004_ (_15361_, _15360_, _07269_);
  or _67005_ (_15362_, _09264_, _07270_);
  and _67006_ (_15363_, _15362_, _15361_);
  or _67007_ (_15364_, _15363_, _07276_);
  and _67008_ (_15365_, _08786_, _08598_);
  nor _67009_ (_15366_, _08786_, _08598_);
  or _67010_ (_15367_, _15366_, _15365_);
  or _67011_ (_15368_, _15367_, _08782_);
  and _67012_ (_15369_, _15368_, _15364_);
  or _67013_ (_15370_, _15369_, _07274_);
  and _67014_ (_15371_, _15370_, _15354_);
  or _67015_ (_15372_, _15371_, _07692_);
  nor _67016_ (_15373_, _12253_, _06052_);
  nor _67017_ (_15374_, _15373_, _07284_);
  and _67018_ (_15375_, _15374_, _15372_);
  and _67019_ (_15376_, _09479_, _07284_);
  or _67020_ (_15377_, _15376_, _07294_);
  or _67021_ (_15378_, _15377_, _15375_);
  and _67022_ (_15379_, _15378_, _15352_);
  or _67023_ (_15380_, _15379_, _06351_);
  nand _67024_ (_15381_, _08598_, _06351_);
  and _67025_ (_15382_, _15381_, _06349_);
  and _67026_ (_15383_, _15382_, _15380_);
  not _67027_ (_15384_, _12930_);
  and _67028_ (_15385_, _15353_, _15384_);
  and _67029_ (_15386_, _15385_, _06348_);
  or _67030_ (_15387_, _15386_, _15383_);
  and _67031_ (_15388_, _15387_, _06049_);
  nor _67032_ (_15389_, _12254_, _06049_);
  or _67033_ (_15390_, _15389_, _06441_);
  or _67034_ (_15391_, _15390_, _15388_);
  nand _67035_ (_15392_, _08598_, _06441_);
  and _67036_ (_15393_, _15392_, _15391_);
  or _67037_ (_15394_, _15393_, _07309_);
  and _67038_ (_15395_, _09264_, _06366_);
  nand _67039_ (_15396_, _08551_, _07309_);
  or _67040_ (_15397_, _15396_, _15395_);
  and _67041_ (_15398_, _15397_, _08821_);
  and _67042_ (_15399_, _15398_, _15394_);
  or _67043_ (_15400_, _15399_, _15351_);
  and _67044_ (_15401_, _15400_, _07745_);
  and _67045_ (_15402_, _12253_, _06039_);
  or _67046_ (_15403_, _15402_, _08832_);
  or _67047_ (_15404_, _15403_, _15401_);
  and _67048_ (_15405_, _15404_, _15347_);
  or _67049_ (_15406_, _15405_, _08838_);
  or _67050_ (_15407_, _09264_, _15010_);
  and _67051_ (_15408_, _15407_, _08842_);
  and _67052_ (_15409_, _15408_, _15406_);
  nor _67053_ (_15410_, _08880_, _08596_);
  and _67054_ (_15411_, _08989_, \oc8051_golden_model_1.P2INREG [4]);
  and _67055_ (_15412_, _08993_, \oc8051_golden_model_1.P0INREG [4]);
  and _67056_ (_15413_, _08998_, \oc8051_golden_model_1.P1INREG [4]);
  and _67057_ (_15414_, _09002_, \oc8051_golden_model_1.P3INREG [4]);
  or _67058_ (_15415_, _15414_, _15413_);
  or _67059_ (_15416_, _15415_, _15412_);
  or _67060_ (_15417_, _15416_, _15411_);
  and _67061_ (_15418_, _09010_, \oc8051_golden_model_1.SP [4]);
  and _67062_ (_15419_, _09017_, \oc8051_golden_model_1.TL0 [4]);
  or _67063_ (_15420_, _15419_, _15418_);
  or _67064_ (_15421_, _15420_, _15417_);
  and _67065_ (_15422_, _09026_, \oc8051_golden_model_1.IP [4]);
  and _67066_ (_15423_, _09023_, \oc8051_golden_model_1.PSW [4]);
  and _67067_ (_15424_, _09030_, \oc8051_golden_model_1.B [4]);
  and _67068_ (_15425_, _09028_, \oc8051_golden_model_1.ACC [4]);
  or _67069_ (_15426_, _15425_, _15424_);
  or _67070_ (_15427_, _15426_, _15423_);
  or _67071_ (_15428_, _15427_, _15422_);
  and _67072_ (_15429_, _09035_, \oc8051_golden_model_1.SCON [4]);
  and _67073_ (_15430_, _09038_, \oc8051_golden_model_1.SBUF [4]);
  or _67074_ (_15431_, _15430_, _15429_);
  and _67075_ (_15432_, _09041_, \oc8051_golden_model_1.IE [4]);
  or _67076_ (_15433_, _15432_, _15431_);
  or _67077_ (_15434_, _15433_, _15428_);
  or _67078_ (_15435_, _15434_, _15421_);
  and _67079_ (_15436_, _09048_, \oc8051_golden_model_1.TH0 [4]);
  and _67080_ (_15437_, _09052_, \oc8051_golden_model_1.TL1 [4]);
  or _67081_ (_15438_, _15437_, _15436_);
  and _67082_ (_15439_, _09055_, \oc8051_golden_model_1.TCON [4]);
  and _67083_ (_15440_, _09059_, \oc8051_golden_model_1.PCON [4]);
  or _67084_ (_15441_, _15440_, _15439_);
  or _67085_ (_15442_, _15441_, _15438_);
  and _67086_ (_15443_, _09063_, \oc8051_golden_model_1.TMOD [4]);
  and _67087_ (_15444_, _09065_, \oc8051_golden_model_1.DPH [4]);
  or _67088_ (_15445_, _15444_, _15443_);
  and _67089_ (_15446_, _09068_, \oc8051_golden_model_1.DPL [4]);
  and _67090_ (_15447_, _09070_, \oc8051_golden_model_1.TH1 [4]);
  or _67091_ (_15448_, _15447_, _15446_);
  or _67092_ (_15449_, _15448_, _15445_);
  or _67093_ (_15450_, _15449_, _15442_);
  or _67094_ (_15451_, _15450_, _15435_);
  or _67095_ (_15452_, _15451_, _15410_);
  and _67096_ (_15453_, _15452_, _08841_);
  or _67097_ (_15454_, _15453_, _08848_);
  or _67098_ (_15455_, _15454_, _15409_);
  and _67099_ (_15456_, _08848_, _07093_);
  nor _67100_ (_15457_, _15456_, _06279_);
  and _67101_ (_15458_, _15457_, _15455_);
  and _67102_ (_15459_, _08995_, _06279_);
  or _67103_ (_15460_, _15459_, _06275_);
  or _67104_ (_15461_, _15460_, _15458_);
  nor _67105_ (_15462_, _12253_, _06009_);
  nor _67106_ (_15463_, _15462_, _07335_);
  and _67107_ (_15464_, _15463_, _15461_);
  or _67108_ (_15465_, _15464_, _15346_);
  and _67109_ (_15466_, _15465_, _09086_);
  and _67110_ (_15467_, _10590_, _07338_);
  or _67111_ (_15468_, _15467_, _15466_);
  and _67112_ (_15469_, _15468_, _09100_);
  and _67113_ (_15470_, _15343_, _07340_);
  or _67114_ (_15471_, _15470_, _15469_);
  and _67115_ (_15472_, _15471_, _07333_);
  and _67116_ (_15473_, _10571_, _07332_);
  or _67117_ (_15474_, _15473_, _07330_);
  or _67118_ (_15475_, _15474_, _15472_);
  nor _67119_ (_15476_, _12253_, _06018_);
  nor _67120_ (_15477_, _15476_, _09108_);
  and _67121_ (_15478_, _15477_, _15475_);
  and _67122_ (_15479_, _15342_, _09108_);
  or _67123_ (_15480_, _15479_, _09113_);
  or _67124_ (_15481_, _15480_, _15478_);
  nand _67125_ (_15482_, _10589_, _09113_);
  and _67126_ (_15483_, _15482_, _06016_);
  and _67127_ (_15484_, _15483_, _15481_);
  or _67128_ (_15485_, _07177_, _07043_);
  nor _67129_ (_15486_, _06320_, _07038_);
  nor _67130_ (_15487_, _12254_, _06016_);
  or _67131_ (_15488_, _15487_, _15486_);
  or _67132_ (_15489_, _15488_, _15485_);
  or _67133_ (_15490_, _15489_, _15484_);
  nand _67134_ (_15491_, _15490_, _15341_);
  and _67135_ (_15492_, _15491_, _15097_);
  and _67136_ (_15493_, _15340_, _07521_);
  or _67137_ (_15494_, _15493_, _15095_);
  or _67138_ (_15495_, _15494_, _15492_);
  nor _67139_ (_15496_, _09450_, _09265_);
  nor _67140_ (_15497_, _15496_, _09451_);
  or _67141_ (_15498_, _15497_, _15096_);
  nand _67142_ (_15499_, _15498_, _15495_);
  and _67143_ (_15500_, _15499_, _14943_);
  nor _67144_ (_15501_, _15497_, _14943_);
  or _67145_ (_15502_, _15501_, _15500_);
  and _67146_ (_15503_, _15502_, _09458_);
  and _67147_ (_15504_, _15367_, _07359_);
  or _67148_ (_15505_, _15504_, _06503_);
  or _67149_ (_15506_, _15505_, _15503_);
  nand _67150_ (_15507_, _12433_, _06503_);
  and _67151_ (_15508_, _15507_, _13082_);
  and _67152_ (_15509_, _15508_, _15506_);
  and _67153_ (_15510_, _12253_, _05998_);
  or _67154_ (_15511_, _15510_, _06272_);
  or _67155_ (_15512_, _15511_, _15509_);
  or _67156_ (_15513_, _15348_, _06273_);
  and _67157_ (_15514_, _15513_, _09473_);
  and _67158_ (_15515_, _15514_, _15512_);
  nor _67159_ (_15516_, _09485_, _09479_);
  nor _67160_ (_15517_, _15516_, _09486_);
  and _67161_ (_15518_, _15517_, _09474_);
  or _67162_ (_15519_, _15518_, _07055_);
  or _67163_ (_15520_, _15519_, _15515_);
  and _67164_ (_15521_, _15520_, _15337_);
  or _67165_ (_15522_, _15521_, _07379_);
  nor _67166_ (_15523_, _08599_, _08505_);
  nor _67167_ (_15524_, _15523_, _08600_);
  or _67168_ (_15525_, _15524_, _09495_);
  and _67169_ (_15526_, _15525_, _07631_);
  and _67170_ (_15527_, _15526_, _15522_);
  or _67171_ (_15528_, _15527_, _14560_);
  or _67172_ (_15529_, _14559_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _67173_ (_15530_, _15529_, _14733_);
  and _67174_ (_15531_, _15530_, _15528_);
  and _67175_ (_15532_, _12391_, _06503_);
  not _67176_ (_15533_, _12215_);
  nor _67177_ (_15534_, _15533_, _06503_);
  or _67178_ (_15535_, _15534_, _15532_);
  and _67179_ (_15536_, _15535_, _14732_);
  or _67180_ (_41546_, _15536_, _15531_);
  nor _67181_ (_15537_, _09486_, _09478_);
  nor _67182_ (_15538_, _15537_, _09487_);
  and _67183_ (_15539_, _15538_, _09474_);
  nor _67184_ (_15540_, _12249_, _06016_);
  nor _67185_ (_15541_, _08953_, _08307_);
  and _67186_ (_15542_, _15541_, _07340_);
  nand _67187_ (_15543_, _08832_, _08305_);
  nor _67188_ (_15544_, _13032_, _13031_);
  and _67189_ (_15545_, _13032_, \oc8051_golden_model_1.PSW [7]);
  or _67190_ (_15546_, _15545_, _15544_);
  and _67191_ (_15547_, _15546_, _07308_);
  or _67192_ (_15548_, _15544_, _08629_);
  nor _67193_ (_15549_, _15365_, _08307_);
  or _67194_ (_15550_, _15549_, _08787_);
  and _67195_ (_15551_, _15550_, _07276_);
  or _67196_ (_15552_, _09218_, _07270_);
  nor _67197_ (_15553_, _15338_, _08305_);
  nor _67198_ (_15554_, _15553_, _08679_);
  nor _67199_ (_15555_, _15554_, _08685_);
  nor _67200_ (_15556_, _06816_, _10237_);
  and _67201_ (_15557_, _12248_, _06816_);
  or _67202_ (_15558_, _15557_, _15556_);
  and _67203_ (_15559_, _15558_, _08685_);
  or _67204_ (_15560_, _15559_, _07269_);
  or _67205_ (_15561_, _15560_, _15555_);
  and _67206_ (_15562_, _15561_, _08782_);
  and _67207_ (_15563_, _15562_, _15552_);
  or _67208_ (_15564_, _15563_, _15551_);
  and _67209_ (_15565_, _15564_, _08670_);
  nand _67210_ (_15566_, _13033_, _13031_);
  and _67211_ (_15567_, _15566_, _07274_);
  or _67212_ (_15568_, _15567_, _07692_);
  or _67213_ (_15569_, _15568_, _15565_);
  nor _67214_ (_15570_, _12248_, _06052_);
  nor _67215_ (_15571_, _15570_, _07284_);
  and _67216_ (_15572_, _15571_, _15569_);
  and _67217_ (_15573_, _09478_, _07284_);
  or _67218_ (_15574_, _15573_, _07294_);
  or _67219_ (_15575_, _15574_, _15572_);
  and _67220_ (_15576_, _15575_, _15548_);
  or _67221_ (_15577_, _15576_, _06351_);
  nand _67222_ (_15578_, _08307_, _06351_);
  and _67223_ (_15579_, _15578_, _06349_);
  and _67224_ (_15580_, _15579_, _15577_);
  not _67225_ (_15581_, _13034_);
  and _67226_ (_15582_, _15566_, _15581_);
  and _67227_ (_15583_, _15582_, _06348_);
  or _67228_ (_15584_, _15583_, _15580_);
  and _67229_ (_15585_, _15584_, _06049_);
  nor _67230_ (_15586_, _12249_, _06049_);
  or _67231_ (_15587_, _15586_, _06441_);
  or _67232_ (_15588_, _15587_, _15585_);
  nand _67233_ (_15589_, _08307_, _06441_);
  and _67234_ (_15590_, _15589_, _15588_);
  or _67235_ (_15591_, _15590_, _07309_);
  and _67236_ (_15592_, _09218_, _06366_);
  nand _67237_ (_15593_, _08260_, _07309_);
  or _67238_ (_15594_, _15593_, _15592_);
  and _67239_ (_15595_, _15594_, _08821_);
  and _67240_ (_15596_, _15595_, _15591_);
  or _67241_ (_15597_, _15596_, _15547_);
  and _67242_ (_15598_, _15597_, _07745_);
  and _67243_ (_15599_, _12248_, _06039_);
  or _67244_ (_15600_, _15599_, _08832_);
  or _67245_ (_15601_, _15600_, _15598_);
  and _67246_ (_15602_, _15601_, _15543_);
  or _67247_ (_15603_, _15602_, _08838_);
  or _67248_ (_15604_, _09218_, _15010_);
  and _67249_ (_15605_, _15604_, _08842_);
  and _67250_ (_15606_, _15605_, _15603_);
  nor _67251_ (_15607_, _08880_, _08305_);
  and _67252_ (_15608_, _08989_, \oc8051_golden_model_1.P2INREG [5]);
  and _67253_ (_15609_, _08993_, \oc8051_golden_model_1.P0INREG [5]);
  and _67254_ (_15610_, _08998_, \oc8051_golden_model_1.P1INREG [5]);
  and _67255_ (_15611_, _09002_, \oc8051_golden_model_1.P3INREG [5]);
  or _67256_ (_15612_, _15611_, _15610_);
  or _67257_ (_15613_, _15612_, _15609_);
  or _67258_ (_15614_, _15613_, _15608_);
  and _67259_ (_15615_, _09010_, \oc8051_golden_model_1.SP [5]);
  and _67260_ (_15616_, _09017_, \oc8051_golden_model_1.TL0 [5]);
  or _67261_ (_15617_, _15616_, _15615_);
  or _67262_ (_15618_, _15617_, _15614_);
  and _67263_ (_15619_, _09026_, \oc8051_golden_model_1.IP [5]);
  and _67264_ (_15620_, _09023_, \oc8051_golden_model_1.PSW [5]);
  and _67265_ (_15621_, _09028_, \oc8051_golden_model_1.ACC [5]);
  and _67266_ (_15622_, _09030_, \oc8051_golden_model_1.B [5]);
  or _67267_ (_15623_, _15622_, _15621_);
  or _67268_ (_15624_, _15623_, _15620_);
  or _67269_ (_15625_, _15624_, _15619_);
  and _67270_ (_15626_, _09035_, \oc8051_golden_model_1.SCON [5]);
  and _67271_ (_15627_, _09038_, \oc8051_golden_model_1.SBUF [5]);
  or _67272_ (_15628_, _15627_, _15626_);
  and _67273_ (_15629_, _09041_, \oc8051_golden_model_1.IE [5]);
  or _67274_ (_15630_, _15629_, _15628_);
  or _67275_ (_15631_, _15630_, _15625_);
  or _67276_ (_15632_, _15631_, _15618_);
  and _67277_ (_15633_, _09048_, \oc8051_golden_model_1.TH0 [5]);
  and _67278_ (_15634_, _09052_, \oc8051_golden_model_1.TL1 [5]);
  or _67279_ (_15635_, _15634_, _15633_);
  and _67280_ (_15636_, _09055_, \oc8051_golden_model_1.TCON [5]);
  and _67281_ (_15637_, _09059_, \oc8051_golden_model_1.PCON [5]);
  or _67282_ (_15638_, _15637_, _15636_);
  or _67283_ (_15639_, _15638_, _15635_);
  and _67284_ (_15640_, _09063_, \oc8051_golden_model_1.TMOD [5]);
  and _67285_ (_15641_, _09065_, \oc8051_golden_model_1.DPH [5]);
  or _67286_ (_15642_, _15641_, _15640_);
  and _67287_ (_15643_, _09068_, \oc8051_golden_model_1.DPL [5]);
  and _67288_ (_15644_, _09070_, \oc8051_golden_model_1.TH1 [5]);
  or _67289_ (_15645_, _15644_, _15643_);
  or _67290_ (_15646_, _15645_, _15642_);
  or _67291_ (_15647_, _15646_, _15639_);
  or _67292_ (_15648_, _15647_, _15632_);
  or _67293_ (_15649_, _15648_, _15607_);
  and _67294_ (_15650_, _15649_, _08841_);
  or _67295_ (_15651_, _15650_, _08848_);
  or _67296_ (_15652_, _15651_, _15606_);
  and _67297_ (_15653_, _08848_, _06685_);
  nor _67298_ (_15654_, _15653_, _06279_);
  and _67299_ (_15655_, _15654_, _15652_);
  and _67300_ (_15656_, _08954_, _06279_);
  or _67301_ (_15657_, _15656_, _06275_);
  or _67302_ (_15658_, _15657_, _15655_);
  nor _67303_ (_15659_, _12248_, _06009_);
  nor _67304_ (_15660_, _15659_, _07335_);
  and _67305_ (_15661_, _15660_, _15658_);
  not _67306_ (_15662_, _15541_);
  nand _67307_ (_15663_, _08953_, _08307_);
  and _67308_ (_15664_, _15663_, _15662_);
  and _67309_ (_15665_, _15664_, _07335_);
  or _67310_ (_15666_, _15665_, _07338_);
  or _67311_ (_15667_, _15666_, _15661_);
  or _67312_ (_15668_, _12626_, _09086_);
  and _67313_ (_15669_, _15668_, _09100_);
  and _67314_ (_15670_, _15669_, _15667_);
  or _67315_ (_15671_, _15670_, _15542_);
  and _67316_ (_15672_, _15671_, _07333_);
  and _67317_ (_15673_, _10569_, _07332_);
  or _67318_ (_15674_, _15673_, _07330_);
  or _67319_ (_15675_, _15674_, _15672_);
  nor _67320_ (_15676_, _12248_, _06018_);
  nor _67321_ (_15677_, _15676_, _09108_);
  and _67322_ (_15678_, _15677_, _15675_);
  and _67323_ (_15679_, _15663_, _09108_);
  or _67324_ (_15680_, _15679_, _09113_);
  or _67325_ (_15681_, _15680_, _15678_);
  nand _67326_ (_15682_, _10570_, _09113_);
  and _67327_ (_15683_, _15682_, _06016_);
  and _67328_ (_15684_, _15683_, _15681_);
  nor _67329_ (_15685_, _15684_, _15540_);
  or _67330_ (_15686_, _15685_, _15091_);
  or _67331_ (_15687_, _15554_, _09122_);
  and _67332_ (_15688_, _15687_, _15097_);
  and _67333_ (_15689_, _15688_, _15686_);
  and _67334_ (_15690_, _15554_, _07521_);
  or _67335_ (_15691_, _15690_, _15095_);
  or _67336_ (_15692_, _15691_, _15689_);
  nor _67337_ (_15693_, _09451_, _09219_);
  nor _67338_ (_15694_, _15693_, _09452_);
  or _67339_ (_15695_, _15694_, _15096_);
  nand _67340_ (_15696_, _15695_, _15692_);
  and _67341_ (_15697_, _15696_, _14943_);
  nor _67342_ (_15698_, _15694_, _14943_);
  or _67343_ (_15699_, _15698_, _15697_);
  and _67344_ (_15700_, _15699_, _09458_);
  and _67345_ (_15701_, _15550_, _07359_);
  or _67346_ (_15702_, _15701_, _06503_);
  or _67347_ (_15703_, _15702_, _15700_);
  nand _67348_ (_15704_, _12428_, _06503_);
  and _67349_ (_15705_, _15704_, _13082_);
  and _67350_ (_15706_, _15705_, _15703_);
  and _67351_ (_15707_, _12248_, _05998_);
  or _67352_ (_15708_, _15707_, _06272_);
  or _67353_ (_15709_, _15708_, _15706_);
  or _67354_ (_15710_, _15544_, _06273_);
  and _67355_ (_15711_, _15710_, _09473_);
  and _67356_ (_15712_, _15711_, _15709_);
  or _67357_ (_15713_, _15712_, _15539_);
  and _67358_ (_15714_, _15713_, _07375_);
  or _67359_ (_15715_, _09500_, _09218_);
  nor _67360_ (_15716_, _09501_, _07375_);
  and _67361_ (_15717_, _15716_, _15715_);
  or _67362_ (_15718_, _15717_, _07379_);
  or _67363_ (_15719_, _15718_, _15714_);
  nor _67364_ (_15720_, _08600_, _08308_);
  nor _67365_ (_15721_, _15720_, _08601_);
  or _67366_ (_15722_, _15721_, _09495_);
  and _67367_ (_15723_, _15722_, _07631_);
  and _67368_ (_15724_, _15723_, _15719_);
  or _67369_ (_15725_, _15724_, _14560_);
  or _67370_ (_15726_, _14559_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _67371_ (_15727_, _15726_, _14733_);
  and _67372_ (_15728_, _15727_, _15725_);
  not _67373_ (_15729_, _12210_);
  nor _67374_ (_15730_, _15729_, _06503_);
  and _67375_ (_15731_, _12386_, _06503_);
  or _67376_ (_15732_, _15731_, _15730_);
  and _67377_ (_15733_, _15732_, _09525_);
  and _67378_ (_15734_, _15733_, _14731_);
  or _67379_ (_41548_, _15734_, _15728_);
  nor _67380_ (_15735_, _09501_, _09172_);
  nor _67381_ (_15736_, _15735_, _09502_);
  or _67382_ (_15737_, _15736_, _07375_);
  nor _67383_ (_15738_, _08679_, _08209_);
  nor _67384_ (_15739_, _15738_, _08680_);
  nand _67385_ (_15740_, _15739_, _15091_);
  or _67386_ (_15741_, _12240_, _06009_);
  nand _67387_ (_15742_, _08832_, _08209_);
  nor _67388_ (_15743_, _12980_, _12979_);
  and _67389_ (_15744_, _12980_, \oc8051_golden_model_1.PSW [7]);
  or _67390_ (_15745_, _15744_, _15743_);
  and _67391_ (_15746_, _15745_, _07308_);
  and _67392_ (_15747_, _09477_, _07284_);
  nand _67393_ (_15748_, _15739_, _08687_);
  and _67394_ (_15749_, _12240_, _06816_);
  or _67395_ (_15750_, _06816_, _10193_);
  nand _67396_ (_15751_, _15750_, _08685_);
  or _67397_ (_15752_, _15751_, _15749_);
  and _67398_ (_15753_, _15752_, _15748_);
  or _67399_ (_15754_, _15753_, _07269_);
  or _67400_ (_15755_, _09172_, _07270_);
  and _67401_ (_15756_, _15755_, _15754_);
  and _67402_ (_15757_, _15756_, _08782_);
  nor _67403_ (_15758_, _08787_, _08211_);
  or _67404_ (_15759_, _15758_, _08788_);
  and _67405_ (_15760_, _15759_, _07276_);
  or _67406_ (_15761_, _15760_, _15757_);
  and _67407_ (_15762_, _15761_, _08670_);
  nand _67408_ (_15763_, _12981_, _12979_);
  and _67409_ (_15764_, _15763_, _07274_);
  or _67410_ (_15765_, _15764_, _07692_);
  or _67411_ (_15766_, _15765_, _15762_);
  nor _67412_ (_15767_, _12240_, _06052_);
  nor _67413_ (_15768_, _15767_, _07284_);
  and _67414_ (_15769_, _15768_, _15766_);
  or _67415_ (_15770_, _15769_, _15747_);
  and _67416_ (_15771_, _15770_, _08629_);
  and _67417_ (_15772_, _15743_, _07294_);
  or _67418_ (_15773_, _15772_, _06351_);
  or _67419_ (_15774_, _15773_, _15771_);
  nand _67420_ (_15775_, _08211_, _06351_);
  and _67421_ (_15776_, _15775_, _06349_);
  and _67422_ (_15777_, _15776_, _15774_);
  not _67423_ (_15778_, _12982_);
  and _67424_ (_15779_, _15763_, _15778_);
  and _67425_ (_15780_, _15779_, _06348_);
  or _67426_ (_15781_, _15780_, _15777_);
  and _67427_ (_15782_, _15781_, _06049_);
  nor _67428_ (_15783_, _12241_, _06049_);
  or _67429_ (_15784_, _15783_, _06441_);
  or _67430_ (_15785_, _15784_, _15782_);
  nand _67431_ (_15786_, _08211_, _06441_);
  and _67432_ (_15787_, _15786_, _15785_);
  or _67433_ (_15788_, _15787_, _07309_);
  and _67434_ (_15789_, _09172_, _06366_);
  nand _67435_ (_15790_, _08164_, _07309_);
  or _67436_ (_15791_, _15790_, _15789_);
  and _67437_ (_15792_, _15791_, _08821_);
  and _67438_ (_15793_, _15792_, _15788_);
  or _67439_ (_15794_, _15793_, _15746_);
  and _67440_ (_15795_, _15794_, _07745_);
  and _67441_ (_15796_, _12240_, _06039_);
  or _67442_ (_15797_, _15796_, _08832_);
  or _67443_ (_15798_, _15797_, _15795_);
  and _67444_ (_15799_, _15798_, _15742_);
  or _67445_ (_15800_, _15799_, _08838_);
  or _67446_ (_15801_, _09172_, _15010_);
  and _67447_ (_15802_, _15801_, _08842_);
  and _67448_ (_15803_, _15802_, _15800_);
  nor _67449_ (_15804_, _08880_, _08209_);
  and _67450_ (_15805_, _08989_, \oc8051_golden_model_1.P2INREG [6]);
  and _67451_ (_15806_, _08993_, \oc8051_golden_model_1.P0INREG [6]);
  and _67452_ (_15807_, _08998_, \oc8051_golden_model_1.P1INREG [6]);
  and _67453_ (_15808_, _09002_, \oc8051_golden_model_1.P3INREG [6]);
  or _67454_ (_15809_, _15808_, _15807_);
  or _67455_ (_15810_, _15809_, _15806_);
  or _67456_ (_15811_, _15810_, _15805_);
  and _67457_ (_15812_, _09010_, \oc8051_golden_model_1.SP [6]);
  and _67458_ (_15813_, _09017_, \oc8051_golden_model_1.TL0 [6]);
  or _67459_ (_15814_, _15813_, _15812_);
  or _67460_ (_15815_, _15814_, _15811_);
  and _67461_ (_15816_, _09023_, \oc8051_golden_model_1.PSW [6]);
  and _67462_ (_15817_, _09026_, \oc8051_golden_model_1.IP [6]);
  and _67463_ (_15818_, _09030_, \oc8051_golden_model_1.B [6]);
  and _67464_ (_15819_, _09028_, \oc8051_golden_model_1.ACC [6]);
  or _67465_ (_15820_, _15819_, _15818_);
  or _67466_ (_15821_, _15820_, _15817_);
  or _67467_ (_15822_, _15821_, _15816_);
  and _67468_ (_15823_, _09035_, \oc8051_golden_model_1.SCON [6]);
  and _67469_ (_15824_, _09038_, \oc8051_golden_model_1.SBUF [6]);
  or _67470_ (_15825_, _15824_, _15823_);
  and _67471_ (_15826_, _09041_, \oc8051_golden_model_1.IE [6]);
  or _67472_ (_15827_, _15826_, _15825_);
  or _67473_ (_15828_, _15827_, _15822_);
  or _67474_ (_15829_, _15828_, _15815_);
  and _67475_ (_15830_, _09048_, \oc8051_golden_model_1.TH0 [6]);
  and _67476_ (_15831_, _09052_, \oc8051_golden_model_1.TL1 [6]);
  or _67477_ (_15832_, _15831_, _15830_);
  and _67478_ (_15833_, _09055_, \oc8051_golden_model_1.TCON [6]);
  and _67479_ (_15834_, _09059_, \oc8051_golden_model_1.PCON [6]);
  or _67480_ (_15835_, _15834_, _15833_);
  or _67481_ (_15836_, _15835_, _15832_);
  and _67482_ (_15837_, _09063_, \oc8051_golden_model_1.TMOD [6]);
  and _67483_ (_15838_, _09065_, \oc8051_golden_model_1.DPH [6]);
  or _67484_ (_15839_, _15838_, _15837_);
  and _67485_ (_15840_, _09068_, \oc8051_golden_model_1.DPL [6]);
  and _67486_ (_15841_, _09070_, \oc8051_golden_model_1.TH1 [6]);
  or _67487_ (_15842_, _15841_, _15840_);
  or _67488_ (_15843_, _15842_, _15839_);
  or _67489_ (_15844_, _15843_, _15836_);
  or _67490_ (_15845_, _15844_, _15829_);
  or _67491_ (_15846_, _15845_, _15804_);
  and _67492_ (_15847_, _15846_, _08841_);
  or _67493_ (_15848_, _15847_, _08848_);
  or _67494_ (_15849_, _15848_, _15803_);
  and _67495_ (_15850_, _08848_, _06397_);
  nor _67496_ (_15851_, _15850_, _06279_);
  and _67497_ (_15852_, _15851_, _15849_);
  not _67498_ (_15853_, _08918_);
  and _67499_ (_15854_, _15853_, _06279_);
  or _67500_ (_15855_, _15854_, _06275_);
  or _67501_ (_15856_, _15855_, _15852_);
  and _67502_ (_15857_, _15856_, _15741_);
  or _67503_ (_15858_, _15857_, _07335_);
  nand _67504_ (_15859_, _08918_, _08211_);
  nor _67505_ (_15860_, _08918_, _08211_);
  not _67506_ (_15861_, _15860_);
  and _67507_ (_15862_, _15861_, _15859_);
  or _67508_ (_15863_, _15862_, _07336_);
  and _67509_ (_15864_, _15863_, _09086_);
  and _67510_ (_15865_, _15864_, _15858_);
  nor _67511_ (_15866_, _10596_, _07340_);
  nor _67512_ (_15867_, _15866_, _07341_);
  or _67513_ (_15868_, _15867_, _15865_);
  or _67514_ (_15869_, _15860_, _09100_);
  and _67515_ (_15870_, _15869_, _07333_);
  and _67516_ (_15871_, _15870_, _15868_);
  and _67517_ (_15872_, _10568_, _07332_);
  or _67518_ (_15873_, _15872_, _07330_);
  or _67519_ (_15874_, _15873_, _15871_);
  nor _67520_ (_15875_, _12240_, _06018_);
  nor _67521_ (_15876_, _15875_, _09108_);
  and _67522_ (_15877_, _15876_, _15874_);
  and _67523_ (_15878_, _15859_, _09108_);
  or _67524_ (_15879_, _15878_, _09113_);
  or _67525_ (_15880_, _15879_, _15877_);
  nand _67526_ (_15881_, _10595_, _09113_);
  and _67527_ (_15882_, _15881_, _06016_);
  and _67528_ (_15883_, _15882_, _15880_);
  nor _67529_ (_15884_, _12241_, _06016_);
  or _67530_ (_15885_, _15884_, _15486_);
  or _67531_ (_15886_, _15885_, _15485_);
  or _67532_ (_15887_, _15886_, _15883_);
  nand _67533_ (_15888_, _15887_, _15740_);
  and _67534_ (_15889_, _15888_, _15097_);
  and _67535_ (_15890_, _15739_, _07521_);
  or _67536_ (_15891_, _15890_, _15095_);
  or _67537_ (_15892_, _15891_, _15889_);
  nor _67538_ (_15893_, _09452_, _09173_);
  nor _67539_ (_15894_, _15893_, _09453_);
  or _67540_ (_15895_, _15894_, _15096_);
  nand _67541_ (_15896_, _15895_, _15892_);
  and _67542_ (_15897_, _15896_, _14943_);
  nor _67543_ (_15898_, _15894_, _14943_);
  or _67544_ (_15899_, _15898_, _15897_);
  and _67545_ (_15900_, _15899_, _09458_);
  and _67546_ (_15901_, _15759_, _07359_);
  or _67547_ (_15902_, _15901_, _06503_);
  or _67548_ (_15903_, _15902_, _15900_);
  nand _67549_ (_15904_, _12420_, _06503_);
  and _67550_ (_15905_, _15904_, _13082_);
  and _67551_ (_15906_, _15905_, _15903_);
  and _67552_ (_15907_, _12240_, _05998_);
  or _67553_ (_15908_, _15907_, _06272_);
  or _67554_ (_15909_, _15908_, _15906_);
  or _67555_ (_15910_, _15743_, _06273_);
  and _67556_ (_15911_, _15910_, _09473_);
  and _67557_ (_15912_, _15911_, _15909_);
  nor _67558_ (_15913_, _09487_, _09477_);
  nor _67559_ (_15914_, _15913_, _09488_);
  and _67560_ (_15915_, _15914_, _09474_);
  or _67561_ (_15916_, _15915_, _07055_);
  or _67562_ (_15917_, _15916_, _15912_);
  and _67563_ (_15918_, _15917_, _15737_);
  or _67564_ (_15919_, _15918_, _07379_);
  nor _67565_ (_15920_, _08601_, _08212_);
  nor _67566_ (_15921_, _15920_, _08602_);
  or _67567_ (_15922_, _15921_, _09495_);
  and _67568_ (_15923_, _15922_, _07631_);
  and _67569_ (_15924_, _15923_, _15919_);
  or _67570_ (_15925_, _15924_, _14560_);
  or _67571_ (_15926_, _14559_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _67572_ (_15927_, _15926_, _14733_);
  and _67573_ (_15928_, _15927_, _15925_);
  and _67574_ (_15929_, _12381_, _06503_);
  not _67575_ (_15930_, _12205_);
  nor _67576_ (_15931_, _15930_, _06503_);
  or _67577_ (_15932_, _15931_, _15929_);
  and _67578_ (_15933_, _15932_, _09525_);
  and _67579_ (_15934_, _15933_, _14731_);
  or _67580_ (_41549_, _15934_, _15928_);
  or _67581_ (_15935_, _14560_, _09510_);
  or _67582_ (_15936_, _14559_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _67583_ (_15937_, _15936_, _14733_);
  and _67584_ (_15938_, _15937_, _15935_);
  and _67585_ (_15939_, _14732_, _09567_);
  or _67586_ (_41550_, _15939_, _15938_);
  and _67587_ (_15940_, _14554_, _07542_);
  and _67588_ (_15941_, _15940_, _14557_);
  not _67589_ (_15942_, _15941_);
  or _67590_ (_15943_, _15942_, _14727_);
  or _67591_ (_15944_, _15941_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _67592_ (_15945_, _14730_, _07684_);
  and _67593_ (_15946_, _15945_, _09525_);
  not _67594_ (_15947_, _15946_);
  and _67595_ (_15948_, _15947_, _15944_);
  and _67596_ (_15949_, _15948_, _15943_);
  and _67597_ (_15950_, _09525_, _07684_);
  and _67598_ (_15951_, _15950_, _14730_);
  and _67599_ (_15952_, _15951_, _14740_);
  or _67600_ (_41554_, _15952_, _15949_);
  or _67601_ (_15953_, _15942_, _14929_);
  or _67602_ (_15954_, _15941_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _67603_ (_15955_, _15954_, _15947_);
  and _67604_ (_15956_, _15955_, _15953_);
  and _67605_ (_15957_, _15951_, _14938_);
  or _67606_ (_41556_, _15957_, _15956_);
  or _67607_ (_15958_, _15942_, _15132_);
  or _67608_ (_15959_, _15941_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _67609_ (_15960_, _15959_, _15947_);
  and _67610_ (_15961_, _15960_, _15958_);
  and _67611_ (_15962_, _15945_, _15140_);
  or _67612_ (_41557_, _15962_, _15961_);
  or _67613_ (_15963_, _15942_, _15324_);
  or _67614_ (_15964_, _15941_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _67615_ (_15965_, _15964_, _15947_);
  and _67616_ (_15966_, _15965_, _15963_);
  and _67617_ (_15967_, _15951_, _15333_);
  or _67618_ (_41558_, _15967_, _15966_);
  or _67619_ (_15968_, _15942_, _15527_);
  or _67620_ (_15969_, _15941_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _67621_ (_15970_, _15969_, _15947_);
  and _67622_ (_15971_, _15970_, _15968_);
  and _67623_ (_15972_, _15946_, _15535_);
  or _67624_ (_41559_, _15972_, _15971_);
  or _67625_ (_15973_, _15942_, _15724_);
  or _67626_ (_15974_, _15941_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _67627_ (_15975_, _15974_, _15947_);
  and _67628_ (_15976_, _15975_, _15973_);
  and _67629_ (_15977_, _15945_, _15733_);
  or _67630_ (_41560_, _15977_, _15976_);
  or _67631_ (_15978_, _15942_, _15924_);
  or _67632_ (_15979_, _15941_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _67633_ (_15980_, _15979_, _15947_);
  and _67634_ (_15981_, _15980_, _15978_);
  and _67635_ (_15982_, _15951_, _15933_);
  or _67636_ (_41562_, _15982_, _15981_);
  or _67637_ (_15983_, _15942_, _09511_);
  or _67638_ (_15984_, _15941_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _67639_ (_15985_, _15984_, _15947_);
  and _67640_ (_15986_, _15985_, _15983_);
  and _67641_ (_15987_, _15946_, _09567_);
  or _67642_ (_41563_, _15987_, _15986_);
  not _67643_ (_15988_, _07382_);
  and _67644_ (_15989_, _07633_, _15988_);
  and _67645_ (_15990_, _15989_, _14557_);
  not _67646_ (_15991_, _15990_);
  or _67647_ (_15992_, _15991_, _14727_);
  or _67648_ (_15993_, _15990_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _67649_ (_15994_, _14730_, _08695_);
  nand _67650_ (_15995_, _15994_, _09525_);
  and _67651_ (_15996_, _15995_, _15993_);
  and _67652_ (_15997_, _15996_, _15992_);
  and _67653_ (_15998_, _09525_, _08695_);
  and _67654_ (_15999_, _15998_, _14730_);
  and _67655_ (_16000_, _15999_, _14740_);
  or _67656_ (_41567_, _16000_, _15997_);
  or _67657_ (_16001_, _15991_, _14929_);
  nor _67658_ (_16002_, _15990_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor _67659_ (_16003_, _16002_, _15999_);
  and _67660_ (_16004_, _16003_, _16001_);
  and _67661_ (_16005_, _15994_, _14938_);
  or _67662_ (_41568_, _16005_, _16004_);
  or _67663_ (_16006_, _15991_, _15132_);
  or _67664_ (_16007_, _15990_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _67665_ (_16008_, _16007_, _15995_);
  and _67666_ (_16009_, _16008_, _16006_);
  and _67667_ (_16010_, _15994_, _15140_);
  or _67668_ (_41570_, _16010_, _16009_);
  or _67669_ (_16011_, _15991_, _15324_);
  or _67670_ (_16012_, _15990_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _67671_ (_16013_, _16012_, _15995_);
  and _67672_ (_16014_, _16013_, _16011_);
  and _67673_ (_16015_, _15999_, _15333_);
  or _67674_ (_41571_, _16015_, _16014_);
  or _67675_ (_16016_, _15991_, _15527_);
  or _67676_ (_16017_, _15990_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _67677_ (_16018_, _16017_, _15995_);
  and _67678_ (_16019_, _16018_, _16016_);
  and _67679_ (_16020_, _15999_, _15535_);
  or _67680_ (_41572_, _16020_, _16019_);
  or _67681_ (_16021_, _15991_, _15724_);
  or _67682_ (_16022_, _15990_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _67683_ (_16023_, _16022_, _15995_);
  and _67684_ (_16024_, _16023_, _16021_);
  and _67685_ (_16025_, _15994_, _15733_);
  or _67686_ (_41573_, _16025_, _16024_);
  or _67687_ (_16026_, _15991_, _15924_);
  or _67688_ (_16027_, _15990_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _67689_ (_16028_, _16027_, _15995_);
  and _67690_ (_16029_, _16028_, _16026_);
  and _67691_ (_16030_, _15999_, _15933_);
  or _67692_ (_41574_, _16030_, _16029_);
  or _67693_ (_16031_, _15991_, _09511_);
  nor _67694_ (_16032_, _15990_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _67695_ (_16033_, _16032_, _15999_);
  and _67696_ (_16034_, _16033_, _16031_);
  and _67697_ (_16035_, _15994_, _09568_);
  or _67698_ (_41576_, _16035_, _16034_);
  and _67699_ (_16036_, _14557_, _07634_);
  or _67700_ (_16037_, _16036_, \oc8051_golden_model_1.IRAM[3] [0]);
  not _67701_ (_16038_, _16036_);
  or _67702_ (_16039_, _16038_, _14727_);
  and _67703_ (_16040_, _14730_, _07386_);
  and _67704_ (_16041_, _16040_, _09525_);
  not _67705_ (_16042_, _16041_);
  and _67706_ (_16043_, _16042_, _16039_);
  and _67707_ (_16044_, _16043_, _16037_);
  and _67708_ (_16045_, _16040_, _14740_);
  or _67709_ (_41579_, _16045_, _16044_);
  nor _67710_ (_16046_, _16036_, _07400_);
  and _67711_ (_16047_, _16036_, _14929_);
  or _67712_ (_16048_, _16047_, _16046_);
  and _67713_ (_16049_, _16048_, _16042_);
  and _67714_ (_16050_, _16040_, _14938_);
  or _67715_ (_41581_, _16050_, _16049_);
  or _67716_ (_16051_, _16038_, _15132_);
  or _67717_ (_16052_, _16036_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _67718_ (_16053_, _16052_, _16042_);
  and _67719_ (_16054_, _16053_, _16051_);
  and _67720_ (_16055_, _16040_, _15140_);
  or _67721_ (_41582_, _16055_, _16054_);
  or _67722_ (_16056_, _16036_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _67723_ (_16057_, _16056_, _16042_);
  or _67724_ (_16058_, _16038_, _15324_);
  and _67725_ (_16059_, _16058_, _16057_);
  and _67726_ (_16060_, _16040_, _15333_);
  or _67727_ (_41583_, _16060_, _16059_);
  or _67728_ (_16061_, _16036_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _67729_ (_16062_, _16061_, _16042_);
  or _67730_ (_16063_, _16038_, _15527_);
  and _67731_ (_16064_, _16063_, _16062_);
  and _67732_ (_16065_, _16041_, _15535_);
  or _67733_ (_41584_, _16065_, _16064_);
  or _67734_ (_16066_, _16036_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _67735_ (_16067_, _16066_, _16042_);
  or _67736_ (_16068_, _16038_, _15724_);
  and _67737_ (_16069_, _16068_, _16067_);
  and _67738_ (_16070_, _16040_, _15733_);
  or _67739_ (_41585_, _16070_, _16069_);
  or _67740_ (_16071_, _16036_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _67741_ (_16072_, _16071_, _16042_);
  or _67742_ (_16073_, _16038_, _15924_);
  and _67743_ (_16074_, _16073_, _16072_);
  and _67744_ (_16075_, _16040_, _15933_);
  or _67745_ (_41587_, _16075_, _16074_);
  or _67746_ (_16076_, _16036_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _67747_ (_16077_, _16076_, _16042_);
  or _67748_ (_16078_, _16038_, _09511_);
  and _67749_ (_16079_, _16078_, _16077_);
  and _67750_ (_16080_, _16041_, _09567_);
  or _67751_ (_41588_, _16080_, _16079_);
  and _67752_ (_16081_, _07941_, _07798_);
  and _67753_ (_16082_, _16081_, _14555_);
  not _67754_ (_16083_, _16082_);
  or _67755_ (_16084_, _16083_, _14727_);
  not _67756_ (_16085_, _09518_);
  and _67757_ (_16086_, _09526_, _16085_);
  and _67758_ (_16087_, _16086_, _07387_);
  not _67759_ (_16088_, _16087_);
  or _67760_ (_16089_, _16082_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _67761_ (_16090_, _16089_, _16088_);
  and _67762_ (_16091_, _16090_, _16084_);
  and _67763_ (_16092_, _16087_, _14740_);
  or _67764_ (_41592_, _16092_, _16091_);
  or _67765_ (_16093_, _16083_, _14929_);
  or _67766_ (_16094_, _16082_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _67767_ (_16095_, _16094_, _16088_);
  and _67768_ (_16096_, _16095_, _16093_);
  and _67769_ (_16097_, _16087_, _14938_);
  or _67770_ (_41593_, _16097_, _16096_);
  or _67771_ (_16098_, _16083_, _15132_);
  or _67772_ (_16099_, _16082_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _67773_ (_16100_, _16099_, _16088_);
  and _67774_ (_16101_, _16100_, _16098_);
  and _67775_ (_16102_, _16087_, _15140_);
  or _67776_ (_41594_, _16102_, _16101_);
  or _67777_ (_16103_, _16083_, _15324_);
  or _67778_ (_16104_, _16082_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _67779_ (_16105_, _16104_, _16088_);
  and _67780_ (_16106_, _16105_, _16103_);
  and _67781_ (_16107_, _16087_, _15333_);
  or _67782_ (_41595_, _16107_, _16106_);
  or _67783_ (_16108_, _16083_, _15527_);
  or _67784_ (_16109_, _16082_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _67785_ (_16110_, _16109_, _16088_);
  and _67786_ (_16111_, _16110_, _16108_);
  and _67787_ (_16112_, _15535_, _09525_);
  and _67788_ (_16113_, _16112_, _16087_);
  or _67789_ (_41596_, _16113_, _16111_);
  or _67790_ (_16114_, _16083_, _15724_);
  or _67791_ (_16115_, _16082_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _67792_ (_16116_, _16115_, _16088_);
  and _67793_ (_16117_, _16116_, _16114_);
  and _67794_ (_16118_, _16087_, _15733_);
  or _67795_ (_41597_, _16118_, _16117_);
  or _67796_ (_16119_, _16083_, _15924_);
  or _67797_ (_16120_, _16082_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _67798_ (_16121_, _16120_, _16088_);
  and _67799_ (_16122_, _16121_, _16119_);
  and _67800_ (_16123_, _16087_, _15933_);
  or _67801_ (_41598_, _16123_, _16122_);
  or _67802_ (_16124_, _16082_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _67803_ (_16125_, _16083_, _09511_);
  and _67804_ (_16126_, _16125_, _16124_);
  or _67805_ (_16127_, _16126_, _16087_);
  or _67806_ (_16128_, _16088_, _09568_);
  and _67807_ (_41601_, _16128_, _16127_);
  and _67808_ (_16129_, _16081_, _15940_);
  not _67809_ (_16130_, _16129_);
  or _67810_ (_16131_, _16130_, _14727_);
  and _67811_ (_16132_, _16086_, _07684_);
  not _67812_ (_16133_, _16132_);
  or _67813_ (_16134_, _16129_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _67814_ (_16135_, _16134_, _16133_);
  and _67815_ (_16136_, _16135_, _16131_);
  and _67816_ (_16137_, _16132_, _14740_);
  or _67817_ (_41604_, _16137_, _16136_);
  or _67818_ (_16138_, _16130_, _14929_);
  or _67819_ (_16139_, _16129_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _67820_ (_16140_, _16139_, _16133_);
  and _67821_ (_16141_, _16140_, _16138_);
  and _67822_ (_16142_, _16132_, _14938_);
  or _67823_ (_41605_, _16142_, _16141_);
  or _67824_ (_16143_, _16130_, _15132_);
  or _67825_ (_16144_, _16129_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _67826_ (_16145_, _16144_, _16133_);
  and _67827_ (_16146_, _16145_, _16143_);
  and _67828_ (_16147_, _16132_, _15140_);
  or _67829_ (_41607_, _16147_, _16146_);
  or _67830_ (_16148_, _16130_, _15324_);
  or _67831_ (_16149_, _16129_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _67832_ (_16150_, _16149_, _16133_);
  and _67833_ (_16151_, _16150_, _16148_);
  and _67834_ (_16152_, _16132_, _15333_);
  or _67835_ (_41608_, _16152_, _16151_);
  or _67836_ (_16153_, _16130_, _15527_);
  or _67837_ (_16154_, _16129_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _67838_ (_16155_, _16154_, _16133_);
  and _67839_ (_16156_, _16155_, _16153_);
  and _67840_ (_16157_, _16132_, _16112_);
  or _67841_ (_41609_, _16157_, _16156_);
  or _67842_ (_16158_, _16130_, _15724_);
  or _67843_ (_16159_, _16129_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _67844_ (_16160_, _16159_, _16133_);
  and _67845_ (_16161_, _16160_, _16158_);
  and _67846_ (_16162_, _16132_, _15733_);
  or _67847_ (_41610_, _16162_, _16161_);
  or _67848_ (_16163_, _16130_, _15924_);
  or _67849_ (_16164_, _16129_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _67850_ (_16165_, _16164_, _16133_);
  and _67851_ (_16166_, _16165_, _16163_);
  and _67852_ (_16167_, _16132_, _15933_);
  or _67853_ (_41611_, _16167_, _16166_);
  or _67854_ (_16168_, _16130_, _09511_);
  or _67855_ (_16169_, _16129_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _67856_ (_16170_, _16169_, _16133_);
  and _67857_ (_16171_, _16170_, _16168_);
  and _67858_ (_16172_, _16132_, _09568_);
  or _67859_ (_41613_, _16172_, _16171_);
  and _67860_ (_16173_, _16081_, _15989_);
  not _67861_ (_16174_, _16173_);
  or _67862_ (_16175_, _16174_, _14727_);
  and _67863_ (_16176_, _16086_, _08695_);
  not _67864_ (_16177_, _16176_);
  or _67865_ (_16178_, _16173_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _67866_ (_16179_, _16178_, _16177_);
  and _67867_ (_16180_, _16179_, _16175_);
  and _67868_ (_16181_, _16176_, _14740_);
  or _67869_ (_41616_, _16181_, _16180_);
  or _67870_ (_16182_, _16174_, _14929_);
  or _67871_ (_16183_, _16173_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _67872_ (_16184_, _16183_, _16177_);
  and _67873_ (_16185_, _16184_, _16182_);
  and _67874_ (_16186_, _16176_, _14938_);
  or _67875_ (_41618_, _16186_, _16185_);
  or _67876_ (_16187_, _16174_, _15132_);
  or _67877_ (_16188_, _16173_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _67878_ (_16189_, _16188_, _16177_);
  and _67879_ (_16190_, _16189_, _16187_);
  and _67880_ (_16191_, _16176_, _15140_);
  or _67881_ (_41619_, _16191_, _16190_);
  or _67882_ (_16192_, _16174_, _15324_);
  or _67883_ (_16193_, _16173_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _67884_ (_16194_, _16193_, _16177_);
  and _67885_ (_16195_, _16194_, _16192_);
  and _67886_ (_16196_, _16176_, _15333_);
  or _67887_ (_41620_, _16196_, _16195_);
  or _67888_ (_16197_, _16174_, _15527_);
  or _67889_ (_16198_, _16173_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _67890_ (_16199_, _16198_, _16177_);
  and _67891_ (_16200_, _16199_, _16197_);
  and _67892_ (_16201_, _16176_, _16112_);
  or _67893_ (_41621_, _16201_, _16200_);
  or _67894_ (_16202_, _16174_, _15724_);
  or _67895_ (_16203_, _16173_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _67896_ (_16204_, _16203_, _16177_);
  and _67897_ (_16205_, _16204_, _16202_);
  and _67898_ (_16206_, _16176_, _15733_);
  or _67899_ (_41622_, _16206_, _16205_);
  or _67900_ (_16207_, _16174_, _15924_);
  or _67901_ (_16208_, _16173_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _67902_ (_16209_, _16208_, _16177_);
  and _67903_ (_16210_, _16209_, _16207_);
  and _67904_ (_16211_, _16176_, _15933_);
  or _67905_ (_41624_, _16211_, _16210_);
  nor _67906_ (_16212_, _16173_, _08064_);
  and _67907_ (_16213_, _16173_, _09511_);
  or _67908_ (_16214_, _16213_, _16212_);
  and _67909_ (_16215_, _16214_, _16177_);
  and _67910_ (_16216_, _16176_, _09568_);
  or _67911_ (_41625_, _16216_, _16215_);
  and _67912_ (_16217_, _16086_, _07386_);
  not _67913_ (_16218_, _16217_);
  or _67914_ (_16219_, _16218_, _14740_);
  and _67915_ (_16220_, _16081_, _07634_);
  and _67916_ (_16221_, _16220_, _14727_);
  nor _67917_ (_16222_, _16220_, _07211_);
  or _67918_ (_16223_, _16222_, _16217_);
  or _67919_ (_16224_, _16223_, _16221_);
  and _67920_ (_41628_, _16224_, _16219_);
  nor _67921_ (_16225_, _16220_, _07408_);
  and _67922_ (_16226_, _16220_, _14929_);
  or _67923_ (_16227_, _16226_, _16225_);
  and _67924_ (_16228_, _16227_, _16218_);
  and _67925_ (_16229_, _16217_, _14938_);
  or _67926_ (_41630_, _16229_, _16228_);
  or _67927_ (_16230_, _16220_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _67928_ (_16231_, _16230_, _16218_);
  not _67929_ (_16232_, _16220_);
  or _67930_ (_16233_, _16232_, _15132_);
  and _67931_ (_16234_, _16233_, _16231_);
  and _67932_ (_16235_, _16217_, _15140_);
  or _67933_ (_41631_, _16235_, _16234_);
  or _67934_ (_16236_, _16220_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _67935_ (_16237_, _16236_, _16218_);
  or _67936_ (_16238_, _16232_, _15324_);
  and _67937_ (_16239_, _16238_, _16237_);
  and _67938_ (_16240_, _16217_, _15333_);
  or _67939_ (_41632_, _16240_, _16239_);
  or _67940_ (_16241_, _16220_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _67941_ (_16242_, _16241_, _16218_);
  or _67942_ (_16243_, _16232_, _15527_);
  and _67943_ (_16244_, _16243_, _16242_);
  and _67944_ (_16245_, _16217_, _16112_);
  or _67945_ (_41633_, _16245_, _16244_);
  or _67946_ (_16246_, _16220_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _67947_ (_16247_, _16246_, _16218_);
  or _67948_ (_16248_, _16232_, _15724_);
  and _67949_ (_16249_, _16248_, _16247_);
  and _67950_ (_16250_, _16217_, _15733_);
  or _67951_ (_41634_, _16250_, _16249_);
  or _67952_ (_16251_, _16220_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _67953_ (_16252_, _16251_, _16218_);
  or _67954_ (_16253_, _16232_, _15924_);
  and _67955_ (_16254_, _16253_, _16252_);
  and _67956_ (_16255_, _16217_, _15933_);
  or _67957_ (_41636_, _16255_, _16254_);
  or _67958_ (_16256_, _16218_, _09568_);
  or _67959_ (_16257_, _16220_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _67960_ (_16258_, _16232_, _09511_);
  and _67961_ (_16259_, _16258_, _16257_);
  or _67962_ (_16260_, _16259_, _16217_);
  and _67963_ (_41637_, _16260_, _16256_);
  and _67964_ (_16261_, _14556_, _07940_);
  and _67965_ (_16262_, _16261_, _14555_);
  not _67966_ (_16263_, _16262_);
  or _67967_ (_16264_, _16263_, _14727_);
  not _67968_ (_16265_, _09521_);
  and _67969_ (_16266_, _09531_, _16265_);
  and _67970_ (_16267_, _16266_, _07387_);
  nor _67971_ (_16268_, _16262_, \oc8051_golden_model_1.IRAM[8] [0]);
  nor _67972_ (_16269_, _16268_, _16267_);
  and _67973_ (_16270_, _16269_, _16264_);
  and _67974_ (_16271_, _16267_, _14740_);
  or _67975_ (_41641_, _16271_, _16270_);
  or _67976_ (_16272_, _16263_, _14929_);
  nand _67977_ (_16273_, _09531_, _09516_);
  or _67978_ (_16274_, _16262_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _67979_ (_16275_, _16274_, _16273_);
  and _67980_ (_16276_, _16275_, _16272_);
  and _67981_ (_16277_, _16267_, _14938_);
  or _67982_ (_41642_, _16277_, _16276_);
  or _67983_ (_16278_, _16263_, _15132_);
  or _67984_ (_16279_, _16262_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _67985_ (_16280_, _16279_, _16273_);
  and _67986_ (_16281_, _16280_, _16278_);
  and _67987_ (_16282_, _16267_, _15140_);
  or _67988_ (_41644_, _16282_, _16281_);
  or _67989_ (_16283_, _16263_, _15324_);
  or _67990_ (_16284_, _16262_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _67991_ (_16285_, _16284_, _16273_);
  and _67992_ (_16286_, _16285_, _16283_);
  and _67993_ (_16287_, _16267_, _15333_);
  or _67994_ (_41645_, _16287_, _16286_);
  or _67995_ (_16288_, _16263_, _15527_);
  or _67996_ (_16289_, _16262_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _67997_ (_16290_, _16289_, _16273_);
  and _67998_ (_16291_, _16290_, _16288_);
  and _67999_ (_16292_, _16267_, _16112_);
  or _68000_ (_41646_, _16292_, _16291_);
  or _68001_ (_16293_, _16263_, _15724_);
  or _68002_ (_16294_, _16262_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _68003_ (_16295_, _16294_, _16273_);
  and _68004_ (_16296_, _16295_, _16293_);
  and _68005_ (_16297_, _16267_, _15733_);
  or _68006_ (_41647_, _16297_, _16296_);
  or _68007_ (_16298_, _16263_, _15924_);
  or _68008_ (_16299_, _16262_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _68009_ (_16300_, _16299_, _16273_);
  and _68010_ (_16301_, _16300_, _16298_);
  and _68011_ (_16302_, _16267_, _15933_);
  or _68012_ (_41648_, _16302_, _16301_);
  or _68013_ (_16303_, _16263_, _09511_);
  nor _68014_ (_16304_, _16262_, \oc8051_golden_model_1.IRAM[8] [7]);
  nor _68015_ (_16305_, _16304_, _16267_);
  and _68016_ (_16306_, _16305_, _16303_);
  and _68017_ (_16307_, _16267_, _09568_);
  or _68018_ (_41649_, _16307_, _16306_);
  and _68019_ (_16308_, _16261_, _15940_);
  not _68020_ (_16309_, _16308_);
  or _68021_ (_16310_, _16309_, _14727_);
  and _68022_ (_16311_, _16266_, _07684_);
  nor _68023_ (_16312_, _16308_, \oc8051_golden_model_1.IRAM[9] [0]);
  nor _68024_ (_16313_, _16312_, _16311_);
  and _68025_ (_16314_, _16313_, _16310_);
  and _68026_ (_16315_, _16311_, _14740_);
  or _68027_ (_41652_, _16315_, _16314_);
  or _68028_ (_16316_, _16309_, _14929_);
  nand _68029_ (_16317_, _09531_, _07685_);
  or _68030_ (_16318_, _16308_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _68031_ (_16319_, _16318_, _16317_);
  and _68032_ (_16320_, _16319_, _16316_);
  and _68033_ (_16321_, _16311_, _14938_);
  or _68034_ (_41653_, _16321_, _16320_);
  or _68035_ (_16322_, _16309_, _15132_);
  or _68036_ (_16323_, _16308_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _68037_ (_16324_, _16323_, _16317_);
  and _68038_ (_16325_, _16324_, _16322_);
  and _68039_ (_16326_, _16311_, _15140_);
  or _68040_ (_41656_, _16326_, _16325_);
  or _68041_ (_16327_, _16309_, _15324_);
  or _68042_ (_16328_, _16308_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _68043_ (_16329_, _16328_, _16317_);
  and _68044_ (_16330_, _16329_, _16327_);
  and _68045_ (_16331_, _16311_, _15333_);
  or _68046_ (_41657_, _16331_, _16330_);
  or _68047_ (_16332_, _16309_, _15527_);
  or _68048_ (_16333_, _16308_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _68049_ (_16334_, _16333_, _16317_);
  and _68050_ (_16335_, _16334_, _16332_);
  and _68051_ (_16336_, _16311_, _16112_);
  or _68052_ (_41658_, _16336_, _16335_);
  or _68053_ (_16337_, _16309_, _15724_);
  or _68054_ (_16338_, _16308_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _68055_ (_16339_, _16338_, _16317_);
  and _68056_ (_16340_, _16339_, _16337_);
  and _68057_ (_16341_, _16311_, _15733_);
  or _68058_ (_41659_, _16341_, _16340_);
  or _68059_ (_16342_, _16309_, _15924_);
  or _68060_ (_16343_, _16308_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _68061_ (_16344_, _16343_, _16317_);
  and _68062_ (_16345_, _16344_, _16342_);
  and _68063_ (_16346_, _16311_, _15933_);
  or _68064_ (_41660_, _16346_, _16345_);
  or _68065_ (_16347_, _16309_, _09511_);
  nor _68066_ (_16348_, _16308_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor _68067_ (_16349_, _16348_, _16311_);
  and _68068_ (_16350_, _16349_, _16347_);
  and _68069_ (_16351_, _16311_, _09568_);
  or _68070_ (_41662_, _16351_, _16350_);
  and _68071_ (_16352_, _16261_, _15989_);
  not _68072_ (_16353_, _16352_);
  or _68073_ (_16354_, _16353_, _14727_);
  and _68074_ (_16355_, _16266_, _08695_);
  not _68075_ (_16356_, _16355_);
  or _68076_ (_16357_, _16352_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _68077_ (_16358_, _16357_, _16356_);
  and _68078_ (_16359_, _16358_, _16354_);
  and _68079_ (_16360_, _16355_, _14740_);
  or _68080_ (_41665_, _16360_, _16359_);
  or _68081_ (_16361_, _16353_, _14929_);
  or _68082_ (_16362_, _16352_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _68083_ (_16363_, _16362_, _16356_);
  and _68084_ (_16364_, _16363_, _16361_);
  and _68085_ (_16365_, _16355_, _14938_);
  or _68086_ (_41667_, _16365_, _16364_);
  or _68087_ (_16366_, _16353_, _15132_);
  or _68088_ (_16367_, _16352_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _68089_ (_16368_, _16367_, _16356_);
  and _68090_ (_16369_, _16368_, _16366_);
  and _68091_ (_16370_, _16355_, _15140_);
  or _68092_ (_41668_, _16370_, _16369_);
  or _68093_ (_16371_, _16353_, _15324_);
  or _68094_ (_16372_, _16352_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _68095_ (_16373_, _16372_, _16356_);
  and _68096_ (_16374_, _16373_, _16371_);
  and _68097_ (_16375_, _16355_, _15333_);
  or _68098_ (_41669_, _16375_, _16374_);
  or _68099_ (_16376_, _16353_, _15527_);
  or _68100_ (_16377_, _16352_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _68101_ (_16378_, _16377_, _16356_);
  and _68102_ (_16379_, _16378_, _16376_);
  and _68103_ (_16380_, _16355_, _16112_);
  or _68104_ (_41670_, _16380_, _16379_);
  or _68105_ (_16381_, _16353_, _15724_);
  or _68106_ (_16382_, _16352_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _68107_ (_16383_, _16382_, _16356_);
  and _68108_ (_16384_, _16383_, _16381_);
  and _68109_ (_16385_, _16355_, _15733_);
  or _68110_ (_41671_, _16385_, _16384_);
  or _68111_ (_16386_, _16353_, _15924_);
  or _68112_ (_16387_, _16352_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _68113_ (_16388_, _16387_, _16356_);
  and _68114_ (_16389_, _16388_, _16386_);
  and _68115_ (_16390_, _16355_, _15933_);
  or _68116_ (_41673_, _16390_, _16389_);
  or _68117_ (_16391_, _16353_, _09511_);
  or _68118_ (_16392_, _16352_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _68119_ (_16393_, _16392_, _16356_);
  and _68120_ (_16394_, _16393_, _16391_);
  and _68121_ (_16395_, _16355_, _09568_);
  or _68122_ (_41674_, _16395_, _16394_);
  and _68123_ (_16396_, _16266_, _07386_);
  not _68124_ (_16397_, _16396_);
  or _68125_ (_16398_, _16397_, _14739_);
  and _68126_ (_16399_, _16261_, _07634_);
  and _68127_ (_16400_, _16399_, _14727_);
  not _68128_ (_16401_, _16399_);
  and _68129_ (_16402_, _16401_, \oc8051_golden_model_1.IRAM[11] [0]);
  or _68130_ (_16403_, _16402_, _16396_);
  or _68131_ (_16404_, _16403_, _16400_);
  and _68132_ (_41677_, _16404_, _16398_);
  nor _68133_ (_16405_, _16399_, _07422_);
  and _68134_ (_16406_, _16399_, _14929_);
  or _68135_ (_16407_, _16406_, _16405_);
  and _68136_ (_16408_, _16407_, _16397_);
  and _68137_ (_16409_, _16396_, _14938_);
  or _68138_ (_41679_, _16409_, _16408_);
  not _68139_ (_16410_, _07542_);
  and _68140_ (_16411_, _14554_, _16410_);
  and _68141_ (_16412_, _16261_, _16411_);
  or _68142_ (_16413_, _16412_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _68143_ (_16414_, _16413_, _16397_);
  or _68144_ (_16415_, _16401_, _15132_);
  and _68145_ (_16416_, _16415_, _16414_);
  and _68146_ (_16417_, _16396_, _15140_);
  or _68147_ (_41680_, _16417_, _16416_);
  or _68148_ (_16418_, _16412_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _68149_ (_16419_, _16418_, _16397_);
  or _68150_ (_16420_, _16401_, _15324_);
  and _68151_ (_16421_, _16420_, _16419_);
  and _68152_ (_16422_, _16396_, _15333_);
  or _68153_ (_41681_, _16422_, _16421_);
  or _68154_ (_16423_, _16412_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _68155_ (_16424_, _16423_, _16397_);
  or _68156_ (_16425_, _16401_, _15527_);
  and _68157_ (_16426_, _16425_, _16424_);
  and _68158_ (_16427_, _16396_, _16112_);
  or _68159_ (_41682_, _16427_, _16426_);
  or _68160_ (_16428_, _16412_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _68161_ (_16429_, _16428_, _16397_);
  or _68162_ (_16430_, _16401_, _15724_);
  and _68163_ (_16431_, _16430_, _16429_);
  and _68164_ (_16432_, _16396_, _15733_);
  or _68165_ (_41683_, _16432_, _16431_);
  or _68166_ (_16433_, _16412_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _68167_ (_16434_, _16433_, _16397_);
  or _68168_ (_16435_, _16401_, _15924_);
  and _68169_ (_16436_, _16435_, _16434_);
  and _68170_ (_16437_, _16396_, _15933_);
  or _68171_ (_41684_, _16437_, _16436_);
  nor _68172_ (_16438_, _16399_, _08078_);
  and _68173_ (_16439_, _16399_, _09511_);
  or _68174_ (_16440_, _16439_, _16438_);
  and _68175_ (_16441_, _16440_, _16397_);
  and _68176_ (_16442_, _16396_, _09568_);
  or _68177_ (_41685_, _16442_, _16441_);
  not _68178_ (_16443_, _14555_);
  nor _68179_ (_16444_, _16443_, _07943_);
  not _68180_ (_16445_, _16444_);
  or _68181_ (_16446_, _16445_, _14727_);
  or _68182_ (_16447_, _16444_, \oc8051_golden_model_1.IRAM[12] [0]);
  not _68183_ (_16448_, _07387_);
  or _68184_ (_16449_, _09528_, _16448_);
  and _68185_ (_16450_, _16449_, _16447_);
  and _68186_ (_16451_, _16450_, _16446_);
  and _68187_ (_16452_, _09532_, _07387_);
  and _68188_ (_16453_, _16452_, _14740_);
  or _68189_ (_41689_, _16453_, _16451_);
  not _68190_ (_16454_, _16452_);
  or _68191_ (_16455_, _16444_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _68192_ (_16456_, _16455_, _16454_);
  or _68193_ (_16457_, _16445_, _14929_);
  and _68194_ (_16458_, _16457_, _16456_);
  and _68195_ (_16459_, _16452_, _14938_);
  or _68196_ (_41690_, _16459_, _16458_);
  or _68197_ (_16460_, _16444_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _68198_ (_16461_, _16460_, _16454_);
  or _68199_ (_16462_, _16445_, _15132_);
  and _68200_ (_16463_, _16462_, _16461_);
  and _68201_ (_16464_, _16452_, _15140_);
  or _68202_ (_41691_, _16464_, _16463_);
  or _68203_ (_16465_, _16444_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _68204_ (_16466_, _16465_, _16454_);
  or _68205_ (_16467_, _16445_, _15324_);
  and _68206_ (_16468_, _16467_, _16466_);
  and _68207_ (_16469_, _16452_, _15333_);
  or _68208_ (_41692_, _16469_, _16468_);
  or _68209_ (_16470_, _16444_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _68210_ (_16471_, _16470_, _16454_);
  or _68211_ (_16472_, _16445_, _15527_);
  and _68212_ (_16473_, _16472_, _16471_);
  and _68213_ (_16474_, _16452_, _16112_);
  or _68214_ (_41694_, _16474_, _16473_);
  or _68215_ (_16475_, _16444_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _68216_ (_16476_, _16475_, _16454_);
  or _68217_ (_16477_, _16445_, _15724_);
  and _68218_ (_16478_, _16477_, _16476_);
  and _68219_ (_16479_, _16452_, _15733_);
  or _68220_ (_41695_, _16479_, _16478_);
  or _68221_ (_16480_, _16444_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _68222_ (_16481_, _16480_, _16454_);
  or _68223_ (_16482_, _16445_, _15924_);
  and _68224_ (_16483_, _16482_, _16481_);
  and _68225_ (_16484_, _16452_, _15933_);
  or _68226_ (_41696_, _16484_, _16483_);
  nor _68227_ (_16485_, _16444_, _08097_);
  and _68228_ (_16486_, _16444_, _09511_);
  or _68229_ (_16487_, _16486_, _16485_);
  and _68230_ (_16488_, _16487_, _16449_);
  and _68231_ (_16489_, _16452_, _09568_);
  or _68232_ (_41697_, _16489_, _16488_);
  not _68233_ (_16490_, _07684_);
  or _68234_ (_16491_, _09528_, _16490_);
  or _68235_ (_16492_, _16491_, _14740_);
  not _68236_ (_16493_, _15940_);
  nor _68237_ (_16494_, _16493_, _07943_);
  and _68238_ (_16495_, _16494_, _14727_);
  or _68239_ (_16496_, _16494_, _07242_);
  nand _68240_ (_16497_, _16496_, _16491_);
  or _68241_ (_16498_, _16497_, _16495_);
  and _68242_ (_41700_, _16498_, _16492_);
  and _68243_ (_16499_, _09532_, _07684_);
  not _68244_ (_16500_, _16499_);
  or _68245_ (_16501_, _16494_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _68246_ (_16502_, _16501_, _16500_);
  not _68247_ (_16503_, _16494_);
  or _68248_ (_16504_, _16503_, _14929_);
  and _68249_ (_16505_, _16504_, _16502_);
  and _68250_ (_16506_, _16499_, _14938_);
  or _68251_ (_41701_, _16506_, _16505_);
  or _68252_ (_16507_, _16494_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _68253_ (_16508_, _16507_, _16500_);
  or _68254_ (_16509_, _16503_, _15132_);
  and _68255_ (_16510_, _16509_, _16508_);
  and _68256_ (_16511_, _16499_, _15140_);
  or _68257_ (_41702_, _16511_, _16510_);
  or _68258_ (_16512_, _16494_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _68259_ (_16513_, _16512_, _16500_);
  or _68260_ (_16514_, _16503_, _15324_);
  and _68261_ (_16515_, _16514_, _16513_);
  and _68262_ (_16516_, _16499_, _15333_);
  or _68263_ (_41703_, _16516_, _16515_);
  or _68264_ (_16517_, _16494_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _68265_ (_16518_, _16517_, _16500_);
  or _68266_ (_16519_, _16503_, _15527_);
  and _68267_ (_16520_, _16519_, _16518_);
  and _68268_ (_16521_, _16499_, _16112_);
  or _68269_ (_41705_, _16521_, _16520_);
  or _68270_ (_16522_, _16494_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _68271_ (_16523_, _16522_, _16500_);
  or _68272_ (_16524_, _16503_, _15724_);
  and _68273_ (_16525_, _16524_, _16523_);
  and _68274_ (_16526_, _16499_, _15733_);
  or _68275_ (_41706_, _16526_, _16525_);
  or _68276_ (_16527_, _16494_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _68277_ (_16528_, _16527_, _16500_);
  or _68278_ (_16529_, _16503_, _15924_);
  and _68279_ (_16530_, _16529_, _16528_);
  and _68280_ (_16531_, _16499_, _15933_);
  or _68281_ (_41707_, _16531_, _16530_);
  nor _68282_ (_16532_, _16494_, _08099_);
  and _68283_ (_16533_, _16494_, _09511_);
  or _68284_ (_16534_, _16533_, _16532_);
  and _68285_ (_16535_, _16534_, _16491_);
  and _68286_ (_16536_, _16499_, _09568_);
  or _68287_ (_41708_, _16536_, _16535_);
  not _68288_ (_16537_, _08695_);
  or _68289_ (_16538_, _09528_, _16537_);
  or _68290_ (_16539_, _16538_, _14740_);
  not _68291_ (_16540_, _15989_);
  nor _68292_ (_16541_, _16540_, _07943_);
  and _68293_ (_16542_, _16541_, _14727_);
  or _68294_ (_16543_, _16541_, _07237_);
  nand _68295_ (_16544_, _16543_, _16538_);
  or _68296_ (_16545_, _16544_, _16542_);
  and _68297_ (_41712_, _16545_, _16539_);
  nor _68298_ (_16546_, _16541_, _07436_);
  and _68299_ (_16547_, _16541_, _14929_);
  or _68300_ (_16548_, _16547_, _16546_);
  and _68301_ (_16549_, _16548_, _16538_);
  and _68302_ (_16550_, _09532_, _08695_);
  and _68303_ (_16551_, _16550_, _14938_);
  or _68304_ (_41713_, _16551_, _16549_);
  not _68305_ (_16552_, _16550_);
  or _68306_ (_16553_, _16541_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _68307_ (_16554_, _16553_, _16552_);
  not _68308_ (_16555_, _16541_);
  or _68309_ (_16556_, _16555_, _15132_);
  and _68310_ (_16557_, _16556_, _16554_);
  and _68311_ (_16558_, _16550_, _15140_);
  or _68312_ (_41714_, _16558_, _16557_);
  or _68313_ (_16559_, _16541_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _68314_ (_16560_, _16559_, _16552_);
  or _68315_ (_16561_, _16555_, _15324_);
  and _68316_ (_16562_, _16561_, _16560_);
  and _68317_ (_16563_, _16550_, _15333_);
  or _68318_ (_41716_, _16563_, _16562_);
  or _68319_ (_16564_, _16541_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _68320_ (_16565_, _16564_, _16552_);
  or _68321_ (_16566_, _16555_, _15527_);
  and _68322_ (_16567_, _16566_, _16565_);
  and _68323_ (_16568_, _16550_, _16112_);
  or _68324_ (_41717_, _16568_, _16567_);
  or _68325_ (_16569_, _16541_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _68326_ (_16570_, _16569_, _16552_);
  or _68327_ (_16571_, _16555_, _15724_);
  and _68328_ (_16572_, _16571_, _16570_);
  and _68329_ (_16573_, _16550_, _15733_);
  or _68330_ (_41718_, _16573_, _16572_);
  or _68331_ (_16574_, _16555_, _15924_);
  or _68332_ (_16575_, _16541_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _68333_ (_16576_, _16575_, _16552_);
  and _68334_ (_16577_, _16576_, _16574_);
  and _68335_ (_16578_, _16550_, _15933_);
  or _68336_ (_41719_, _16578_, _16577_);
  nor _68337_ (_16579_, _16541_, _08093_);
  and _68338_ (_16580_, _16541_, _09511_);
  or _68339_ (_16581_, _16580_, _16579_);
  and _68340_ (_16582_, _16581_, _16538_);
  and _68341_ (_16583_, _16550_, _09568_);
  or _68342_ (_41720_, _16583_, _16582_);
  or _68343_ (_16584_, _14740_, _09529_);
  and _68344_ (_16585_, _14727_, _07944_);
  or _68345_ (_16586_, _07944_, _07235_);
  nand _68346_ (_16587_, _16586_, _09529_);
  or _68347_ (_16588_, _16587_, _16585_);
  and _68348_ (_41724_, _16588_, _16584_);
  nor _68349_ (_16589_, _07944_, _07434_);
  and _68350_ (_16590_, _14929_, _07944_);
  or _68351_ (_16591_, _16590_, _16589_);
  and _68352_ (_16592_, _16591_, _09529_);
  and _68353_ (_16593_, _14938_, _09533_);
  or _68354_ (_41725_, _16593_, _16592_);
  not _68355_ (_16594_, _09533_);
  or _68356_ (_16595_, _07944_, \oc8051_golden_model_1.IRAM[15] [2]);
  and _68357_ (_16596_, _16595_, _16594_);
  not _68358_ (_16597_, _07944_);
  or _68359_ (_16598_, _15132_, _16597_);
  and _68360_ (_16599_, _16598_, _16596_);
  and _68361_ (_16600_, _15140_, _09533_);
  or _68362_ (_41726_, _16600_, _16599_);
  or _68363_ (_16601_, _15324_, _16597_);
  or _68364_ (_16602_, _07944_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _68365_ (_16603_, _16602_, _16594_);
  and _68366_ (_16604_, _16603_, _16601_);
  and _68367_ (_16605_, _15333_, _09533_);
  or _68368_ (_41728_, _16605_, _16604_);
  or _68369_ (_16606_, _07944_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _68370_ (_16607_, _16606_, _16594_);
  or _68371_ (_16608_, _15527_, _16597_);
  and _68372_ (_16609_, _16608_, _16607_);
  and _68373_ (_16610_, _16112_, _09533_);
  or _68374_ (_41729_, _16610_, _16609_);
  or _68375_ (_16611_, _15724_, _16597_);
  or _68376_ (_16612_, _07944_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _68377_ (_16613_, _16612_, _16594_);
  and _68378_ (_16614_, _16613_, _16611_);
  and _68379_ (_16615_, _15733_, _09533_);
  or _68380_ (_41730_, _16615_, _16614_);
  or _68381_ (_16616_, _07944_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _68382_ (_16617_, _16616_, _16594_);
  or _68383_ (_16618_, _15924_, _16597_);
  and _68384_ (_16619_, _16618_, _16617_);
  and _68385_ (_16620_, _15933_, _09533_);
  or _68386_ (_41731_, _16620_, _16619_);
  nor _68387_ (_16621_, _01442_, _10179_);
  nor _68388_ (_16622_, _08025_, _10179_);
  and _68389_ (_16623_, _08025_, _09008_);
  or _68390_ (_16624_, _16623_, _16622_);
  or _68391_ (_16625_, _16624_, _06278_);
  and _68392_ (_16626_, _08025_, _07250_);
  or _68393_ (_16627_, _16626_, _16622_);
  or _68394_ (_16628_, _16627_, _06327_);
  or _68395_ (_16629_, _16627_, _06772_);
  nor _68396_ (_16630_, _08453_, _09574_);
  or _68397_ (_16631_, _16630_, _16622_);
  or _68398_ (_16632_, _16631_, _07275_);
  and _68399_ (_16633_, _08025_, \oc8051_golden_model_1.ACC [0]);
  or _68400_ (_16634_, _16633_, _16622_);
  and _68401_ (_16635_, _16634_, _07259_);
  nor _68402_ (_16636_, _07259_, _10179_);
  or _68403_ (_16637_, _16636_, _06474_);
  or _68404_ (_16638_, _16637_, _16635_);
  and _68405_ (_16639_, _16638_, _06357_);
  and _68406_ (_16640_, _16639_, _16632_);
  nor _68407_ (_16641_, _08637_, _10179_);
  and _68408_ (_16642_, _14581_, _08637_);
  or _68409_ (_16643_, _16642_, _16641_);
  and _68410_ (_16644_, _16643_, _06356_);
  or _68411_ (_16645_, _16644_, _16640_);
  or _68412_ (_16646_, _16645_, _06410_);
  and _68413_ (_16647_, _16646_, _16629_);
  or _68414_ (_16648_, _16647_, _06417_);
  or _68415_ (_16649_, _16634_, _06426_);
  and _68416_ (_16650_, _16649_, _06353_);
  and _68417_ (_16651_, _16650_, _16648_);
  and _68418_ (_16652_, _16622_, _06352_);
  or _68419_ (_16653_, _16652_, _06345_);
  or _68420_ (_16654_, _16653_, _16651_);
  or _68421_ (_16655_, _16631_, _06346_);
  and _68422_ (_16656_, _16655_, _16654_);
  or _68423_ (_16657_, _16656_, _09606_);
  nor _68424_ (_16658_, _10115_, _10113_);
  nor _68425_ (_16659_, _16658_, _10116_);
  or _68426_ (_16660_, _16659_, _09612_);
  and _68427_ (_16661_, _16660_, _06340_);
  and _68428_ (_16662_, _16661_, _16657_);
  nand _68429_ (_16663_, _07967_, _10967_);
  or _68430_ (_16664_, _16641_, _16663_);
  and _68431_ (_16665_, _16664_, _06339_);
  and _68432_ (_16666_, _16665_, _16643_);
  or _68433_ (_16667_, _16666_, _10153_);
  or _68434_ (_16668_, _16667_, _16662_);
  and _68435_ (_16669_, _16668_, _16628_);
  or _68436_ (_16670_, _16669_, _09572_);
  and _68437_ (_16671_, _09447_, _08025_);
  not _68438_ (_16672_, _14025_);
  or _68439_ (_16673_, _16622_, _16672_);
  or _68440_ (_16674_, _16673_, _16671_);
  and _68441_ (_16675_, _16674_, _16670_);
  or _68442_ (_16676_, _16675_, _06037_);
  and _68443_ (_16677_, _14666_, _08025_);
  or _68444_ (_16678_, _16622_, _06313_);
  or _68445_ (_16679_, _16678_, _16677_);
  and _68446_ (_16680_, _16679_, _10172_);
  and _68447_ (_16681_, _16680_, _16676_);
  nand _68448_ (_16682_, _10511_, _06071_);
  or _68449_ (_16683_, _10505_, _10452_);
  or _68450_ (_16684_, _10511_, _16683_);
  and _68451_ (_16685_, _16684_, _10166_);
  and _68452_ (_16686_, _16685_, _16682_);
  or _68453_ (_16687_, _16686_, _06277_);
  or _68454_ (_16688_, _16687_, _16681_);
  and _68455_ (_16689_, _16688_, _16625_);
  or _68456_ (_16690_, _16689_, _06502_);
  and _68457_ (_16691_, _14566_, _08025_);
  or _68458_ (_16692_, _16622_, _07334_);
  or _68459_ (_16693_, _16692_, _16691_);
  and _68460_ (_16694_, _16693_, _07337_);
  and _68461_ (_16695_, _16694_, _16690_);
  nor _68462_ (_16696_, _12622_, _09574_);
  or _68463_ (_16697_, _16696_, _16622_);
  and _68464_ (_16698_, _16633_, _08453_);
  nor _68465_ (_16699_, _16698_, _07337_);
  and _68466_ (_16700_, _16699_, _16697_);
  or _68467_ (_16701_, _16700_, _16695_);
  and _68468_ (_16702_, _16701_, _07339_);
  nand _68469_ (_16703_, _16624_, _06507_);
  nor _68470_ (_16704_, _16703_, _16630_);
  or _68471_ (_16705_, _16704_, _06610_);
  or _68472_ (_16706_, _16705_, _16702_);
  or _68473_ (_16707_, _16698_, _16622_);
  or _68474_ (_16708_, _16707_, _07331_);
  and _68475_ (_16709_, _16708_, _16706_);
  or _68476_ (_16710_, _16709_, _06509_);
  and _68477_ (_16711_, _14563_, _08025_);
  or _68478_ (_16712_, _16622_, _09107_);
  or _68479_ (_16713_, _16712_, _16711_);
  and _68480_ (_16714_, _16713_, _09112_);
  and _68481_ (_16715_, _16714_, _16710_);
  and _68482_ (_16716_, _16697_, _06602_);
  or _68483_ (_16717_, _16716_, _06639_);
  or _68484_ (_16718_, _16717_, _16715_);
  or _68485_ (_16719_, _16631_, _07048_);
  and _68486_ (_16720_, _16719_, _16718_);
  or _68487_ (_16721_, _16720_, _05989_);
  or _68488_ (_16722_, _16622_, _05990_);
  and _68489_ (_16723_, _16722_, _16721_);
  or _68490_ (_16724_, _16723_, _06646_);
  or _68491_ (_16725_, _16631_, _06651_);
  and _68492_ (_16726_, _16725_, _01442_);
  and _68493_ (_16727_, _16726_, _16724_);
  or _68494_ (_16728_, _16727_, _16621_);
  and _68495_ (_44115_, _16728_, _43634_);
  nor _68496_ (_16729_, _01442_, _10173_);
  nor _68497_ (_16730_, _08025_, _10173_);
  nor _68498_ (_16731_, _10578_, _09574_);
  or _68499_ (_16732_, _16731_, _16730_);
  or _68500_ (_16733_, _16732_, _09112_);
  or _68501_ (_16734_, _08025_, \oc8051_golden_model_1.B [1]);
  nand _68502_ (_16735_, _08025_, _07160_);
  and _68503_ (_16736_, _16735_, _06277_);
  and _68504_ (_16737_, _16736_, _16734_);
  nor _68505_ (_16738_, _08637_, _10173_);
  and _68506_ (_16739_, _14767_, _08637_);
  or _68507_ (_16740_, _16739_, _16738_);
  or _68508_ (_16741_, _16738_, _14782_);
  and _68509_ (_16742_, _16741_, _16740_);
  or _68510_ (_16743_, _16742_, _06346_);
  nor _68511_ (_16744_, _09574_, _07448_);
  or _68512_ (_16745_, _16744_, _16730_);
  and _68513_ (_16746_, _16745_, _06410_);
  or _68514_ (_16747_, _16740_, _06357_);
  and _68515_ (_16748_, _14744_, _08025_);
  not _68516_ (_16749_, _16748_);
  and _68517_ (_16750_, _16749_, _16734_);
  and _68518_ (_16751_, _16750_, _06474_);
  nor _68519_ (_16752_, _07259_, _10173_);
  and _68520_ (_16753_, _08025_, \oc8051_golden_model_1.ACC [1]);
  or _68521_ (_16754_, _16753_, _16730_);
  and _68522_ (_16755_, _16754_, _07259_);
  or _68523_ (_16756_, _16755_, _16752_);
  and _68524_ (_16757_, _16756_, _07275_);
  or _68525_ (_16758_, _16757_, _06356_);
  or _68526_ (_16759_, _16758_, _16751_);
  and _68527_ (_16760_, _16759_, _16747_);
  and _68528_ (_16761_, _16760_, _06772_);
  or _68529_ (_16762_, _16761_, _16746_);
  or _68530_ (_16763_, _16762_, _06417_);
  or _68531_ (_16764_, _16754_, _06426_);
  and _68532_ (_16765_, _16764_, _06353_);
  and _68533_ (_16766_, _16765_, _16763_);
  and _68534_ (_16767_, _14754_, _08637_);
  or _68535_ (_16768_, _16767_, _16738_);
  and _68536_ (_16769_, _16768_, _06352_);
  or _68537_ (_16770_, _16769_, _06345_);
  or _68538_ (_16771_, _16770_, _16766_);
  and _68539_ (_16772_, _16771_, _16743_);
  or _68540_ (_16773_, _16772_, _09606_);
  nor _68541_ (_16774_, _10118_, _10060_);
  nor _68542_ (_16775_, _16774_, _10119_);
  or _68543_ (_16776_, _16775_, _09612_);
  and _68544_ (_16777_, _16776_, _06340_);
  and _68545_ (_16778_, _16777_, _16773_);
  and _68546_ (_16779_, _14796_, _08637_);
  or _68547_ (_16780_, _16779_, _16738_);
  and _68548_ (_16781_, _16780_, _06339_);
  or _68549_ (_16782_, _16781_, _10153_);
  or _68550_ (_16783_, _16782_, _16778_);
  or _68551_ (_16784_, _16745_, _06327_);
  and _68552_ (_16785_, _16784_, _16783_);
  or _68553_ (_16786_, _16785_, _09572_);
  and _68554_ (_16787_, _09402_, _08025_);
  or _68555_ (_16788_, _16730_, _06333_);
  or _68556_ (_16789_, _16788_, _16787_);
  and _68557_ (_16790_, _16789_, _06313_);
  and _68558_ (_16791_, _16790_, _16786_);
  or _68559_ (_16792_, _14851_, _09574_);
  and _68560_ (_16793_, _16734_, _06037_);
  and _68561_ (_16794_, _16793_, _16792_);
  or _68562_ (_16795_, _16794_, _10166_);
  or _68563_ (_16796_, _16795_, _16791_);
  nor _68564_ (_16797_, _10506_, _10504_);
  or _68565_ (_16798_, _16797_, _10507_);
  nor _68566_ (_16799_, _16798_, _10511_);
  and _68567_ (_16800_, _10511_, _10449_);
  or _68568_ (_16801_, _16800_, _16799_);
  or _68569_ (_16802_, _16801_, _10172_);
  and _68570_ (_16803_, _16802_, _06278_);
  and _68571_ (_16804_, _16803_, _16796_);
  or _68572_ (_16805_, _16804_, _16737_);
  and _68573_ (_16806_, _16805_, _07334_);
  or _68574_ (_16807_, _14749_, _09574_);
  and _68575_ (_16808_, _16734_, _06502_);
  and _68576_ (_16809_, _16808_, _16807_);
  or _68577_ (_16810_, _16809_, _06615_);
  or _68578_ (_16811_, _16810_, _16806_);
  and _68579_ (_16812_, _10579_, _08025_);
  or _68580_ (_16813_, _16812_, _16730_);
  or _68581_ (_16814_, _16813_, _07337_);
  and _68582_ (_16815_, _16814_, _07339_);
  and _68583_ (_16816_, _16815_, _16811_);
  or _68584_ (_16817_, _14747_, _09574_);
  and _68585_ (_16818_, _16734_, _06507_);
  and _68586_ (_16819_, _16818_, _16817_);
  or _68587_ (_16820_, _16819_, _06610_);
  or _68588_ (_16821_, _16820_, _16816_);
  and _68589_ (_16822_, _16753_, _08404_);
  or _68590_ (_16823_, _16730_, _07331_);
  or _68591_ (_16824_, _16823_, _16822_);
  and _68592_ (_16825_, _16824_, _09107_);
  and _68593_ (_16826_, _16825_, _16821_);
  or _68594_ (_16827_, _16735_, _08404_);
  and _68595_ (_16828_, _16734_, _06509_);
  and _68596_ (_16829_, _16828_, _16827_);
  or _68597_ (_16830_, _16829_, _06602_);
  or _68598_ (_16831_, _16830_, _16826_);
  and _68599_ (_16832_, _16831_, _16733_);
  or _68600_ (_16833_, _16832_, _06639_);
  or _68601_ (_16834_, _16750_, _07048_);
  and _68602_ (_16835_, _16834_, _05990_);
  and _68603_ (_16836_, _16835_, _16833_);
  and _68604_ (_16837_, _16768_, _05989_);
  or _68605_ (_16838_, _16837_, _06646_);
  or _68606_ (_16839_, _16838_, _16836_);
  or _68607_ (_16840_, _16730_, _06651_);
  or _68608_ (_16841_, _16840_, _16748_);
  and _68609_ (_16842_, _16841_, _01442_);
  and _68610_ (_16843_, _16842_, _16839_);
  or _68611_ (_16844_, _16843_, _16729_);
  and _68612_ (_44116_, _16844_, _43634_);
  nor _68613_ (_16845_, _01442_, _10326_);
  nor _68614_ (_16846_, _08025_, _10326_);
  and _68615_ (_16847_, _08025_, _09057_);
  or _68616_ (_16848_, _16847_, _16846_);
  or _68617_ (_16849_, _16848_, _06278_);
  nor _68618_ (_16850_, _09574_, _07854_);
  or _68619_ (_16851_, _16850_, _16846_);
  or _68620_ (_16852_, _16851_, _06327_);
  nor _68621_ (_16853_, _08637_, _10326_);
  and _68622_ (_16854_, _14955_, _08637_);
  or _68623_ (_16855_, _16854_, _16853_);
  or _68624_ (_16856_, _16853_, _14986_);
  and _68625_ (_16857_, _16856_, _16855_);
  or _68626_ (_16858_, _16857_, _06346_);
  and _68627_ (_16859_, _14959_, _08025_);
  or _68628_ (_16860_, _16859_, _16846_);
  and _68629_ (_16861_, _16860_, _06474_);
  nor _68630_ (_16862_, _07259_, _10326_);
  and _68631_ (_16863_, _08025_, \oc8051_golden_model_1.ACC [2]);
  or _68632_ (_16864_, _16863_, _16846_);
  and _68633_ (_16865_, _16864_, _07259_);
  or _68634_ (_16866_, _16865_, _16862_);
  and _68635_ (_16867_, _16866_, _07275_);
  or _68636_ (_16868_, _16867_, _06356_);
  or _68637_ (_16869_, _16868_, _16861_);
  or _68638_ (_16870_, _16855_, _06357_);
  and _68639_ (_16871_, _16870_, _06772_);
  and _68640_ (_16872_, _16871_, _16869_);
  and _68641_ (_16873_, _16851_, _06410_);
  or _68642_ (_16874_, _16873_, _06417_);
  or _68643_ (_16875_, _16874_, _16872_);
  or _68644_ (_16876_, _16864_, _06426_);
  and _68645_ (_16877_, _16876_, _06353_);
  and _68646_ (_16878_, _16877_, _16875_);
  and _68647_ (_16879_, _14953_, _08637_);
  or _68648_ (_16880_, _16879_, _16853_);
  and _68649_ (_16881_, _16880_, _06352_);
  or _68650_ (_16882_, _16881_, _06345_);
  or _68651_ (_16883_, _16882_, _16878_);
  and _68652_ (_16884_, _16883_, _16858_);
  or _68653_ (_16885_, _16884_, _09606_);
  or _68654_ (_16886_, _10120_, _10015_);
  and _68655_ (_16887_, _16886_, _10121_);
  or _68656_ (_16888_, _16887_, _09612_);
  and _68657_ (_16889_, _16888_, _06340_);
  and _68658_ (_16890_, _16889_, _16885_);
  and _68659_ (_16891_, _15000_, _08637_);
  or _68660_ (_16892_, _16891_, _16853_);
  and _68661_ (_16893_, _16892_, _06339_);
  or _68662_ (_16894_, _16893_, _10153_);
  or _68663_ (_16895_, _16894_, _16890_);
  and _68664_ (_16896_, _16895_, _16852_);
  or _68665_ (_16897_, _16896_, _09572_);
  and _68666_ (_16898_, _09356_, _08025_);
  or _68667_ (_16899_, _16846_, _16672_);
  or _68668_ (_16900_, _16899_, _16898_);
  and _68669_ (_16901_, _16900_, _16897_);
  or _68670_ (_16902_, _16901_, _06037_);
  and _68671_ (_16903_, _15056_, _08025_);
  or _68672_ (_16904_, _16846_, _06313_);
  or _68673_ (_16905_, _16904_, _16903_);
  and _68674_ (_16906_, _16905_, _10172_);
  and _68675_ (_16907_, _16906_, _16902_);
  not _68676_ (_16908_, _10511_);
  or _68677_ (_16909_, _16908_, _10440_);
  nor _68678_ (_16910_, _10507_, _10450_);
  not _68679_ (_16911_, _16910_);
  and _68680_ (_16912_, _16911_, _10443_);
  nor _68681_ (_16913_, _16911_, _10443_);
  nor _68682_ (_16914_, _16913_, _16912_);
  or _68683_ (_16915_, _16914_, _10511_);
  and _68684_ (_16916_, _16915_, _10166_);
  and _68685_ (_16917_, _16916_, _16909_);
  or _68686_ (_16918_, _16917_, _06277_);
  or _68687_ (_16919_, _16918_, _16907_);
  and _68688_ (_16920_, _16919_, _16849_);
  or _68689_ (_16921_, _16920_, _06502_);
  and _68690_ (_16922_, _14948_, _08025_);
  or _68691_ (_16923_, _16846_, _07334_);
  or _68692_ (_16924_, _16923_, _16922_);
  and _68693_ (_16925_, _16924_, _07337_);
  and _68694_ (_16926_, _16925_, _16921_);
  and _68695_ (_16927_, _10583_, _08025_);
  or _68696_ (_16928_, _16927_, _16846_);
  and _68697_ (_16929_, _16928_, _06615_);
  or _68698_ (_16930_, _16929_, _16926_);
  and _68699_ (_16931_, _16930_, _07339_);
  or _68700_ (_16932_, _16846_, _08503_);
  and _68701_ (_16933_, _16848_, _06507_);
  and _68702_ (_16934_, _16933_, _16932_);
  or _68703_ (_16935_, _16934_, _16931_);
  and _68704_ (_16936_, _16935_, _07331_);
  and _68705_ (_16937_, _16864_, _06610_);
  and _68706_ (_16938_, _16937_, _16932_);
  or _68707_ (_16939_, _16938_, _06509_);
  or _68708_ (_16940_, _16939_, _16936_);
  and _68709_ (_16941_, _14945_, _08025_);
  or _68710_ (_16942_, _16846_, _09107_);
  or _68711_ (_16943_, _16942_, _16941_);
  and _68712_ (_16944_, _16943_, _09112_);
  and _68713_ (_16945_, _16944_, _16940_);
  nor _68714_ (_16946_, _10582_, _09574_);
  or _68715_ (_16947_, _16946_, _16846_);
  and _68716_ (_16948_, _16947_, _06602_);
  or _68717_ (_16949_, _16948_, _06639_);
  or _68718_ (_16950_, _16949_, _16945_);
  or _68719_ (_16951_, _16860_, _07048_);
  and _68720_ (_16952_, _16951_, _05990_);
  and _68721_ (_16953_, _16952_, _16950_);
  and _68722_ (_16954_, _16880_, _05989_);
  or _68723_ (_16955_, _16954_, _06646_);
  or _68724_ (_16956_, _16955_, _16953_);
  and _68725_ (_16957_, _15129_, _08025_);
  or _68726_ (_16958_, _16846_, _06651_);
  or _68727_ (_16959_, _16958_, _16957_);
  and _68728_ (_16960_, _16959_, _01442_);
  and _68729_ (_16961_, _16960_, _16956_);
  or _68730_ (_16962_, _16961_, _16845_);
  and _68731_ (_44117_, _16962_, _43634_);
  nor _68732_ (_16963_, _01442_, _10215_);
  nor _68733_ (_16964_, _08025_, _10215_);
  nor _68734_ (_16965_, _10574_, _09574_);
  or _68735_ (_16966_, _16965_, _16964_);
  and _68736_ (_16967_, _08025_, \oc8051_golden_model_1.ACC [3]);
  nand _68737_ (_16968_, _16967_, _08359_);
  and _68738_ (_16969_, _16968_, _06615_);
  and _68739_ (_16970_, _16969_, _16966_);
  and _68740_ (_16971_, _08025_, _09014_);
  or _68741_ (_16972_, _16971_, _16964_);
  or _68742_ (_16973_, _16972_, _06278_);
  and _68743_ (_16974_, _15251_, _08025_);
  or _68744_ (_16975_, _16974_, _16964_);
  and _68745_ (_16976_, _16975_, _06037_);
  nor _68746_ (_16977_, _08637_, _10215_);
  and _68747_ (_16978_, _15150_, _08637_);
  or _68748_ (_16979_, _16978_, _16977_);
  or _68749_ (_16980_, _16977_, _15180_);
  and _68750_ (_16981_, _16980_, _16979_);
  or _68751_ (_16982_, _16981_, _06346_);
  and _68752_ (_16983_, _15153_, _08025_);
  or _68753_ (_16984_, _16983_, _16964_);
  or _68754_ (_16985_, _16984_, _07275_);
  or _68755_ (_16986_, _16967_, _16964_);
  and _68756_ (_16987_, _16986_, _07259_);
  nor _68757_ (_16988_, _07259_, _10215_);
  or _68758_ (_16989_, _16988_, _06474_);
  or _68759_ (_16990_, _16989_, _16987_);
  and _68760_ (_16991_, _16990_, _06357_);
  and _68761_ (_16992_, _16991_, _16985_);
  and _68762_ (_16993_, _16979_, _06356_);
  or _68763_ (_16994_, _16993_, _06410_);
  or _68764_ (_16995_, _16994_, _16992_);
  nor _68765_ (_16996_, _09574_, _07680_);
  or _68766_ (_16997_, _16996_, _16964_);
  or _68767_ (_16998_, _16997_, _06772_);
  and _68768_ (_16999_, _16998_, _16995_);
  or _68769_ (_17000_, _16999_, _06417_);
  or _68770_ (_17001_, _16986_, _06426_);
  and _68771_ (_17002_, _17001_, _06353_);
  and _68772_ (_17003_, _17002_, _17000_);
  and _68773_ (_17004_, _15148_, _08637_);
  or _68774_ (_17005_, _17004_, _16977_);
  and _68775_ (_17006_, _17005_, _06352_);
  or _68776_ (_17007_, _17006_, _06345_);
  or _68777_ (_17008_, _17007_, _17003_);
  and _68778_ (_17009_, _17008_, _16982_);
  or _68779_ (_17010_, _17009_, _09606_);
  nor _68780_ (_17011_, _10123_, _09957_);
  nor _68781_ (_17012_, _17011_, _10124_);
  or _68782_ (_17013_, _17012_, _09612_);
  and _68783_ (_17014_, _17013_, _06340_);
  and _68784_ (_17015_, _17014_, _17010_);
  and _68785_ (_17016_, _15197_, _08637_);
  or _68786_ (_17017_, _17016_, _16977_);
  and _68787_ (_17018_, _17017_, _06339_);
  or _68788_ (_17019_, _17018_, _10153_);
  or _68789_ (_17020_, _17019_, _17015_);
  or _68790_ (_17021_, _16997_, _06327_);
  and _68791_ (_17022_, _17021_, _17020_);
  or _68792_ (_17023_, _17022_, _09572_);
  and _68793_ (_17024_, _09310_, _08025_);
  or _68794_ (_17025_, _16964_, _06333_);
  or _68795_ (_17026_, _17025_, _17024_);
  and _68796_ (_17027_, _17026_, _06313_);
  and _68797_ (_17028_, _17027_, _17023_);
  or _68798_ (_17029_, _17028_, _16976_);
  and _68799_ (_17030_, _17029_, _10172_);
  nor _68800_ (_17031_, _16912_, _10442_);
  nor _68801_ (_17032_, _17031_, _10434_);
  and _68802_ (_17033_, _17031_, _10434_);
  or _68803_ (_17034_, _17033_, _17032_);
  or _68804_ (_17035_, _17034_, _10511_);
  or _68805_ (_17036_, _16908_, _10431_);
  and _68806_ (_17037_, _17036_, _10166_);
  and _68807_ (_17038_, _17037_, _17035_);
  or _68808_ (_17039_, _17038_, _06277_);
  or _68809_ (_17040_, _17039_, _17030_);
  and _68810_ (_17041_, _17040_, _16973_);
  or _68811_ (_17042_, _17041_, _06502_);
  and _68812_ (_17043_, _15266_, _08025_);
  or _68813_ (_17044_, _16964_, _07334_);
  or _68814_ (_17045_, _17044_, _17043_);
  and _68815_ (_17046_, _17045_, _07337_);
  and _68816_ (_17047_, _17046_, _17042_);
  or _68817_ (_17048_, _17047_, _16970_);
  and _68818_ (_17049_, _17048_, _07339_);
  or _68819_ (_17050_, _16964_, _08359_);
  and _68820_ (_17051_, _16972_, _06507_);
  and _68821_ (_17052_, _17051_, _17050_);
  or _68822_ (_17053_, _17052_, _17049_);
  and _68823_ (_17054_, _17053_, _07331_);
  and _68824_ (_17055_, _16986_, _06610_);
  and _68825_ (_17056_, _17055_, _17050_);
  or _68826_ (_17057_, _17056_, _06509_);
  or _68827_ (_17058_, _17057_, _17054_);
  and _68828_ (_17059_, _15263_, _08025_);
  or _68829_ (_17060_, _16964_, _09107_);
  or _68830_ (_17061_, _17060_, _17059_);
  and _68831_ (_17062_, _17061_, _09112_);
  and _68832_ (_17063_, _17062_, _17058_);
  and _68833_ (_17064_, _16966_, _06602_);
  or _68834_ (_17065_, _17064_, _06639_);
  or _68835_ (_17066_, _17065_, _17063_);
  or _68836_ (_17067_, _16984_, _07048_);
  and _68837_ (_17068_, _17067_, _05990_);
  and _68838_ (_17069_, _17068_, _17066_);
  and _68839_ (_17070_, _17005_, _05989_);
  or _68840_ (_17071_, _17070_, _06646_);
  or _68841_ (_17072_, _17071_, _17069_);
  and _68842_ (_17073_, _15321_, _08025_);
  or _68843_ (_17074_, _16964_, _06651_);
  or _68844_ (_17075_, _17074_, _17073_);
  and _68845_ (_17076_, _17075_, _01442_);
  and _68846_ (_17077_, _17076_, _17072_);
  or _68847_ (_17078_, _17077_, _16963_);
  and _68848_ (_44118_, _17078_, _43634_);
  nor _68849_ (_17079_, _01442_, _10305_);
  nor _68850_ (_17080_, _08025_, _10305_);
  nor _68851_ (_17081_, _10589_, _09574_);
  or _68852_ (_17082_, _17081_, _17080_);
  and _68853_ (_17083_, _08025_, \oc8051_golden_model_1.ACC [4]);
  nand _68854_ (_17084_, _17083_, _08599_);
  and _68855_ (_17085_, _17084_, _06615_);
  and _68856_ (_17086_, _17085_, _17082_);
  and _68857_ (_17087_, _08995_, _08025_);
  or _68858_ (_17088_, _17087_, _17080_);
  or _68859_ (_17089_, _17088_, _06278_);
  and _68860_ (_17090_, _15452_, _08025_);
  or _68861_ (_17091_, _17090_, _17080_);
  and _68862_ (_17092_, _17091_, _06037_);
  nor _68863_ (_17093_, _08596_, _09574_);
  or _68864_ (_17094_, _17093_, _17080_);
  or _68865_ (_17095_, _17094_, _06327_);
  nor _68866_ (_17096_, _08637_, _10305_);
  and _68867_ (_17097_, _15348_, _08637_);
  or _68868_ (_17098_, _17097_, _17096_);
  and _68869_ (_17099_, _17098_, _06352_);
  and _68870_ (_17100_, _15367_, _08025_);
  or _68871_ (_17101_, _17100_, _17080_);
  or _68872_ (_17102_, _17101_, _07275_);
  or _68873_ (_17103_, _17083_, _17080_);
  and _68874_ (_17104_, _17103_, _07259_);
  nor _68875_ (_17105_, _07259_, _10305_);
  or _68876_ (_17106_, _17105_, _06474_);
  or _68877_ (_17107_, _17106_, _17104_);
  and _68878_ (_17108_, _17107_, _06357_);
  and _68879_ (_17109_, _17108_, _17102_);
  and _68880_ (_17110_, _15353_, _08637_);
  or _68881_ (_17111_, _17110_, _17096_);
  and _68882_ (_17112_, _17111_, _06356_);
  or _68883_ (_17113_, _17112_, _06410_);
  or _68884_ (_17114_, _17113_, _17109_);
  or _68885_ (_17115_, _17094_, _06772_);
  and _68886_ (_17116_, _17115_, _17114_);
  or _68887_ (_17117_, _17116_, _06417_);
  or _68888_ (_17118_, _17103_, _06426_);
  and _68889_ (_17119_, _17118_, _06353_);
  and _68890_ (_17120_, _17119_, _17117_);
  or _68891_ (_17121_, _17120_, _17099_);
  and _68892_ (_17122_, _17121_, _06346_);
  or _68893_ (_17123_, _17096_, _15384_);
  and _68894_ (_17124_, _17111_, _06345_);
  and _68895_ (_17125_, _17124_, _17123_);
  or _68896_ (_17126_, _17125_, _09606_);
  or _68897_ (_17127_, _17126_, _17122_);
  or _68898_ (_17128_, _10127_, _10125_);
  and _68899_ (_17129_, _17128_, _10128_);
  or _68900_ (_17130_, _17129_, _09612_);
  and _68901_ (_17131_, _17130_, _06340_);
  and _68902_ (_17132_, _17131_, _17127_);
  and _68903_ (_17133_, _15350_, _08637_);
  or _68904_ (_17134_, _17133_, _17096_);
  and _68905_ (_17135_, _17134_, _06339_);
  or _68906_ (_17136_, _17135_, _10153_);
  or _68907_ (_17137_, _17136_, _17132_);
  and _68908_ (_17138_, _17137_, _17095_);
  or _68909_ (_17139_, _17138_, _09572_);
  and _68910_ (_17140_, _09264_, _08025_);
  or _68911_ (_17141_, _17080_, _06333_);
  or _68912_ (_17142_, _17141_, _17140_);
  and _68913_ (_17143_, _17142_, _06313_);
  and _68914_ (_17144_, _17143_, _17139_);
  or _68915_ (_17145_, _17144_, _17092_);
  and _68916_ (_17146_, _17145_, _10172_);
  or _68917_ (_17147_, _16908_, _10465_);
  nor _68918_ (_17148_, _17031_, _10433_);
  or _68919_ (_17149_, _17148_, _10432_);
  nand _68920_ (_17150_, _17149_, _10468_);
  or _68921_ (_17151_, _17149_, _10468_);
  and _68922_ (_17152_, _17151_, _17150_);
  or _68923_ (_17153_, _17152_, _10511_);
  and _68924_ (_17154_, _17153_, _10166_);
  and _68925_ (_17155_, _17154_, _17147_);
  or _68926_ (_17156_, _17155_, _06277_);
  or _68927_ (_17157_, _17156_, _17146_);
  and _68928_ (_17158_, _17157_, _17089_);
  or _68929_ (_17159_, _17158_, _06502_);
  and _68930_ (_17160_, _15345_, _08025_);
  or _68931_ (_17161_, _17080_, _07334_);
  or _68932_ (_17162_, _17161_, _17160_);
  and _68933_ (_17163_, _17162_, _07337_);
  and _68934_ (_17164_, _17163_, _17159_);
  or _68935_ (_17165_, _17164_, _17086_);
  and _68936_ (_17166_, _17165_, _07339_);
  or _68937_ (_17167_, _17080_, _08599_);
  and _68938_ (_17168_, _17088_, _06507_);
  and _68939_ (_17169_, _17168_, _17167_);
  or _68940_ (_17170_, _17169_, _17166_);
  and _68941_ (_17171_, _17170_, _07331_);
  and _68942_ (_17172_, _17103_, _06610_);
  and _68943_ (_17173_, _17172_, _17167_);
  or _68944_ (_17174_, _17173_, _06509_);
  or _68945_ (_17175_, _17174_, _17171_);
  and _68946_ (_17176_, _15342_, _08025_);
  or _68947_ (_17177_, _17080_, _09107_);
  or _68948_ (_17178_, _17177_, _17176_);
  and _68949_ (_17179_, _17178_, _09112_);
  and _68950_ (_17180_, _17179_, _17175_);
  and _68951_ (_17181_, _17082_, _06602_);
  or _68952_ (_17182_, _17181_, _06639_);
  or _68953_ (_17183_, _17182_, _17180_);
  or _68954_ (_17184_, _17101_, _07048_);
  and _68955_ (_17185_, _17184_, _05990_);
  and _68956_ (_17186_, _17185_, _17183_);
  and _68957_ (_17187_, _17098_, _05989_);
  or _68958_ (_17188_, _17187_, _06646_);
  or _68959_ (_17189_, _17188_, _17186_);
  and _68960_ (_17190_, _15524_, _08025_);
  or _68961_ (_17191_, _17080_, _06651_);
  or _68962_ (_17192_, _17191_, _17190_);
  and _68963_ (_17193_, _17192_, _01442_);
  and _68964_ (_17194_, _17193_, _17189_);
  or _68965_ (_17195_, _17194_, _17079_);
  and _68966_ (_44119_, _17195_, _43634_);
  nor _68967_ (_17196_, _01442_, _10296_);
  nor _68968_ (_17197_, _08025_, _10296_);
  and _68969_ (_17198_, _15649_, _08025_);
  or _68970_ (_17199_, _17198_, _17197_);
  and _68971_ (_17200_, _17199_, _06037_);
  nor _68972_ (_17201_, _08305_, _09574_);
  or _68973_ (_17202_, _17201_, _17197_);
  or _68974_ (_17203_, _17202_, _06327_);
  nor _68975_ (_17204_, _08637_, _10296_);
  and _68976_ (_17205_, _15544_, _08637_);
  or _68977_ (_17206_, _17205_, _17204_);
  and _68978_ (_17207_, _17206_, _06352_);
  and _68979_ (_17208_, _15550_, _08025_);
  or _68980_ (_17209_, _17208_, _17197_);
  or _68981_ (_17210_, _17209_, _07275_);
  and _68982_ (_17211_, _08025_, \oc8051_golden_model_1.ACC [5]);
  or _68983_ (_17212_, _17211_, _17197_);
  and _68984_ (_17213_, _17212_, _07259_);
  nor _68985_ (_17214_, _07259_, _10296_);
  or _68986_ (_17215_, _17214_, _06474_);
  or _68987_ (_17216_, _17215_, _17213_);
  and _68988_ (_17217_, _17216_, _06357_);
  and _68989_ (_17218_, _17217_, _17210_);
  and _68990_ (_17219_, _15566_, _08637_);
  or _68991_ (_17220_, _17219_, _17204_);
  and _68992_ (_17221_, _17220_, _06356_);
  or _68993_ (_17222_, _17221_, _06410_);
  or _68994_ (_17223_, _17222_, _17218_);
  or _68995_ (_17224_, _17202_, _06772_);
  and _68996_ (_17225_, _17224_, _17223_);
  or _68997_ (_17226_, _17225_, _06417_);
  or _68998_ (_17227_, _17212_, _06426_);
  and _68999_ (_17228_, _17227_, _06353_);
  and _69000_ (_17229_, _17228_, _17226_);
  or _69001_ (_17230_, _17229_, _17207_);
  and _69002_ (_17231_, _17230_, _06346_);
  or _69003_ (_17232_, _17204_, _15581_);
  and _69004_ (_17233_, _17220_, _06345_);
  and _69005_ (_17234_, _17233_, _17232_);
  or _69006_ (_17235_, _17234_, _09606_);
  or _69007_ (_17236_, _17235_, _17231_);
  nor _69008_ (_17237_, _10130_, _09831_);
  nor _69009_ (_17238_, _17237_, _10131_);
  or _69010_ (_17239_, _17238_, _09612_);
  and _69011_ (_17240_, _17239_, _06340_);
  and _69012_ (_17241_, _17240_, _17236_);
  and _69013_ (_17242_, _15546_, _08637_);
  or _69014_ (_17243_, _17242_, _17204_);
  and _69015_ (_17244_, _17243_, _06339_);
  or _69016_ (_17245_, _17244_, _10153_);
  or _69017_ (_17246_, _17245_, _17241_);
  and _69018_ (_17247_, _17246_, _17203_);
  or _69019_ (_17248_, _17247_, _09572_);
  and _69020_ (_17249_, _09218_, _08025_);
  or _69021_ (_17250_, _17197_, _06333_);
  or _69022_ (_17251_, _17250_, _17249_);
  and _69023_ (_17252_, _17251_, _06313_);
  and _69024_ (_17253_, _17252_, _17248_);
  or _69025_ (_17254_, _17253_, _17200_);
  and _69026_ (_17255_, _17254_, _10172_);
  or _69027_ (_17256_, _16908_, _10475_);
  not _69028_ (_17257_, _10467_);
  and _69029_ (_17258_, _17150_, _17257_);
  nor _69030_ (_17259_, _17258_, _10478_);
  and _69031_ (_17260_, _17258_, _10478_);
  or _69032_ (_17261_, _17260_, _17259_);
  or _69033_ (_17262_, _17261_, _10511_);
  and _69034_ (_17263_, _17262_, _10166_);
  and _69035_ (_17264_, _17263_, _17256_);
  or _69036_ (_17265_, _17264_, _06277_);
  or _69037_ (_17266_, _17265_, _17255_);
  and _69038_ (_17267_, _08954_, _08025_);
  or _69039_ (_17268_, _17267_, _17197_);
  or _69040_ (_17269_, _17268_, _06278_);
  and _69041_ (_17270_, _17269_, _17266_);
  or _69042_ (_17271_, _17270_, _06502_);
  and _69043_ (_17272_, _15664_, _08025_);
  or _69044_ (_17273_, _17197_, _07334_);
  or _69045_ (_17274_, _17273_, _17272_);
  and _69046_ (_17275_, _17274_, _07337_);
  and _69047_ (_17276_, _17275_, _17271_);
  and _69048_ (_17277_, _12626_, _08025_);
  or _69049_ (_17278_, _17277_, _17197_);
  and _69050_ (_17279_, _17278_, _06615_);
  or _69051_ (_17280_, _17279_, _17276_);
  and _69052_ (_17281_, _17280_, _07339_);
  or _69053_ (_17282_, _17197_, _08308_);
  and _69054_ (_17283_, _17268_, _06507_);
  and _69055_ (_17284_, _17283_, _17282_);
  or _69056_ (_17285_, _17284_, _17281_);
  and _69057_ (_17286_, _17285_, _07331_);
  and _69058_ (_17287_, _17212_, _06610_);
  and _69059_ (_17288_, _17287_, _17282_);
  or _69060_ (_17289_, _17288_, _06509_);
  or _69061_ (_17290_, _17289_, _17286_);
  and _69062_ (_17291_, _15663_, _08025_);
  or _69063_ (_17292_, _17197_, _09107_);
  or _69064_ (_17293_, _17292_, _17291_);
  and _69065_ (_17294_, _17293_, _09112_);
  and _69066_ (_17295_, _17294_, _17290_);
  nor _69067_ (_17296_, _10570_, _09574_);
  or _69068_ (_17297_, _17296_, _17197_);
  and _69069_ (_17298_, _17297_, _06602_);
  or _69070_ (_17299_, _17298_, _06639_);
  or _69071_ (_17300_, _17299_, _17295_);
  or _69072_ (_17301_, _17209_, _07048_);
  and _69073_ (_17302_, _17301_, _05990_);
  and _69074_ (_17303_, _17302_, _17300_);
  and _69075_ (_17304_, _17206_, _05989_);
  or _69076_ (_17305_, _17304_, _06646_);
  or _69077_ (_17306_, _17305_, _17303_);
  and _69078_ (_17307_, _15721_, _08025_);
  or _69079_ (_17308_, _17197_, _06651_);
  or _69080_ (_17309_, _17308_, _17307_);
  and _69081_ (_17310_, _17309_, _01442_);
  and _69082_ (_17311_, _17310_, _17306_);
  or _69083_ (_17312_, _17311_, _17196_);
  and _69084_ (_44121_, _17312_, _43634_);
  nor _69085_ (_17313_, _01442_, _10483_);
  nor _69086_ (_17314_, _08025_, _10483_);
  and _69087_ (_17315_, _15853_, _08025_);
  or _69088_ (_17316_, _17315_, _17314_);
  or _69089_ (_17317_, _17316_, _06278_);
  and _69090_ (_17318_, _15846_, _08025_);
  or _69091_ (_17319_, _17318_, _17314_);
  and _69092_ (_17320_, _17319_, _06037_);
  nor _69093_ (_17321_, _08209_, _09574_);
  or _69094_ (_17322_, _17321_, _17314_);
  or _69095_ (_17323_, _17322_, _06327_);
  nor _69096_ (_17324_, _08637_, _10483_);
  and _69097_ (_17325_, _15743_, _08637_);
  or _69098_ (_17326_, _17325_, _17324_);
  and _69099_ (_17327_, _17326_, _06352_);
  and _69100_ (_17328_, _15759_, _08025_);
  or _69101_ (_17329_, _17328_, _17314_);
  or _69102_ (_17330_, _17329_, _07275_);
  and _69103_ (_17331_, _08025_, \oc8051_golden_model_1.ACC [6]);
  or _69104_ (_17332_, _17331_, _17314_);
  and _69105_ (_17333_, _17332_, _07259_);
  nor _69106_ (_17334_, _07259_, _10483_);
  or _69107_ (_17335_, _17334_, _06474_);
  or _69108_ (_17336_, _17335_, _17333_);
  and _69109_ (_17337_, _17336_, _06357_);
  and _69110_ (_17338_, _17337_, _17330_);
  and _69111_ (_17339_, _15763_, _08637_);
  or _69112_ (_17340_, _17339_, _17324_);
  and _69113_ (_17341_, _17340_, _06356_);
  or _69114_ (_17342_, _17341_, _06410_);
  or _69115_ (_17343_, _17342_, _17338_);
  or _69116_ (_17344_, _17322_, _06772_);
  and _69117_ (_17345_, _17344_, _17343_);
  or _69118_ (_17346_, _17345_, _06417_);
  or _69119_ (_17347_, _17332_, _06426_);
  and _69120_ (_17348_, _17347_, _06353_);
  and _69121_ (_17349_, _17348_, _17346_);
  or _69122_ (_17350_, _17349_, _17327_);
  and _69123_ (_17351_, _17350_, _06346_);
  or _69124_ (_17352_, _17324_, _15778_);
  and _69125_ (_17353_, _17340_, _06345_);
  and _69126_ (_17354_, _17353_, _17352_);
  or _69127_ (_17355_, _17354_, _09606_);
  or _69128_ (_17356_, _17355_, _17351_);
  nor _69129_ (_17357_, _10145_, _10132_);
  nor _69130_ (_17359_, _17357_, _10146_);
  or _69131_ (_17360_, _17359_, _09612_);
  and _69132_ (_17361_, _17360_, _06340_);
  and _69133_ (_17362_, _17361_, _17356_);
  and _69134_ (_17363_, _15745_, _08637_);
  or _69135_ (_17364_, _17363_, _17324_);
  and _69136_ (_17365_, _17364_, _06339_);
  or _69137_ (_17366_, _17365_, _10153_);
  or _69138_ (_17367_, _17366_, _17362_);
  and _69139_ (_17368_, _17367_, _17323_);
  or _69140_ (_17370_, _17368_, _09572_);
  and _69141_ (_17371_, _09172_, _08025_);
  or _69142_ (_17372_, _17314_, _06333_);
  or _69143_ (_17373_, _17372_, _17371_);
  and _69144_ (_17374_, _17373_, _06313_);
  and _69145_ (_17375_, _17374_, _17370_);
  or _69146_ (_17376_, _17375_, _17320_);
  and _69147_ (_17377_, _17376_, _10172_);
  nor _69148_ (_17378_, _17258_, _10476_);
  or _69149_ (_17379_, _17378_, _10477_);
  or _69150_ (_17381_, _17379_, _10491_);
  nand _69151_ (_17382_, _17379_, _10491_);
  and _69152_ (_17383_, _17382_, _17381_);
  or _69153_ (_17384_, _17383_, _10511_);
  or _69154_ (_17385_, _16908_, _10488_);
  and _69155_ (_17386_, _17385_, _10166_);
  and _69156_ (_17387_, _17386_, _17384_);
  or _69157_ (_17388_, _17387_, _06277_);
  or _69158_ (_17389_, _17388_, _17377_);
  and _69159_ (_17390_, _17389_, _17317_);
  or _69160_ (_17392_, _17390_, _06502_);
  and _69161_ (_17393_, _15862_, _08025_);
  or _69162_ (_17394_, _17314_, _07334_);
  or _69163_ (_17395_, _17394_, _17393_);
  and _69164_ (_17396_, _17395_, _07337_);
  and _69165_ (_17397_, _17396_, _17392_);
  and _69166_ (_17398_, _10596_, _08025_);
  or _69167_ (_17399_, _17398_, _17314_);
  and _69168_ (_17400_, _17399_, _06615_);
  or _69169_ (_17401_, _17400_, _17397_);
  and _69170_ (_17403_, _17401_, _07339_);
  or _69171_ (_17404_, _17314_, _08212_);
  and _69172_ (_17405_, _17316_, _06507_);
  and _69173_ (_17406_, _17405_, _17404_);
  or _69174_ (_17407_, _17406_, _17403_);
  and _69175_ (_17408_, _17407_, _07331_);
  and _69176_ (_17409_, _17332_, _06610_);
  and _69177_ (_17410_, _17409_, _17404_);
  or _69178_ (_17411_, _17410_, _06509_);
  or _69179_ (_17412_, _17411_, _17408_);
  and _69180_ (_17414_, _15859_, _08025_);
  or _69181_ (_17415_, _17314_, _09107_);
  or _69182_ (_17416_, _17415_, _17414_);
  and _69183_ (_17417_, _17416_, _09112_);
  and _69184_ (_17418_, _17417_, _17412_);
  nor _69185_ (_17419_, _10595_, _09574_);
  or _69186_ (_17420_, _17419_, _17314_);
  and _69187_ (_17421_, _17420_, _06602_);
  or _69188_ (_17422_, _17421_, _06639_);
  or _69189_ (_17423_, _17422_, _17418_);
  or _69190_ (_17424_, _17329_, _07048_);
  and _69191_ (_17425_, _17424_, _05990_);
  and _69192_ (_17426_, _17425_, _17423_);
  and _69193_ (_17427_, _17326_, _05989_);
  or _69194_ (_17428_, _17427_, _06646_);
  or _69195_ (_17429_, _17428_, _17426_);
  and _69196_ (_17430_, _15921_, _08025_);
  or _69197_ (_17431_, _17314_, _06651_);
  or _69198_ (_17432_, _17431_, _17430_);
  and _69199_ (_17433_, _17432_, _01442_);
  and _69200_ (_17434_, _17433_, _17429_);
  or _69201_ (_17435_, _17434_, _17313_);
  and _69202_ (_44122_, _17435_, _43634_);
  nor _69203_ (_17436_, _01442_, _06071_);
  nand _69204_ (_17437_, _10564_, _08688_);
  nor _69205_ (_17438_, _09447_, \oc8051_golden_model_1.ACC [0]);
  nor _69206_ (_17439_, _11313_, _17438_);
  or _69207_ (_17440_, _11292_, _17439_);
  nor _69208_ (_17441_, _07250_, \oc8051_golden_model_1.ACC [0]);
  nor _69209_ (_17442_, _17441_, _11271_);
  and _69210_ (_17443_, _10614_, _06360_);
  or _69211_ (_17444_, _17443_, _11246_);
  and _69212_ (_17445_, _17444_, _17442_);
  nor _69213_ (_17446_, _12641_, _10967_);
  and _69214_ (_17447_, _12641_, _10967_);
  or _69215_ (_17448_, _17447_, _17446_);
  or _69216_ (_17449_, _11218_, _17448_);
  nor _69217_ (_17450_, _17441_, _06984_);
  or _69218_ (_17451_, _17450_, _11104_);
  not _69219_ (_17452_, _10609_);
  and _69220_ (_17453_, _14566_, _08017_);
  nor _69221_ (_17454_, _08017_, _06071_);
  or _69222_ (_17455_, _17454_, _07334_);
  or _69223_ (_17456_, _17455_, _17453_);
  and _69224_ (_17457_, _06329_, _06501_);
  nand _69225_ (_17458_, _06310_, _06031_);
  and _69226_ (_17459_, _08017_, _07250_);
  or _69227_ (_17460_, _17459_, _17454_);
  or _69228_ (_17461_, _17460_, _06327_);
  not _69229_ (_17462_, _10696_);
  or _69230_ (_17463_, _17462_, _07250_);
  and _69231_ (_17464_, _10711_, _07250_);
  nor _69232_ (_17465_, _06855_, _06071_);
  and _69233_ (_17466_, _06855_, _06071_);
  or _69234_ (_17467_, _17466_, _17465_);
  and _69235_ (_17468_, _17467_, _10714_);
  or _69236_ (_17469_, _17468_, _17464_);
  and _69237_ (_17470_, _17469_, _07270_);
  or _69238_ (_17471_, _17470_, _09447_);
  or _69239_ (_17472_, _17469_, _10703_);
  and _69240_ (_17473_, _17472_, _06062_);
  or _69241_ (_17474_, _17473_, _07269_);
  and _69242_ (_17475_, _17474_, _07275_);
  and _69243_ (_17476_, _17475_, _17471_);
  nor _69244_ (_17477_, _08453_, _10619_);
  or _69245_ (_17478_, _17477_, _17454_);
  and _69246_ (_17479_, _17478_, _06474_);
  or _69247_ (_17480_, _17479_, _06356_);
  or _69248_ (_17481_, _17480_, _17476_);
  and _69249_ (_17482_, _14581_, _08645_);
  nor _69250_ (_17483_, _08645_, _06071_);
  or _69251_ (_17484_, _17483_, _06357_);
  or _69252_ (_17485_, _17484_, _17482_);
  and _69253_ (_17486_, _17485_, _06772_);
  and _69254_ (_17487_, _17486_, _17481_);
  and _69255_ (_17488_, _17460_, _06410_);
  or _69256_ (_17489_, _17488_, _10696_);
  or _69257_ (_17490_, _17489_, _17487_);
  and _69258_ (_17491_, _17490_, _17463_);
  or _69259_ (_17492_, _17491_, _07289_);
  or _69260_ (_17493_, _09447_, _07290_);
  and _69261_ (_17494_, _17493_, _06426_);
  and _69262_ (_17495_, _17494_, _17492_);
  and _69263_ (_17496_, _08453_, _06417_);
  or _69264_ (_17497_, _17496_, _10694_);
  or _69265_ (_17498_, _17497_, _17495_);
  nand _69266_ (_17499_, _10694_, _10204_);
  and _69267_ (_17500_, _17499_, _17498_);
  or _69268_ (_17501_, _17500_, _06352_);
  or _69269_ (_17502_, _17454_, _06353_);
  and _69270_ (_17503_, _17502_, _06346_);
  and _69271_ (_17504_, _17503_, _17501_);
  and _69272_ (_17505_, _17478_, _06345_);
  or _69273_ (_17506_, _17505_, _09606_);
  or _69274_ (_17507_, _17506_, _17504_);
  nand _69275_ (_17508_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand _69276_ (_17509_, _17508_, _09606_);
  and _69277_ (_17510_, _17509_, _10784_);
  and _69278_ (_17511_, _17510_, _17507_);
  nor _69279_ (_17512_, _10834_, _06071_);
  or _69280_ (_17513_, _17512_, _10835_);
  and _69281_ (_17514_, _17513_, _12338_);
  or _69282_ (_17515_, _17514_, _17511_);
  and _69283_ (_17516_, _17515_, _10854_);
  nor _69284_ (_17517_, _10902_, _06071_);
  or _69285_ (_17518_, _17517_, _10903_);
  and _69286_ (_17519_, _17518_, _10853_);
  or _69287_ (_17520_, _17519_, _06453_);
  or _69288_ (_17521_, _17520_, _17516_);
  nor _69289_ (_17522_, _10672_, _06071_);
  or _69290_ (_17523_, _17522_, _10673_);
  or _69291_ (_17524_, _17523_, _06458_);
  and _69292_ (_17525_, _17524_, _10624_);
  and _69293_ (_17526_, _17525_, _17521_);
  and _69294_ (_17527_, _17448_, _10623_);
  or _69295_ (_17528_, _17527_, _06042_);
  or _69296_ (_17529_, _17528_, _17526_);
  nand _69297_ (_17530_, _06310_, _06042_);
  and _69298_ (_17531_, _17530_, _06340_);
  and _69299_ (_17532_, _17531_, _17529_);
  and _69300_ (_17533_, _14612_, _08645_);
  or _69301_ (_17534_, _17533_, _17483_);
  and _69302_ (_17535_, _17534_, _06339_);
  or _69303_ (_17536_, _17535_, _10153_);
  or _69304_ (_17537_, _17536_, _17532_);
  and _69305_ (_17538_, _17537_, _17461_);
  or _69306_ (_17539_, _17538_, _09572_);
  and _69307_ (_17540_, _09447_, _08017_);
  or _69308_ (_17541_, _17454_, _06333_);
  or _69309_ (_17542_, _17541_, _17540_);
  and _69310_ (_17543_, _17542_, _06313_);
  and _69311_ (_17544_, _17543_, _17539_);
  and _69312_ (_17545_, _14666_, _08017_);
  or _69313_ (_17546_, _17545_, _17454_);
  and _69314_ (_17547_, _17546_, _06037_);
  or _69315_ (_17548_, _17547_, _10166_);
  or _69316_ (_17549_, _17548_, _17544_);
  nand _69317_ (_17550_, _10511_, _10166_);
  and _69318_ (_17551_, _17550_, _17549_);
  or _69319_ (_17552_, _17551_, _06031_);
  and _69320_ (_17553_, _17552_, _17458_);
  or _69321_ (_17554_, _17553_, _06277_);
  and _69322_ (_17555_, _08017_, _09008_);
  or _69323_ (_17556_, _17555_, _17454_);
  or _69324_ (_17557_, _17556_, _06278_);
  and _69325_ (_17558_, _17557_, _11029_);
  and _69326_ (_17559_, _17558_, _17554_);
  nor _69327_ (_17560_, _11029_, _06310_);
  or _69328_ (_17561_, _17560_, _17559_);
  and _69329_ (_17562_, _17561_, _11040_);
  and _69330_ (_17563_, _11048_, _11040_);
  not _69331_ (_17564_, _17563_);
  not _69332_ (_17565_, _11048_);
  or _69333_ (_17566_, _17565_, _17442_);
  and _69334_ (_17567_, _17566_, _17564_);
  or _69335_ (_17568_, _17567_, _11042_);
  or _69336_ (_17569_, _17568_, _17562_);
  not _69337_ (_17570_, _06966_);
  or _69338_ (_17571_, _17442_, _17570_);
  and _69339_ (_17572_, _06331_, _06501_);
  and _69340_ (_17573_, _06480_, _06501_);
  not _69341_ (_17574_, _17573_);
  and _69342_ (_17575_, _17574_, _11048_);
  nor _69343_ (_17576_, _17575_, _17442_);
  nor _69344_ (_17577_, _17576_, _17572_);
  and _69345_ (_17578_, _17577_, _17571_);
  and _69346_ (_17579_, _17578_, _17569_);
  and _69347_ (_17580_, _17572_, _17439_);
  nor _69348_ (_17581_, _17580_, _17579_);
  or _69349_ (_17582_, _17581_, _17457_);
  nand _69350_ (_17583_, _17439_, _17457_);
  nand _69351_ (_17584_, _17583_, _17582_);
  or _69352_ (_17585_, _17584_, _06613_);
  nand _69353_ (_17586_, _12623_, _06613_);
  and _69354_ (_17587_, _17586_, _11071_);
  and _69355_ (_17588_, _17587_, _17585_);
  and _69356_ (_17589_, _11064_, _12641_);
  or _69357_ (_17590_, _17589_, _06502_);
  or _69358_ (_17591_, _17590_, _17588_);
  and _69359_ (_17592_, _17591_, _17456_);
  or _69360_ (_17593_, _17592_, _06615_);
  or _69361_ (_17594_, _17454_, _07337_);
  and _69362_ (_17595_, _10616_, _06973_);
  and _69363_ (_17596_, _17595_, _17594_);
  and _69364_ (_17597_, _17596_, _17593_);
  not _69365_ (_17598_, _17595_);
  and _69366_ (_17599_, _17598_, _11271_);
  or _69367_ (_17600_, _17599_, _06976_);
  or _69368_ (_17601_, _17600_, _17597_);
  or _69369_ (_17602_, _11313_, _10611_);
  and _69370_ (_17603_, _17602_, _06609_);
  and _69371_ (_17604_, _17603_, _17601_);
  or _69372_ (_17605_, _11089_, _10577_);
  and _69373_ (_17606_, _17605_, _12323_);
  or _69374_ (_17607_, _17606_, _17604_);
  or _69375_ (_17608_, _11090_, _11351_);
  and _69376_ (_17609_, _17608_, _07339_);
  and _69377_ (_17610_, _17609_, _17607_);
  nand _69378_ (_17611_, _17556_, _06507_);
  nor _69379_ (_17612_, _17611_, _17477_);
  or _69380_ (_17613_, _17612_, _17610_);
  and _69381_ (_17614_, _17613_, _17452_);
  nor _69382_ (_17615_, _17441_, _17452_);
  or _69383_ (_17616_, _17615_, _11102_);
  or _69384_ (_17617_, _17616_, _17614_);
  and _69385_ (_17618_, _17617_, _17451_);
  nor _69386_ (_17619_, _17441_, _06985_);
  or _69387_ (_17620_, _17619_, _06987_);
  nor _69388_ (_17621_, _17620_, _17618_);
  and _69389_ (_17622_, _17438_, _06987_);
  or _69390_ (_17623_, _17622_, _06604_);
  or _69391_ (_17624_, _17623_, _17621_);
  not _69392_ (_17625_, _11114_);
  or _69393_ (_17626_, _12622_, _06605_);
  and _69394_ (_17627_, _17626_, _17625_);
  and _69395_ (_17628_, _17627_, _17624_);
  and _69396_ (_17629_, _11114_, _12640_);
  or _69397_ (_17630_, _17629_, _17628_);
  and _69398_ (_17631_, _17630_, _09107_);
  and _69399_ (_17632_, _14563_, _08017_);
  or _69400_ (_17633_, _17454_, _09107_);
  or _69401_ (_17634_, _17633_, _17632_);
  nand _69402_ (_17635_, _17634_, _11127_);
  nor _69403_ (_17636_, _17635_, _17631_);
  or _69404_ (_17637_, _11129_, _17513_);
  and _69405_ (_17638_, _17637_, _12839_);
  or _69406_ (_17639_, _17638_, _17636_);
  or _69407_ (_17640_, _11158_, _17518_);
  and _69408_ (_17641_, _17640_, _06601_);
  and _69409_ (_17642_, _17641_, _17639_);
  or _69410_ (_17643_, _11186_, _17523_);
  and _69411_ (_17644_, _17643_, _11188_);
  or _69412_ (_17645_, _17644_, _17642_);
  and _69413_ (_17646_, _17645_, _17449_);
  or _69414_ (_17647_, _17646_, _11216_);
  and _69415_ (_17648_, _11216_, _10967_);
  or _69416_ (_17649_, _17648_, _17443_);
  nor _69417_ (_17650_, _17649_, _11246_);
  and _69418_ (_17651_, _17650_, _17647_);
  or _69419_ (_17652_, _17651_, _17445_);
  and _69420_ (_17653_, _17652_, _07018_);
  and _69421_ (_17654_, _17442_, _07017_);
  or _69422_ (_17655_, _17654_, _11290_);
  or _69423_ (_17656_, _17655_, _17653_);
  and _69424_ (_17657_, _17656_, _17440_);
  or _69425_ (_17658_, _17657_, _06363_);
  nand _69426_ (_17659_, _12623_, _06363_);
  and _69427_ (_17660_, _17659_, _10567_);
  and _69428_ (_17661_, _17660_, _17658_);
  and _69429_ (_17662_, _12641_, _10566_);
  or _69430_ (_17663_, _17662_, _10564_);
  or _69431_ (_17664_, _17663_, _17661_);
  and _69432_ (_17665_, _17664_, _17437_);
  or _69433_ (_17666_, _17665_, _06639_);
  or _69434_ (_17667_, _17478_, _07048_);
  and _69435_ (_17668_, _17667_, _11378_);
  and _69436_ (_17669_, _17668_, _17666_);
  nor _69437_ (_17670_, _11382_, _06071_);
  nor _69438_ (_17671_, _17670_, _13072_);
  or _69439_ (_17672_, _17671_, _17669_);
  nand _69440_ (_17673_, _11382_, _06097_);
  and _69441_ (_17674_, _17673_, _05990_);
  and _69442_ (_17675_, _17674_, _17672_);
  and _69443_ (_17676_, _17454_, _05989_);
  or _69444_ (_17677_, _17676_, _06646_);
  or _69445_ (_17678_, _17677_, _17675_);
  or _69446_ (_17679_, _17478_, _06651_);
  and _69447_ (_17680_, _17679_, _11401_);
  and _69448_ (_17681_, _17680_, _17678_);
  nor _69449_ (_17682_, _11407_, _06071_);
  nor _69450_ (_17683_, _17682_, _13095_);
  or _69451_ (_17684_, _17683_, _17681_);
  nand _69452_ (_17685_, _11407_, _06097_);
  and _69453_ (_17686_, _17685_, _01442_);
  and _69454_ (_17687_, _17686_, _17684_);
  or _69455_ (_17688_, _17687_, _17436_);
  and _69456_ (_44123_, _17688_, _43634_);
  nor _69457_ (_17689_, _01442_, _06097_);
  and _69458_ (_17690_, _06331_, _06360_);
  not _69459_ (_17691_, _17690_);
  nor _69460_ (_17692_, _11313_, _11312_);
  nor _69461_ (_17693_, _17692_, _11314_);
  or _69462_ (_17694_, _17693_, _17691_);
  nand _69463_ (_17695_, _11269_, _10609_);
  and _69464_ (_17696_, _06785_, _06506_);
  nor _69465_ (_17697_, _08017_, _06097_);
  or _69466_ (_17698_, _17697_, _07337_);
  nor _69467_ (_17699_, _10619_, _07448_);
  or _69468_ (_17700_, _17699_, _17697_);
  or _69469_ (_17701_, _17700_, _06327_);
  not _69470_ (_17702_, _11312_);
  nor _69471_ (_17703_, _10896_, _06071_);
  or _69472_ (_17704_, _17703_, _10901_);
  nand _69473_ (_17705_, _17704_, _17702_);
  or _69474_ (_17706_, _17704_, _17702_);
  and _69475_ (_17707_, _17706_, _10853_);
  and _69476_ (_17708_, _17707_, _17705_);
  nand _69477_ (_17709_, _10696_, _07448_);
  nor _69478_ (_17710_, _10712_, _07448_);
  nor _69479_ (_17711_, _06855_, _06097_);
  and _69480_ (_17712_, _06855_, _06097_);
  or _69481_ (_17713_, _17712_, _17711_);
  and _69482_ (_17714_, _17713_, _10714_);
  or _69483_ (_17715_, _17714_, _17710_);
  or _69484_ (_17716_, _17715_, _10703_);
  and _69485_ (_17717_, _17716_, _06062_);
  or _69486_ (_17718_, _17717_, _07269_);
  and _69487_ (_17719_, _17715_, _07270_);
  or _69488_ (_17720_, _17719_, _09402_);
  and _69489_ (_17721_, _17720_, _17718_);
  or _69490_ (_17722_, _17721_, _06474_);
  or _69491_ (_17723_, _08017_, \oc8051_golden_model_1.ACC [1]);
  and _69492_ (_17724_, _14744_, _08017_);
  not _69493_ (_17725_, _17724_);
  and _69494_ (_17726_, _17725_, _17723_);
  or _69495_ (_17727_, _17726_, _07275_);
  and _69496_ (_17728_, _17727_, _17722_);
  or _69497_ (_17729_, _17728_, _10729_);
  nor _69498_ (_17730_, _10733_, \oc8051_golden_model_1.PSW [6]);
  nor _69499_ (_17731_, _17730_, \oc8051_golden_model_1.ACC [1]);
  and _69500_ (_17732_, _17730_, \oc8051_golden_model_1.ACC [1]);
  nor _69501_ (_17733_, _17732_, _17731_);
  nand _69502_ (_17734_, _17733_, _10729_);
  and _69503_ (_17735_, _17734_, _06418_);
  and _69504_ (_17736_, _17735_, _17729_);
  nor _69505_ (_17737_, _08645_, _06097_);
  and _69506_ (_17738_, _14767_, _08645_);
  or _69507_ (_17739_, _17738_, _17737_);
  and _69508_ (_17740_, _17739_, _06356_);
  and _69509_ (_17741_, _17700_, _06410_);
  or _69510_ (_17742_, _17741_, _10696_);
  or _69511_ (_17743_, _17742_, _17740_);
  or _69512_ (_17744_, _17743_, _17736_);
  and _69513_ (_17745_, _17744_, _17709_);
  or _69514_ (_17746_, _17745_, _07289_);
  or _69515_ (_17747_, _09402_, _07290_);
  and _69516_ (_17748_, _17747_, _06426_);
  and _69517_ (_17749_, _17748_, _17746_);
  nor _69518_ (_17750_, _08403_, _06426_);
  or _69519_ (_17751_, _17750_, _10694_);
  or _69520_ (_17752_, _17751_, _17749_);
  nand _69521_ (_17753_, _10694_, _10237_);
  and _69522_ (_17754_, _17753_, _17752_);
  or _69523_ (_17755_, _17754_, _06352_);
  and _69524_ (_17756_, _14754_, _08645_);
  or _69525_ (_17757_, _17756_, _17737_);
  or _69526_ (_17758_, _17757_, _06353_);
  and _69527_ (_17759_, _17758_, _06346_);
  and _69528_ (_17760_, _17759_, _17755_);
  or _69529_ (_17761_, _17737_, _14782_);
  and _69530_ (_17762_, _17739_, _06345_);
  and _69531_ (_17763_, _17762_, _17761_);
  or _69532_ (_17764_, _17763_, _17760_);
  and _69533_ (_17765_, _17764_, _09612_);
  nor _69534_ (_17766_, _10094_, _10093_);
  nor _69535_ (_17767_, _17766_, _10095_);
  and _69536_ (_17768_, _17767_, _09606_);
  or _69537_ (_17769_, _17768_, _12338_);
  or _69538_ (_17770_, _17769_, _17765_);
  nor _69539_ (_17771_, _10787_, _06071_);
  or _69540_ (_17772_, _17771_, _10833_);
  nor _69541_ (_17773_, _17772_, _11270_);
  and _69542_ (_17774_, _17772_, _11270_);
  or _69543_ (_17775_, _17774_, _17773_);
  or _69544_ (_17776_, _17775_, _10784_);
  and _69545_ (_17777_, _17776_, _10854_);
  and _69546_ (_17778_, _17777_, _17770_);
  or _69547_ (_17779_, _17778_, _17708_);
  and _69548_ (_17780_, _17779_, _06458_);
  nor _69549_ (_17781_, _10666_, _06071_);
  or _69550_ (_17782_, _17781_, _10671_);
  or _69551_ (_17783_, _17782_, _12621_);
  nand _69552_ (_17784_, _17782_, _12621_);
  and _69553_ (_17785_, _17784_, _06453_);
  and _69554_ (_17786_, _17785_, _17783_);
  or _69555_ (_17787_, _17786_, _17780_);
  and _69556_ (_17788_, _17787_, _10624_);
  nor _69557_ (_17789_, _06310_, \oc8051_golden_model_1.ACC [0]);
  not _69558_ (_17790_, _17789_);
  and _69559_ (_17791_, _11354_, _17790_);
  nor _69560_ (_17792_, _11354_, _17790_);
  or _69561_ (_17793_, _17792_, _17791_);
  nor _69562_ (_17794_, _17446_, _17793_);
  and _69563_ (_17795_, _12642_, \oc8051_golden_model_1.PSW [7]);
  or _69564_ (_17796_, _17795_, _17794_);
  and _69565_ (_17797_, _17796_, _10623_);
  or _69566_ (_17798_, _17797_, _06042_);
  or _69567_ (_17799_, _17798_, _17788_);
  nand _69568_ (_17800_, _07127_, _06042_);
  and _69569_ (_17801_, _17800_, _06340_);
  and _69570_ (_17802_, _17801_, _17799_);
  and _69571_ (_17803_, _14796_, _08645_);
  or _69572_ (_17804_, _17803_, _17737_);
  and _69573_ (_17805_, _17804_, _06339_);
  or _69574_ (_17806_, _17805_, _10153_);
  or _69575_ (_17807_, _17806_, _17802_);
  and _69576_ (_17808_, _17807_, _17701_);
  or _69577_ (_17809_, _17808_, _09572_);
  and _69578_ (_17810_, _09402_, _08017_);
  or _69579_ (_17811_, _17697_, _06333_);
  or _69580_ (_17812_, _17811_, _17810_);
  and _69581_ (_17813_, _17812_, _06313_);
  and _69582_ (_17814_, _17813_, _17809_);
  or _69583_ (_17815_, _14851_, _10619_);
  and _69584_ (_17816_, _17723_, _06037_);
  and _69585_ (_17817_, _17816_, _17815_);
  or _69586_ (_17818_, _17817_, _10166_);
  or _69587_ (_17819_, _17818_, _17814_);
  nand _69588_ (_17820_, _10421_, _10166_);
  and _69589_ (_17821_, _17820_, _17819_);
  or _69590_ (_17822_, _17821_, _06031_);
  nand _69591_ (_17823_, _07127_, _06031_);
  and _69592_ (_17824_, _17823_, _06278_);
  and _69593_ (_17825_, _17824_, _17822_);
  nand _69594_ (_17826_, _08017_, _07160_);
  and _69595_ (_17827_, _17826_, _06277_);
  and _69596_ (_17828_, _17827_, _17723_);
  or _69597_ (_17829_, _17828_, _11028_);
  or _69598_ (_17830_, _17829_, _17825_);
  nand _69599_ (_17831_, _11028_, _07127_);
  and _69600_ (_17832_, _17563_, _11043_);
  and _69601_ (_17833_, _17832_, _17831_);
  and _69602_ (_17834_, _17833_, _17830_);
  not _69603_ (_17835_, _17832_);
  and _69604_ (_17836_, _17835_, _11270_);
  or _69605_ (_17837_, _17836_, _11052_);
  or _69606_ (_17838_, _17837_, _17834_);
  or _69607_ (_17839_, _11060_, _11312_);
  and _69608_ (_17840_, _17839_, _17838_);
  or _69609_ (_17841_, _17840_, _06613_);
  or _69610_ (_17842_, _10579_, _06614_);
  and _69611_ (_17843_, _17842_, _11071_);
  and _69612_ (_17844_, _17843_, _17841_);
  nor _69613_ (_17845_, _11071_, _11354_);
  or _69614_ (_17846_, _17845_, _17844_);
  and _69615_ (_17847_, _17846_, _07334_);
  or _69616_ (_17848_, _14749_, _10619_);
  and _69617_ (_17849_, _17723_, _06502_);
  and _69618_ (_17850_, _17849_, _17848_);
  or _69619_ (_17851_, _17850_, _06615_);
  or _69620_ (_17852_, _17851_, _17847_);
  and _69621_ (_17853_, _17852_, _17698_);
  or _69622_ (_17854_, _17853_, _17696_);
  nand _69623_ (_17855_, _06323_, _06506_);
  nor _69624_ (_17856_, _06319_, _06017_);
  not _69625_ (_17857_, _17856_);
  not _69626_ (_17858_, _06828_);
  and _69627_ (_17859_, _11268_, _17858_);
  or _69628_ (_17860_, _17859_, _17857_);
  and _69629_ (_17861_, _17860_, _17855_);
  and _69630_ (_17862_, _17861_, _17854_);
  and _69631_ (_17863_, _06315_, _06506_);
  not _69632_ (_17864_, _17855_);
  or _69633_ (_17865_, _17864_, _06828_);
  and _69634_ (_17866_, _17865_, _11268_);
  or _69635_ (_17867_, _17866_, _17863_);
  or _69636_ (_17868_, _17867_, _17862_);
  not _69637_ (_17869_, _17863_);
  or _69638_ (_17870_, _17869_, _11268_);
  and _69639_ (_17871_, _17870_, _10611_);
  and _69640_ (_17872_, _17871_, _17868_);
  and _69641_ (_17873_, _11309_, _06976_);
  or _69642_ (_17874_, _17873_, _06608_);
  or _69643_ (_17875_, _17874_, _17872_);
  or _69644_ (_17876_, _10576_, _06609_);
  and _69645_ (_17877_, _17876_, _11090_);
  and _69646_ (_17878_, _17877_, _17875_);
  and _69647_ (_17879_, _11089_, _11350_);
  or _69648_ (_17880_, _17879_, _17878_);
  and _69649_ (_17881_, _17880_, _07339_);
  or _69650_ (_17882_, _14747_, _10619_);
  and _69651_ (_17883_, _17723_, _06507_);
  and _69652_ (_17884_, _17883_, _17882_);
  or _69653_ (_17885_, _17884_, _10609_);
  or _69654_ (_17886_, _17885_, _17881_);
  and _69655_ (_17887_, _17886_, _17695_);
  or _69656_ (_17888_, _17887_, _11102_);
  nor _69657_ (_17889_, _11269_, _06984_);
  or _69658_ (_17890_, _17889_, _11104_);
  and _69659_ (_17891_, _17890_, _17888_);
  nor _69660_ (_17892_, _11269_, _06985_);
  or _69661_ (_17893_, _17892_, _06987_);
  or _69662_ (_17894_, _17893_, _17891_);
  nand _69663_ (_17895_, _11311_, _06987_);
  and _69664_ (_17896_, _17895_, _06605_);
  and _69665_ (_17897_, _17896_, _17894_);
  nor _69666_ (_17898_, _10578_, _06605_);
  or _69667_ (_17899_, _17898_, _11114_);
  or _69668_ (_17900_, _17899_, _17897_);
  and _69669_ (_17901_, _11114_, _06097_);
  nand _69670_ (_17902_, _17901_, _07127_);
  and _69671_ (_17903_, _17902_, _09107_);
  and _69672_ (_17904_, _17903_, _17900_);
  or _69673_ (_17905_, _17826_, _08404_);
  and _69674_ (_17906_, _17723_, _06509_);
  and _69675_ (_17907_, _17906_, _17905_);
  or _69676_ (_17908_, _17907_, _11122_);
  or _69677_ (_17909_, _17908_, _17904_);
  nor _69678_ (_17910_, _11139_, _11138_);
  nor _69679_ (_17911_, _17910_, _11140_);
  or _69680_ (_17912_, _17911_, _11123_);
  and _69681_ (_17913_, _17912_, _11126_);
  and _69682_ (_17914_, _17913_, _17909_);
  not _69683_ (_17915_, _11126_);
  and _69684_ (_17916_, _17911_, _17915_);
  or _69685_ (_17917_, _17916_, _17914_);
  and _69686_ (_17918_, _17917_, _11158_);
  nor _69687_ (_17919_, _11167_, _11166_);
  nor _69688_ (_17920_, _17919_, _11168_);
  and _69689_ (_17921_, _17920_, _07002_);
  and _69690_ (_17922_, _06331_, _06511_);
  and _69691_ (_17923_, _17920_, _17922_);
  or _69692_ (_17924_, _17923_, _06600_);
  or _69693_ (_17925_, _17924_, _17921_);
  or _69694_ (_17926_, _17925_, _17918_);
  nor _69695_ (_17927_, _11197_, _11196_);
  nor _69696_ (_17928_, _17927_, _11198_);
  or _69697_ (_17929_, _17928_, _06601_);
  and _69698_ (_17930_, _17929_, _11218_);
  and _69699_ (_17931_, _17930_, _17926_);
  or _69700_ (_17932_, _11226_, _10974_);
  nor _69701_ (_17933_, _11227_, _11218_);
  and _69702_ (_17934_, _17933_, _17932_);
  or _69703_ (_17935_, _17934_, _11216_);
  or _69704_ (_17936_, _17935_, _17931_);
  nand _69705_ (_17937_, _11216_, _06071_);
  and _69706_ (_17938_, _17937_, _11248_);
  and _69707_ (_17939_, _17938_, _17936_);
  or _69708_ (_17940_, _11271_, _11270_);
  nor _69709_ (_17941_, _11272_, _11248_);
  and _69710_ (_17942_, _17941_, _17940_);
  or _69711_ (_17943_, _17942_, _17690_);
  or _69712_ (_17944_, _17943_, _17939_);
  and _69713_ (_17945_, _17944_, _17694_);
  or _69714_ (_17946_, _17945_, _07019_);
  or _69715_ (_17947_, _17693_, _07020_);
  and _69716_ (_17948_, _17947_, _06364_);
  and _69717_ (_17949_, _17948_, _17946_);
  nor _69718_ (_17950_, _10579_, _10577_);
  nor _69719_ (_17951_, _17950_, _10580_);
  and _69720_ (_17952_, _17951_, _06363_);
  or _69721_ (_17953_, _17952_, _10566_);
  or _69722_ (_17954_, _17953_, _17949_);
  nor _69723_ (_17955_, _11355_, _11351_);
  nor _69724_ (_17956_, _17955_, _11356_);
  or _69725_ (_17957_, _17956_, _10567_);
  and _69726_ (_17958_, _17957_, _13049_);
  and _69727_ (_17959_, _17958_, _17954_);
  and _69728_ (_17960_, _10564_, \oc8051_golden_model_1.ACC [0]);
  or _69729_ (_17961_, _17960_, _06639_);
  or _69730_ (_17962_, _17961_, _17959_);
  or _69731_ (_17963_, _17726_, _07048_);
  and _69732_ (_17964_, _17963_, _11378_);
  and _69733_ (_17965_, _17964_, _17962_);
  nor _69734_ (_17966_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor _69735_ (_17967_, _11408_, _17966_);
  nor _69736_ (_17968_, _17967_, _11378_);
  or _69737_ (_17969_, _17968_, _17965_);
  or _69738_ (_17970_, _17969_, _11382_);
  nand _69739_ (_17971_, _11382_, _10280_);
  and _69740_ (_17972_, _17971_, _05990_);
  and _69741_ (_17973_, _17972_, _17970_);
  and _69742_ (_17974_, _17757_, _05989_);
  or _69743_ (_17975_, _17974_, _06646_);
  or _69744_ (_17976_, _17975_, _17973_);
  or _69745_ (_17977_, _17697_, _06651_);
  or _69746_ (_17978_, _17977_, _17724_);
  and _69747_ (_17979_, _17978_, _11401_);
  and _69748_ (_17980_, _17979_, _17976_);
  and _69749_ (_17981_, _17967_, _11400_);
  or _69750_ (_17983_, _17981_, _11407_);
  or _69751_ (_17984_, _17983_, _17980_);
  nand _69752_ (_17985_, _11407_, _10280_);
  and _69753_ (_17986_, _17985_, _01442_);
  and _69754_ (_17987_, _17986_, _17984_);
  or _69755_ (_17988_, _17987_, _17689_);
  and _69756_ (_44125_, _17988_, _43634_);
  nor _69757_ (_17989_, _01442_, _10280_);
  nand _69758_ (_17990_, _10564_, _06097_);
  and _69759_ (_17991_, _10584_, _10581_);
  nor _69760_ (_17992_, _17991_, _10585_);
  or _69761_ (_17993_, _17992_, _06364_);
  and _69762_ (_17994_, _17993_, _10567_);
  nand _69763_ (_17995_, _11114_, _11348_);
  or _69764_ (_17996_, _11306_, _10611_);
  or _69765_ (_17997_, _10583_, _06614_);
  and _69766_ (_17998_, _17997_, _11071_);
  nand _69767_ (_17999_, _06727_, _06031_);
  nor _69768_ (_18000_, _08017_, _10280_);
  nor _69769_ (_18001_, _10619_, _07854_);
  or _69770_ (_18002_, _18001_, _18000_);
  or _69771_ (_18003_, _18002_, _06327_);
  nand _69772_ (_18004_, _10696_, _07854_);
  nor _69773_ (_18005_, _10712_, _07854_);
  nor _69774_ (_18006_, _06855_, _10280_);
  and _69775_ (_18007_, _06855_, _10280_);
  or _69776_ (_18008_, _18007_, _18006_);
  and _69777_ (_18009_, _18008_, _10714_);
  or _69778_ (_18010_, _18009_, _18005_);
  or _69779_ (_18011_, _18010_, _10703_);
  and _69780_ (_18012_, _18011_, _06062_);
  or _69781_ (_18013_, _18012_, _07269_);
  and _69782_ (_18014_, _18010_, _07270_);
  or _69783_ (_18015_, _18014_, _09356_);
  and _69784_ (_18016_, _18015_, _18013_);
  and _69785_ (_18017_, _18016_, _07275_);
  and _69786_ (_18018_, _14959_, _08017_);
  or _69787_ (_18019_, _18018_, _18000_);
  and _69788_ (_18020_, _18019_, _06474_);
  or _69789_ (_18021_, _18020_, _10729_);
  or _69790_ (_18022_, _18021_, _18017_);
  nor _69791_ (_18023_, _17731_, _10280_);
  and _69792_ (_18024_, _10732_, \oc8051_golden_model_1.PSW [6]);
  nor _69793_ (_18025_, _18024_, _18023_);
  nand _69794_ (_18026_, _18025_, _10729_);
  and _69795_ (_18027_, _18026_, _06418_);
  and _69796_ (_18028_, _18027_, _18022_);
  nor _69797_ (_18029_, _08645_, _10280_);
  and _69798_ (_18030_, _14955_, _08645_);
  or _69799_ (_18031_, _18030_, _18029_);
  and _69800_ (_18032_, _18031_, _06356_);
  and _69801_ (_18033_, _18002_, _06410_);
  or _69802_ (_18034_, _18033_, _10696_);
  or _69803_ (_18035_, _18034_, _18032_);
  or _69804_ (_18036_, _18035_, _18028_);
  and _69805_ (_18037_, _18036_, _18004_);
  or _69806_ (_18038_, _18037_, _07289_);
  or _69807_ (_18039_, _09356_, _07290_);
  and _69808_ (_18040_, _18039_, _06426_);
  and _69809_ (_18041_, _18040_, _18038_);
  nor _69810_ (_18042_, _08502_, _06426_);
  or _69811_ (_18043_, _18042_, _10694_);
  or _69812_ (_18044_, _18043_, _18041_);
  nand _69813_ (_18045_, _10694_, _10193_);
  and _69814_ (_18046_, _18045_, _18044_);
  or _69815_ (_18047_, _18046_, _06352_);
  and _69816_ (_18048_, _14953_, _08645_);
  or _69817_ (_18049_, _18048_, _18029_);
  or _69818_ (_18050_, _18049_, _06353_);
  and _69819_ (_18051_, _18050_, _06346_);
  and _69820_ (_18052_, _18051_, _18047_);
  or _69821_ (_18053_, _18029_, _14986_);
  and _69822_ (_18054_, _18031_, _06345_);
  and _69823_ (_18055_, _18054_, _18053_);
  or _69824_ (_18056_, _18055_, _09606_);
  or _69825_ (_18057_, _18056_, _18052_);
  nor _69826_ (_18058_, _10097_, _10095_);
  or _69827_ (_18059_, _18058_, _10098_);
  nand _69828_ (_18060_, _18059_, _09606_);
  and _69829_ (_18061_, _18060_, _10784_);
  and _69830_ (_18062_, _18061_, _18057_);
  and _69831_ (_18063_, _06331_, _06038_);
  and _69832_ (_18064_, _07448_, \oc8051_golden_model_1.ACC [1]);
  and _69833_ (_18065_, _07250_, _06071_);
  nor _69834_ (_18066_, _18065_, _11270_);
  nor _69835_ (_18067_, _18066_, _18064_);
  nor _69836_ (_18068_, _11266_, _18067_);
  and _69837_ (_18069_, _11266_, _18067_);
  nor _69838_ (_18070_, _18069_, _18068_);
  nor _69839_ (_18071_, _17442_, _11270_);
  and _69840_ (_18072_, _18071_, \oc8051_golden_model_1.PSW [7]);
  or _69841_ (_18073_, _18072_, _18070_);
  nand _69842_ (_18074_, _18072_, _18070_);
  and _69843_ (_18075_, _18074_, _12338_);
  and _69844_ (_18076_, _18075_, _18073_);
  or _69845_ (_18077_, _18076_, _18063_);
  or _69846_ (_18078_, _18077_, _18062_);
  and _69847_ (_18079_, _11310_, \oc8051_golden_model_1.ACC [1]);
  and _69848_ (_18080_, _09447_, _06071_);
  nor _69849_ (_18081_, _18080_, _11312_);
  nor _69850_ (_18082_, _18081_, _18079_);
  nor _69851_ (_18083_, _11308_, _18082_);
  and _69852_ (_18084_, _11308_, _18082_);
  nor _69853_ (_18085_, _18084_, _18083_);
  nor _69854_ (_18086_, _17439_, _11312_);
  not _69855_ (_18087_, _18086_);
  or _69856_ (_18088_, _18087_, _18085_);
  and _69857_ (_18089_, _18088_, \oc8051_golden_model_1.PSW [7]);
  nor _69858_ (_18090_, _18085_, \oc8051_golden_model_1.PSW [7]);
  nor _69859_ (_18091_, _18090_, _18089_);
  and _69860_ (_18092_, _18087_, _18085_);
  or _69861_ (_18093_, _18092_, _18091_);
  and _69862_ (_18094_, _18093_, _06028_);
  or _69863_ (_18095_, _18094_, _10854_);
  and _69864_ (_18096_, _18095_, _18078_);
  and _69865_ (_18097_, _18093_, _06909_);
  or _69866_ (_18098_, _18097_, _06453_);
  or _69867_ (_18099_, _18098_, _18096_);
  and _69868_ (_18100_, _08403_, \oc8051_golden_model_1.ACC [1]);
  and _69869_ (_18101_, _08453_, _06071_);
  nor _69870_ (_18102_, _18101_, _14324_);
  nor _69871_ (_18103_, _18102_, _18100_);
  nor _69872_ (_18104_, _18103_, _10583_);
  and _69873_ (_18105_, _18103_, _10583_);
  nor _69874_ (_18106_, _18105_, _18104_);
  and _69875_ (_18107_, _12624_, \oc8051_golden_model_1.PSW [7]);
  nand _69876_ (_18108_, _18107_, _18106_);
  or _69877_ (_18109_, _18107_, _18106_);
  and _69878_ (_18110_, _18109_, _18108_);
  or _69879_ (_18111_, _18110_, _06458_);
  and _69880_ (_18112_, _18111_, _10624_);
  and _69881_ (_18113_, _18112_, _18099_);
  nor _69882_ (_18114_, _17791_, _11352_);
  nor _69883_ (_18115_, _11349_, _18114_);
  and _69884_ (_18116_, _11349_, _18114_);
  nor _69885_ (_18117_, _18116_, _18115_);
  not _69886_ (_18118_, _17795_);
  or _69887_ (_18119_, _18118_, _18117_);
  nand _69888_ (_18120_, _18118_, _18117_);
  nand _69889_ (_18121_, _18120_, _18119_);
  and _69890_ (_18122_, _18121_, _10623_);
  or _69891_ (_18123_, _18122_, _06042_);
  or _69892_ (_18124_, _18123_, _18113_);
  nand _69893_ (_18125_, _06727_, _06042_);
  and _69894_ (_18126_, _18125_, _06340_);
  and _69895_ (_18127_, _18126_, _18124_);
  and _69896_ (_18128_, _15000_, _08645_);
  or _69897_ (_18129_, _18128_, _18029_);
  and _69898_ (_18130_, _18129_, _06339_);
  or _69899_ (_18131_, _18130_, _10153_);
  or _69900_ (_18132_, _18131_, _18127_);
  and _69901_ (_18133_, _18132_, _18003_);
  or _69902_ (_18134_, _18133_, _09572_);
  and _69903_ (_18135_, _09356_, _08017_);
  or _69904_ (_18136_, _18000_, _06333_);
  or _69905_ (_18137_, _18136_, _18135_);
  and _69906_ (_18138_, _18137_, _06313_);
  and _69907_ (_18139_, _18138_, _18134_);
  and _69908_ (_18140_, _15056_, _08017_);
  or _69909_ (_18141_, _18140_, _18000_);
  and _69910_ (_18142_, _18141_, _06037_);
  or _69911_ (_18143_, _18142_, _10166_);
  or _69912_ (_18144_, _18143_, _18139_);
  or _69913_ (_18145_, _10358_, _10172_);
  and _69914_ (_18146_, _18145_, _18144_);
  or _69915_ (_18147_, _18146_, _06031_);
  and _69916_ (_18148_, _18147_, _17999_);
  or _69917_ (_18149_, _18148_, _06277_);
  and _69918_ (_18150_, _08017_, _09057_);
  or _69919_ (_18151_, _18150_, _18000_);
  or _69920_ (_18152_, _18151_, _06278_);
  and _69921_ (_18153_, _18152_, _11029_);
  nand _69922_ (_18154_, _18153_, _18149_);
  or _69923_ (_18155_, _11029_, _06727_);
  and _69924_ (_18156_, _18155_, _11040_);
  nand _69925_ (_18157_, _18156_, _18154_);
  nor _69926_ (_18158_, _11040_, _11266_);
  nor _69927_ (_18159_, _18158_, _17565_);
  and _69928_ (_18160_, _18159_, _18157_);
  nor _69929_ (_18161_, _17573_, _11266_);
  nor _69930_ (_18162_, _18161_, _17575_);
  or _69931_ (_18163_, _18162_, _06966_);
  or _69932_ (_18164_, _18163_, _18160_);
  or _69933_ (_18165_, _11266_, _11043_);
  and _69934_ (_18166_, _18165_, _11060_);
  and _69935_ (_18167_, _18166_, _18164_);
  and _69936_ (_18168_, _11052_, _11308_);
  or _69937_ (_18169_, _18168_, _06613_);
  or _69938_ (_18170_, _18169_, _18167_);
  and _69939_ (_18171_, _18170_, _17998_);
  and _69940_ (_18172_, _11064_, _11349_);
  or _69941_ (_18173_, _18172_, _06502_);
  or _69942_ (_18174_, _18173_, _18171_);
  and _69943_ (_18175_, _14948_, _08017_);
  or _69944_ (_18176_, _18175_, _18000_);
  or _69945_ (_18177_, _18176_, _07334_);
  and _69946_ (_18178_, _18177_, _18174_);
  or _69947_ (_18179_, _18178_, _06615_);
  or _69948_ (_18180_, _18000_, _07337_);
  and _69949_ (_18181_, _18180_, _17857_);
  and _69950_ (_18182_, _18181_, _18179_);
  and _69951_ (_18183_, _11264_, _17856_);
  or _69952_ (_18184_, _18183_, _17864_);
  or _69953_ (_18185_, _18184_, _18182_);
  or _69954_ (_18186_, _11264_, _17855_);
  and _69955_ (_18187_, _18186_, _17869_);
  and _69956_ (_18188_, _18187_, _18185_);
  and _69957_ (_18189_, _17863_, _11264_);
  or _69958_ (_18190_, _18189_, _06976_);
  or _69959_ (_18191_, _18190_, _18188_);
  and _69960_ (_18192_, _18191_, _17996_);
  or _69961_ (_18193_, _18192_, _06608_);
  or _69962_ (_18194_, _10575_, _06609_);
  and _69963_ (_18195_, _18194_, _11090_);
  and _69964_ (_18196_, _18195_, _18193_);
  and _69965_ (_18197_, _11089_, _11347_);
  or _69966_ (_18198_, _18197_, _18196_);
  and _69967_ (_18199_, _18198_, _07339_);
  and _69968_ (_18200_, _07577_, _06508_);
  nand _69969_ (_18201_, _18151_, _06507_);
  nor _69970_ (_18202_, _18201_, _10582_);
  or _69971_ (_18203_, _18202_, _18200_);
  or _69972_ (_18204_, _18203_, _18199_);
  nand _69973_ (_18205_, _18200_, _11265_);
  and _69974_ (_18206_, _06315_, _06508_);
  not _69975_ (_18207_, _18206_);
  and _69976_ (_18208_, _18207_, _18205_);
  and _69977_ (_18209_, _18208_, _18204_);
  nor _69978_ (_18210_, _18207_, _11265_);
  or _69979_ (_18211_, _18210_, _06987_);
  or _69980_ (_18212_, _18211_, _18209_);
  nand _69981_ (_18213_, _11307_, _06987_);
  and _69982_ (_18214_, _18213_, _06605_);
  and _69983_ (_18215_, _18214_, _18212_);
  nand _69984_ (_18216_, _17625_, _10582_);
  and _69985_ (_18217_, _18216_, _12315_);
  or _69986_ (_18218_, _18217_, _18215_);
  and _69987_ (_18219_, _18218_, _17995_);
  or _69988_ (_18220_, _18219_, _06509_);
  and _69989_ (_18221_, _14945_, _08017_);
  or _69990_ (_18222_, _18000_, _09107_);
  or _69991_ (_18223_, _18222_, _18221_);
  and _69992_ (_18224_, _18223_, _11127_);
  and _69993_ (_18225_, _18224_, _18220_);
  nand _69994_ (_18226_, _11141_, _10827_);
  nor _69995_ (_18227_, _11142_, _11127_);
  and _69996_ (_18228_, _18227_, _18226_);
  or _69997_ (_18229_, _18228_, _17922_);
  or _69998_ (_18230_, _18229_, _18225_);
  not _69999_ (_18231_, _17922_);
  and _70000_ (_18232_, _11169_, _10894_);
  nor _70001_ (_18233_, _18232_, _11170_);
  or _70002_ (_18234_, _18233_, _18231_);
  and _70003_ (_18235_, _18234_, _18230_);
  or _70004_ (_18236_, _18235_, _07002_);
  not _70005_ (_18237_, _07002_);
  or _70006_ (_18238_, _18233_, _18237_);
  and _70007_ (_18239_, _18238_, _06601_);
  and _70008_ (_18240_, _18239_, _18236_);
  nand _70009_ (_18241_, _11199_, _10664_);
  nor _70010_ (_18242_, _11200_, _06601_);
  and _70011_ (_18243_, _18242_, _18241_);
  or _70012_ (_18244_, _18243_, _18240_);
  and _70013_ (_18245_, _18244_, _11218_);
  nand _70014_ (_18246_, _11228_, _10965_);
  nor _70015_ (_18247_, _11229_, _11218_);
  and _70016_ (_18248_, _18247_, _18246_);
  or _70017_ (_18249_, _18248_, _11216_);
  or _70018_ (_18250_, _18249_, _18245_);
  nand _70019_ (_18251_, _11216_, _06097_);
  and _70020_ (_18252_, _18251_, _11248_);
  and _70021_ (_18253_, _18252_, _18250_);
  not _70022_ (_18254_, _11248_);
  and _70023_ (_18255_, _11273_, _11267_);
  nor _70024_ (_18256_, _18255_, _11274_);
  and _70025_ (_18257_, _18256_, _18254_);
  or _70026_ (_18258_, _18257_, _17690_);
  or _70027_ (_18259_, _18258_, _18253_);
  nor _70028_ (_18260_, _11316_, _11308_);
  nor _70029_ (_18261_, _18260_, _11317_);
  and _70030_ (_18262_, _18261_, _07020_);
  or _70031_ (_18263_, _18262_, _11292_);
  and _70032_ (_18264_, _18263_, _18259_);
  and _70033_ (_18265_, _18261_, _07019_);
  or _70034_ (_18266_, _18265_, _06363_);
  or _70035_ (_18267_, _18266_, _18264_);
  and _70036_ (_18268_, _18267_, _17994_);
  or _70037_ (_18269_, _11358_, _11349_);
  nor _70038_ (_18270_, _11359_, _10567_);
  and _70039_ (_18271_, _18270_, _18269_);
  or _70040_ (_18272_, _18271_, _10564_);
  or _70041_ (_18273_, _18272_, _18268_);
  and _70042_ (_18274_, _18273_, _17990_);
  or _70043_ (_18275_, _18274_, _06639_);
  or _70044_ (_18276_, _18019_, _07048_);
  and _70045_ (_18277_, _18276_, _11378_);
  and _70046_ (_18278_, _18277_, _18275_);
  nor _70047_ (_18279_, _17966_, _10280_);
  or _70048_ (_18280_, _18279_, _11383_);
  and _70049_ (_18281_, _18280_, _11377_);
  or _70050_ (_18282_, _18281_, _11382_);
  or _70051_ (_18283_, _18282_, _18278_);
  nand _70052_ (_18284_, _11382_, _10334_);
  and _70053_ (_18285_, _18284_, _05990_);
  and _70054_ (_18286_, _18285_, _18283_);
  and _70055_ (_18287_, _18049_, _05989_);
  or _70056_ (_18288_, _18287_, _06646_);
  or _70057_ (_18289_, _18288_, _18286_);
  and _70058_ (_18290_, _15129_, _08017_);
  or _70059_ (_18291_, _18000_, _06651_);
  or _70060_ (_18292_, _18291_, _18290_);
  and _70061_ (_18293_, _18292_, _11401_);
  and _70062_ (_18294_, _18293_, _18289_);
  nor _70063_ (_18295_, _11408_, \oc8051_golden_model_1.ACC [2]);
  nor _70064_ (_18296_, _18295_, _11409_);
  and _70065_ (_18297_, _18296_, _11400_);
  or _70066_ (_18298_, _18297_, _11407_);
  or _70067_ (_18299_, _18298_, _18294_);
  nand _70068_ (_18300_, _11407_, _10334_);
  and _70069_ (_18301_, _18300_, _01442_);
  and _70070_ (_18302_, _18301_, _18299_);
  or _70071_ (_18303_, _18302_, _17989_);
  and _70072_ (_44126_, _18303_, _43634_);
  nor _70073_ (_18304_, _01442_, _10334_);
  nor _70074_ (_18305_, _11262_, _11263_);
  nor _70075_ (_18306_, _11275_, _18305_);
  and _70076_ (_18307_, _11275_, _18305_);
  or _70077_ (_18308_, _18307_, _18306_);
  and _70078_ (_18309_, _18308_, _07018_);
  or _70079_ (_18310_, _18309_, _11248_);
  and _70080_ (_18311_, _11143_, _10822_);
  nor _70081_ (_18312_, _18311_, _11144_);
  or _70082_ (_18313_, _18312_, _11127_);
  not _70083_ (_18314_, _06789_);
  or _70084_ (_18315_, _11304_, _10611_);
  or _70085_ (_18316_, _11305_, _11304_);
  nand _70086_ (_18317_, _18316_, _17457_);
  and _70087_ (_18318_, _06475_, _06501_);
  not _70088_ (_18319_, _18318_);
  and _70089_ (_18320_, _11047_, _06965_);
  and _70090_ (_18321_, _18320_, _17574_);
  and _70091_ (_18322_, _18321_, _06804_);
  and _70092_ (_18323_, _18322_, _18319_);
  nor _70093_ (_18324_, _18323_, _18305_);
  nand _70094_ (_18325_, _06269_, _06031_);
  nor _70095_ (_18326_, _08017_, _10334_);
  nor _70096_ (_18327_, _10619_, _07680_);
  or _70097_ (_18328_, _18327_, _18326_);
  or _70098_ (_18329_, _18328_, _06327_);
  and _70099_ (_18330_, _06727_, \oc8051_golden_model_1.ACC [2]);
  nor _70100_ (_18331_, _18115_, _18330_);
  nor _70101_ (_18332_, _12638_, _18331_);
  and _70102_ (_18333_, _12638_, _18331_);
  nor _70103_ (_18334_, _18333_, _18332_);
  and _70104_ (_18335_, _18119_, _18334_);
  nor _70105_ (_18336_, _18119_, _18334_);
  or _70106_ (_18337_, _18336_, _10624_);
  or _70107_ (_18338_, _18337_, _18335_);
  and _70108_ (_18339_, _06315_, _06038_);
  not _70109_ (_18340_, _18339_);
  and _70110_ (_18341_, _07854_, \oc8051_golden_model_1.ACC [2]);
  nor _70111_ (_18342_, _18068_, _18341_);
  nor _70112_ (_18343_, _18305_, _18342_);
  and _70113_ (_18344_, _18305_, _18342_);
  nor _70114_ (_18345_, _18344_, _18343_);
  and _70115_ (_18346_, _18345_, \oc8051_golden_model_1.PSW [7]);
  nor _70116_ (_18347_, _18345_, \oc8051_golden_model_1.PSW [7]);
  nor _70117_ (_18348_, _18347_, _18346_);
  and _70118_ (_18349_, _18070_, \oc8051_golden_model_1.PSW [7]);
  nor _70119_ (_18350_, _18071_, _10967_);
  nor _70120_ (_18351_, _18350_, _18349_);
  not _70121_ (_18352_, _18351_);
  and _70122_ (_18353_, _18352_, _18348_);
  nor _70123_ (_18354_, _18352_, _18348_);
  nor _70124_ (_18355_, _18354_, _18353_);
  and _70125_ (_18356_, _18355_, _18340_);
  or _70126_ (_18357_, _18356_, _10784_);
  nand _70127_ (_18358_, _10696_, _07680_);
  nor _70128_ (_18359_, _08645_, _10334_);
  and _70129_ (_18360_, _15150_, _08645_);
  or _70130_ (_18361_, _18360_, _18359_);
  or _70131_ (_18362_, _18361_, _06357_);
  and _70132_ (_18363_, _18362_, _06772_);
  and _70133_ (_18364_, _15153_, _08017_);
  or _70134_ (_18365_, _18364_, _18326_);
  and _70135_ (_18366_, _18365_, _06474_);
  nand _70136_ (_18367_, _10711_, _07680_);
  nand _70137_ (_18368_, _06855_, \oc8051_golden_model_1.ACC [3]);
  not _70138_ (_18369_, _10703_);
  or _70139_ (_18370_, _06855_, \oc8051_golden_model_1.ACC [3]);
  and _70140_ (_18371_, _18370_, _18369_);
  and _70141_ (_18372_, _18371_, _18368_);
  or _70142_ (_18373_, _18372_, _10711_);
  and _70143_ (_18374_, _18373_, _18367_);
  and _70144_ (_18375_, _18374_, _07270_);
  or _70145_ (_18376_, _18375_, _09310_);
  or _70146_ (_18377_, _18374_, _10703_);
  and _70147_ (_18378_, _18377_, _06062_);
  or _70148_ (_18379_, _18378_, _07269_);
  and _70149_ (_18380_, _18379_, _07275_);
  and _70150_ (_18381_, _18380_, _18376_);
  or _70151_ (_18382_, _18381_, _18366_);
  and _70152_ (_18383_, _18382_, _10730_);
  not _70153_ (_18384_, \oc8051_golden_model_1.PSW [6]);
  nor _70154_ (_18385_, _10732_, _18384_);
  nor _70155_ (_18386_, _18385_, \oc8051_golden_model_1.ACC [3]);
  nor _70156_ (_18387_, _18386_, _10733_);
  and _70157_ (_18388_, _18387_, _10729_);
  or _70158_ (_18389_, _18388_, _06356_);
  or _70159_ (_18390_, _18389_, _18383_);
  and _70160_ (_18391_, _18390_, _18363_);
  and _70161_ (_18392_, _18328_, _06410_);
  or _70162_ (_18393_, _18392_, _10696_);
  or _70163_ (_18394_, _18393_, _18391_);
  and _70164_ (_18395_, _18394_, _18358_);
  or _70165_ (_18396_, _18395_, _07289_);
  or _70166_ (_18397_, _09310_, _07290_);
  and _70167_ (_18398_, _18397_, _06426_);
  and _70168_ (_18399_, _18398_, _18396_);
  nor _70169_ (_18400_, _08358_, _06426_);
  or _70170_ (_18401_, _18400_, _10694_);
  or _70171_ (_18402_, _18401_, _18399_);
  nand _70172_ (_18403_, _10694_, _08688_);
  and _70173_ (_18404_, _18403_, _18402_);
  or _70174_ (_18405_, _18404_, _06352_);
  and _70175_ (_18406_, _15148_, _08645_);
  or _70176_ (_18407_, _18406_, _18359_);
  or _70177_ (_18408_, _18407_, _06353_);
  and _70178_ (_18409_, _18408_, _06346_);
  and _70179_ (_18410_, _18409_, _18405_);
  or _70180_ (_18411_, _18359_, _15180_);
  and _70181_ (_18412_, _18361_, _06345_);
  and _70182_ (_18413_, _18412_, _18411_);
  or _70183_ (_18414_, _18413_, _18410_);
  and _70184_ (_18415_, _18414_, _09612_);
  or _70185_ (_18416_, _10100_, _10098_);
  nor _70186_ (_18417_, _10101_, _09612_);
  and _70187_ (_18418_, _18417_, _18416_);
  or _70188_ (_18419_, _18418_, _14389_);
  or _70189_ (_18420_, _18419_, _18415_);
  and _70190_ (_18421_, _18420_, _18357_);
  and _70191_ (_18422_, _18355_, _18339_);
  or _70192_ (_18423_, _18422_, _10853_);
  or _70193_ (_18424_, _18423_, _18421_);
  nor _70194_ (_18425_, _09356_, _10280_);
  nor _70195_ (_18426_, _18083_, _18425_);
  nor _70196_ (_18427_, _18316_, _18426_);
  and _70197_ (_18428_, _18316_, _18426_);
  nor _70198_ (_18429_, _18428_, _18427_);
  nor _70199_ (_18430_, _18429_, _10967_);
  and _70200_ (_18431_, _18429_, _10967_);
  nor _70201_ (_18432_, _18431_, _18430_);
  and _70202_ (_18433_, _18432_, _18089_);
  nor _70203_ (_18434_, _18432_, _18089_);
  nor _70204_ (_18435_, _18434_, _18433_);
  or _70205_ (_18436_, _18435_, _10854_);
  and _70206_ (_18437_, _18436_, _06458_);
  and _70207_ (_18438_, _18437_, _18424_);
  and _70208_ (_18439_, _12625_, \oc8051_golden_model_1.PSW [7]);
  and _70209_ (_18440_, _08502_, \oc8051_golden_model_1.ACC [2]);
  nor _70210_ (_18441_, _18104_, _18440_);
  nor _70211_ (_18442_, _18441_, _12619_);
  and _70212_ (_18443_, _18441_, _12619_);
  nor _70213_ (_18444_, _18443_, _18442_);
  not _70214_ (_18445_, _12624_);
  or _70215_ (_18446_, _18445_, _18106_);
  or _70216_ (_18447_, _18446_, _10967_);
  and _70217_ (_18448_, _18447_, _18444_);
  or _70218_ (_18449_, _18448_, _10623_);
  or _70219_ (_18450_, _18449_, _18439_);
  and _70220_ (_18451_, _18450_, _12337_);
  or _70221_ (_18452_, _18451_, _18438_);
  and _70222_ (_18453_, _18452_, _18338_);
  or _70223_ (_18454_, _18453_, _06042_);
  nand _70224_ (_18455_, _06269_, _06042_);
  and _70225_ (_18456_, _18455_, _06340_);
  and _70226_ (_18457_, _18456_, _18454_);
  and _70227_ (_18458_, _15197_, _08645_);
  or _70228_ (_18459_, _18458_, _18359_);
  and _70229_ (_18460_, _18459_, _06339_);
  or _70230_ (_18461_, _18460_, _10153_);
  or _70231_ (_18462_, _18461_, _18457_);
  and _70232_ (_18463_, _18462_, _18329_);
  or _70233_ (_18464_, _18463_, _09572_);
  and _70234_ (_18465_, _09310_, _08017_);
  or _70235_ (_18466_, _18326_, _06333_);
  or _70236_ (_18467_, _18466_, _18465_);
  and _70237_ (_18468_, _18467_, _06313_);
  and _70238_ (_18469_, _18468_, _18464_);
  and _70239_ (_18470_, _15251_, _08017_);
  or _70240_ (_18471_, _18470_, _18326_);
  and _70241_ (_18472_, _18471_, _06037_);
  or _70242_ (_18473_, _18472_, _10166_);
  or _70243_ (_18474_, _18473_, _18469_);
  or _70244_ (_18475_, _10302_, _10172_);
  and _70245_ (_18476_, _18475_, _18474_);
  or _70246_ (_18477_, _18476_, _06031_);
  and _70247_ (_18478_, _18477_, _18325_);
  or _70248_ (_18479_, _18478_, _06277_);
  and _70249_ (_18480_, _08017_, _09014_);
  or _70250_ (_18481_, _18480_, _18326_);
  or _70251_ (_18482_, _18481_, _06278_);
  and _70252_ (_18483_, _18482_, _11029_);
  nand _70253_ (_18484_, _18483_, _18479_);
  or _70254_ (_18485_, _11029_, _06269_);
  and _70255_ (_18486_, _18485_, _18323_);
  and _70256_ (_18487_, _18486_, _18484_);
  or _70257_ (_18488_, _18487_, _18324_);
  and _70258_ (_18489_, _18488_, _17570_);
  nor _70259_ (_18490_, _18305_, _17570_);
  or _70260_ (_18491_, _18490_, _17572_);
  nor _70261_ (_18492_, _18491_, _18489_);
  nand _70262_ (_18493_, _18316_, _06028_);
  and _70263_ (_18494_, _18493_, _11052_);
  or _70264_ (_18495_, _18494_, _18492_);
  and _70265_ (_18496_, _18495_, _18317_);
  or _70266_ (_18497_, _18496_, _06613_);
  or _70267_ (_18498_, _12619_, _06614_);
  and _70268_ (_18499_, _18498_, _11071_);
  and _70269_ (_18500_, _18499_, _18497_);
  and _70270_ (_18501_, _11064_, _12638_);
  or _70271_ (_18502_, _18501_, _06502_);
  or _70272_ (_18503_, _18502_, _18500_);
  and _70273_ (_18504_, _15266_, _08017_);
  or _70274_ (_18505_, _18504_, _18326_);
  or _70275_ (_18506_, _18505_, _07334_);
  and _70276_ (_18507_, _18506_, _18503_);
  or _70277_ (_18508_, _18507_, _06615_);
  or _70278_ (_18509_, _18326_, _07337_);
  and _70279_ (_18510_, _18509_, _17595_);
  and _70280_ (_18511_, _18510_, _18508_);
  and _70281_ (_18512_, _17598_, _11262_);
  or _70282_ (_18513_, _18512_, _06976_);
  or _70283_ (_18514_, _18513_, _18511_);
  and _70284_ (_18515_, _18514_, _18315_);
  or _70285_ (_18516_, _18515_, _06608_);
  or _70286_ (_18517_, _10573_, _06609_);
  and _70287_ (_18518_, _18517_, _11090_);
  and _70288_ (_18519_, _18518_, _18516_);
  and _70289_ (_18520_, _11089_, _11345_);
  or _70290_ (_18521_, _18520_, _18519_);
  and _70291_ (_18522_, _18521_, _07339_);
  nand _70292_ (_18523_, _18481_, _06507_);
  nor _70293_ (_18524_, _18523_, _10574_);
  or _70294_ (_18525_, _18524_, _18522_);
  and _70295_ (_18526_, _18525_, _18314_);
  nor _70296_ (_18527_, _11263_, _18314_);
  nor _70297_ (_18528_, _06323_, _06792_);
  nor _70298_ (_18529_, _18528_, _06022_);
  or _70299_ (_18530_, _18529_, _18527_);
  or _70300_ (_18531_, _18530_, _18526_);
  nand _70301_ (_18532_, _18529_, _11263_);
  and _70302_ (_18533_, _18532_, _18207_);
  and _70303_ (_18534_, _18533_, _18531_);
  nor _70304_ (_18535_, _18207_, _11263_);
  or _70305_ (_18536_, _18535_, _06987_);
  or _70306_ (_18537_, _18536_, _18534_);
  nand _70307_ (_18538_, _11305_, _06987_);
  and _70308_ (_18539_, _18538_, _06605_);
  and _70309_ (_18540_, _18539_, _18537_);
  nand _70310_ (_18541_, _17625_, _10574_);
  and _70311_ (_18542_, _18541_, _12315_);
  or _70312_ (_18543_, _18542_, _18540_);
  nand _70313_ (_18544_, _11114_, _11346_);
  and _70314_ (_18545_, _18544_, _09107_);
  and _70315_ (_18546_, _18545_, _18543_);
  and _70316_ (_18547_, _15263_, _08017_);
  or _70317_ (_18548_, _18547_, _18326_);
  and _70318_ (_18549_, _18548_, _06509_);
  or _70319_ (_18550_, _18549_, _11130_);
  or _70320_ (_18551_, _18550_, _18546_);
  and _70321_ (_18552_, _18551_, _18313_);
  or _70322_ (_18553_, _18552_, _11129_);
  and _70323_ (_18554_, _11171_, _10888_);
  nor _70324_ (_18555_, _18554_, _11172_);
  or _70325_ (_18556_, _18555_, _11158_);
  and _70326_ (_18557_, _18556_, _06601_);
  and _70327_ (_18558_, _18557_, _18553_);
  and _70328_ (_18559_, _11201_, _10658_);
  nor _70329_ (_18560_, _18559_, _11202_);
  or _70330_ (_18561_, _18560_, _11186_);
  and _70331_ (_18562_, _18561_, _11188_);
  or _70332_ (_18563_, _18562_, _18558_);
  and _70333_ (_18564_, _11230_, _10959_);
  nor _70334_ (_18565_, _18564_, _11231_);
  or _70335_ (_18566_, _18565_, _11218_);
  and _70336_ (_18567_, _18566_, _11217_);
  and _70337_ (_18568_, _18567_, _18563_);
  and _70338_ (_18569_, _11216_, \oc8051_golden_model_1.ACC [2]);
  or _70339_ (_18570_, _18569_, _17444_);
  or _70340_ (_18571_, _18570_, _18568_);
  and _70341_ (_18572_, _18571_, _18310_);
  and _70342_ (_18573_, _18308_, _07017_);
  or _70343_ (_18574_, _18573_, _11290_);
  or _70344_ (_18575_, _18574_, _18572_);
  not _70345_ (_18576_, _11318_);
  nor _70346_ (_18577_, _18576_, _18316_);
  and _70347_ (_18578_, _18576_, _18316_);
  or _70348_ (_18579_, _18578_, _18577_);
  or _70349_ (_18580_, _18579_, _11292_);
  and _70350_ (_18581_, _18580_, _06364_);
  and _70351_ (_18582_, _18581_, _18575_);
  and _70352_ (_18583_, _12619_, _10586_);
  nor _70353_ (_18584_, _12619_, _10586_);
  or _70354_ (_18585_, _18584_, _18583_);
  and _70355_ (_18586_, _18585_, _06363_);
  or _70356_ (_18587_, _18586_, _10566_);
  or _70357_ (_18588_, _18587_, _18582_);
  and _70358_ (_18589_, _11360_, _12638_);
  nor _70359_ (_18590_, _11360_, _12638_);
  or _70360_ (_18591_, _18590_, _18589_);
  or _70361_ (_18592_, _18591_, _10567_);
  and _70362_ (_18593_, _18592_, _13049_);
  and _70363_ (_18594_, _18593_, _18588_);
  and _70364_ (_18595_, _10564_, \oc8051_golden_model_1.ACC [2]);
  or _70365_ (_18596_, _18595_, _06639_);
  or _70366_ (_18597_, _18596_, _18594_);
  or _70367_ (_18598_, _18365_, _07048_);
  and _70368_ (_18599_, _18598_, _11378_);
  and _70369_ (_18600_, _18599_, _18597_);
  nor _70370_ (_18601_, _11383_, _10334_);
  or _70371_ (_18602_, _18601_, _11384_);
  nor _70372_ (_18603_, _18602_, _11382_);
  nor _70373_ (_18604_, _18603_, _13072_);
  or _70374_ (_18605_, _18604_, _18600_);
  nand _70375_ (_18606_, _11382_, _10204_);
  and _70376_ (_18607_, _18606_, _05990_);
  and _70377_ (_18608_, _18607_, _18605_);
  and _70378_ (_18609_, _18407_, _05989_);
  or _70379_ (_18610_, _18609_, _06646_);
  or _70380_ (_18611_, _18610_, _18608_);
  and _70381_ (_18612_, _15321_, _08017_);
  or _70382_ (_18613_, _18326_, _06651_);
  or _70383_ (_18614_, _18613_, _18612_);
  and _70384_ (_18615_, _18614_, _11401_);
  and _70385_ (_18616_, _18615_, _18611_);
  nor _70386_ (_18617_, _11409_, \oc8051_golden_model_1.ACC [3]);
  nor _70387_ (_18618_, _18617_, _11410_);
  and _70388_ (_18619_, _18618_, _11400_);
  or _70389_ (_18620_, _18619_, _11407_);
  or _70390_ (_18621_, _18620_, _18616_);
  nand _70391_ (_18622_, _11407_, _10204_);
  and _70392_ (_18623_, _18622_, _01442_);
  and _70393_ (_18624_, _18623_, _18621_);
  or _70394_ (_18625_, _18624_, _18304_);
  and _70395_ (_44127_, _18625_, _43634_);
  nor _70396_ (_18626_, _01442_, _10204_);
  or _70397_ (_18627_, _10590_, _10588_);
  and _70398_ (_18628_, _10591_, _06363_);
  and _70399_ (_18629_, _18628_, _18627_);
  or _70400_ (_18630_, _11320_, _11303_);
  and _70401_ (_18631_, _18630_, _11321_);
  or _70402_ (_18632_, _18631_, _17691_);
  or _70403_ (_18633_, _11145_, _10816_);
  and _70404_ (_18634_, _18633_, _11146_);
  and _70405_ (_18635_, _18634_, _11130_);
  nand _70406_ (_18636_, _11114_, _11343_);
  or _70407_ (_18637_, _11260_, _17452_);
  or _70408_ (_18638_, _10571_, _06609_);
  and _70409_ (_18639_, _18638_, _11090_);
  and _70410_ (_18640_, _15345_, _08017_);
  nor _70411_ (_18641_, _08017_, _10204_);
  or _70412_ (_18642_, _18641_, _07334_);
  or _70413_ (_18643_, _18642_, _18640_);
  or _70414_ (_18644_, _11060_, _11303_);
  nor _70415_ (_18645_, _11046_, _06802_);
  not _70416_ (_18646_, _18645_);
  or _70417_ (_18647_, _11040_, _11261_);
  nand _70418_ (_18648_, _07093_, _06031_);
  nor _70419_ (_18649_, _08596_, _10619_);
  or _70420_ (_18650_, _18649_, _18641_);
  or _70421_ (_18651_, _18650_, _06327_);
  nor _70422_ (_18652_, _12643_, _10967_);
  or _70423_ (_18653_, _18331_, _14363_);
  and _70424_ (_18654_, _18653_, _14362_);
  nor _70425_ (_18655_, _11344_, _18654_);
  and _70426_ (_18656_, _11344_, _18654_);
  nor _70427_ (_18657_, _18656_, _18655_);
  and _70428_ (_18658_, _18657_, \oc8051_golden_model_1.PSW [7]);
  nor _70429_ (_18659_, _18657_, \oc8051_golden_model_1.PSW [7]);
  nor _70430_ (_18660_, _18659_, _18658_);
  and _70431_ (_18661_, _18660_, _18652_);
  nor _70432_ (_18662_, _18660_, _18652_);
  nor _70433_ (_18663_, _18662_, _18661_);
  or _70434_ (_18664_, _18663_, _10624_);
  or _70435_ (_18665_, _18433_, _18430_);
  or _70436_ (_18666_, _09310_, _10334_);
  and _70437_ (_18667_, _09310_, _10334_);
  or _70438_ (_18668_, _18426_, _18667_);
  and _70439_ (_18669_, _18668_, _18666_);
  nor _70440_ (_18670_, _11303_, _18669_);
  and _70441_ (_18671_, _11303_, _18669_);
  nor _70442_ (_18672_, _18671_, _18670_);
  and _70443_ (_18673_, _18672_, \oc8051_golden_model_1.PSW [7]);
  nor _70444_ (_18674_, _18672_, \oc8051_golden_model_1.PSW [7]);
  nor _70445_ (_18675_, _18674_, _18673_);
  or _70446_ (_18676_, _18675_, _18665_);
  and _70447_ (_18677_, _18675_, _18665_);
  nor _70448_ (_18678_, _18677_, _10854_);
  and _70449_ (_18679_, _18678_, _18676_);
  or _70450_ (_18680_, _18353_, _18346_);
  nor _70451_ (_18681_, _07680_, \oc8051_golden_model_1.ACC [3]);
  nand _70452_ (_18682_, _07680_, \oc8051_golden_model_1.ACC [3]);
  and _70453_ (_18683_, _18682_, _18342_);
  or _70454_ (_18684_, _18683_, _18681_);
  nor _70455_ (_18685_, _11261_, _18684_);
  and _70456_ (_18686_, _11261_, _18684_);
  nor _70457_ (_18687_, _18686_, _18685_);
  and _70458_ (_18688_, _18687_, \oc8051_golden_model_1.PSW [7]);
  nor _70459_ (_18689_, _18687_, \oc8051_golden_model_1.PSW [7]);
  nor _70460_ (_18690_, _18689_, _18688_);
  or _70461_ (_18691_, _18690_, _18680_);
  and _70462_ (_18692_, _18690_, _18680_);
  nor _70463_ (_18693_, _18692_, _10784_);
  and _70464_ (_18694_, _18693_, _18691_);
  nand _70465_ (_18695_, _10696_, _08596_);
  nor _70466_ (_18696_, _08645_, _10204_);
  and _70467_ (_18697_, _15353_, _08645_);
  or _70468_ (_18698_, _18697_, _18696_);
  or _70469_ (_18699_, _18698_, _06357_);
  and _70470_ (_18700_, _18699_, _06772_);
  nand _70471_ (_18701_, _10711_, _08596_);
  nand _70472_ (_18702_, _06855_, \oc8051_golden_model_1.ACC [4]);
  or _70473_ (_18703_, _06855_, \oc8051_golden_model_1.ACC [4]);
  and _70474_ (_18704_, _18703_, _18369_);
  and _70475_ (_18705_, _18704_, _18702_);
  or _70476_ (_18706_, _18705_, _10711_);
  and _70477_ (_18707_, _18706_, _18701_);
  and _70478_ (_18708_, _10703_, _09264_);
  or _70479_ (_18709_, _18708_, _18707_);
  and _70480_ (_18710_, _18709_, _10722_);
  and _70481_ (_18711_, _15367_, _08017_);
  or _70482_ (_18712_, _18711_, _18641_);
  and _70483_ (_18713_, _18712_, _06474_);
  or _70484_ (_18714_, _18713_, _18710_);
  and _70485_ (_18715_, _18714_, _10730_);
  nor _70486_ (_18716_, _10733_, \oc8051_golden_model_1.ACC [4]);
  nor _70487_ (_18717_, _18716_, _10734_);
  and _70488_ (_18718_, _18717_, _10729_);
  or _70489_ (_18719_, _18718_, _06356_);
  or _70490_ (_18720_, _18719_, _18715_);
  and _70491_ (_18721_, _18720_, _18700_);
  and _70492_ (_18722_, _18650_, _06410_);
  or _70493_ (_18723_, _18722_, _10696_);
  or _70494_ (_18724_, _18723_, _18721_);
  and _70495_ (_18725_, _18724_, _18695_);
  or _70496_ (_18726_, _18725_, _07289_);
  or _70497_ (_18727_, _09264_, _07290_);
  and _70498_ (_18728_, _18727_, _06426_);
  and _70499_ (_18729_, _18728_, _18726_);
  nor _70500_ (_18730_, _08598_, _06426_);
  or _70501_ (_18731_, _18730_, _10694_);
  or _70502_ (_18732_, _18731_, _18729_);
  nand _70503_ (_18733_, _10694_, _06071_);
  and _70504_ (_18734_, _18733_, _18732_);
  or _70505_ (_18735_, _18734_, _06352_);
  and _70506_ (_18736_, _15348_, _08645_);
  or _70507_ (_18737_, _18736_, _18696_);
  or _70508_ (_18738_, _18737_, _06353_);
  and _70509_ (_18739_, _18738_, _06346_);
  and _70510_ (_18740_, _18739_, _18735_);
  or _70511_ (_18741_, _18696_, _15384_);
  and _70512_ (_18742_, _18698_, _06345_);
  and _70513_ (_18743_, _18742_, _18741_);
  or _70514_ (_18744_, _18743_, _09606_);
  or _70515_ (_18745_, _18744_, _18740_);
  nor _70516_ (_18746_, _10103_, _10101_);
  nor _70517_ (_18747_, _18746_, _10104_);
  or _70518_ (_18748_, _18747_, _09612_);
  and _70519_ (_18749_, _18748_, _10784_);
  and _70520_ (_18750_, _18749_, _18745_);
  or _70521_ (_18751_, _18750_, _18694_);
  and _70522_ (_18752_, _18751_, _10854_);
  or _70523_ (_18753_, _18752_, _18679_);
  and _70524_ (_18754_, _18753_, _06458_);
  nor _70525_ (_18755_, _12625_, _10967_);
  or _70526_ (_18756_, _18441_, _14321_);
  and _70527_ (_18757_, _18756_, _14319_);
  nor _70528_ (_18758_, _18757_, _10590_);
  and _70529_ (_18759_, _18757_, _10590_);
  nor _70530_ (_18760_, _18759_, _18758_);
  and _70531_ (_18761_, _18760_, \oc8051_golden_model_1.PSW [7]);
  nor _70532_ (_18762_, _18760_, \oc8051_golden_model_1.PSW [7]);
  nor _70533_ (_18763_, _18762_, _18761_);
  or _70534_ (_18764_, _18763_, _18755_);
  and _70535_ (_18765_, _18763_, _18755_);
  nor _70536_ (_18766_, _18765_, _06458_);
  and _70537_ (_18767_, _18766_, _18764_);
  or _70538_ (_18768_, _18767_, _10623_);
  or _70539_ (_18769_, _18768_, _18754_);
  and _70540_ (_18770_, _18769_, _18664_);
  or _70541_ (_18771_, _18770_, _06042_);
  nand _70542_ (_18772_, _07093_, _06042_);
  and _70543_ (_18773_, _18772_, _06340_);
  and _70544_ (_18774_, _18773_, _18771_);
  and _70545_ (_18775_, _15350_, _08645_);
  or _70546_ (_18776_, _18775_, _18696_);
  and _70547_ (_18777_, _18776_, _06339_);
  or _70548_ (_18778_, _18777_, _10153_);
  or _70549_ (_18779_, _18778_, _18774_);
  and _70550_ (_18780_, _18779_, _18651_);
  or _70551_ (_18781_, _18780_, _09572_);
  and _70552_ (_18782_, _09264_, _08017_);
  or _70553_ (_18783_, _18641_, _06333_);
  or _70554_ (_18784_, _18783_, _18782_);
  and _70555_ (_18785_, _18784_, _06313_);
  and _70556_ (_18786_, _18785_, _18781_);
  and _70557_ (_18787_, _15452_, _08017_);
  or _70558_ (_18788_, _18787_, _18641_);
  and _70559_ (_18789_, _18788_, _06037_);
  or _70560_ (_18790_, _18789_, _10166_);
  or _70561_ (_18791_, _18790_, _18786_);
  or _70562_ (_18792_, _10249_, _10172_);
  and _70563_ (_18793_, _18792_, _18791_);
  or _70564_ (_18794_, _18793_, _06031_);
  and _70565_ (_18795_, _18794_, _18648_);
  or _70566_ (_18796_, _18795_, _06277_);
  and _70567_ (_18797_, _08995_, _08017_);
  or _70568_ (_18798_, _18797_, _18641_);
  or _70569_ (_18799_, _18798_, _06278_);
  and _70570_ (_18800_, _18799_, _11029_);
  and _70571_ (_18801_, _18800_, _18796_);
  nor _70572_ (_18802_, _11029_, _07093_);
  or _70573_ (_18803_, _18802_, _11036_);
  or _70574_ (_18804_, _18803_, _18801_);
  and _70575_ (_18805_, _18804_, _18647_);
  or _70576_ (_18806_, _18805_, _18646_);
  nor _70577_ (_18807_, _10708_, _06011_);
  nor _70578_ (_18808_, _18645_, _11261_);
  nor _70579_ (_18809_, _18808_, _18807_);
  and _70580_ (_18810_, _18809_, _18806_);
  and _70581_ (_18811_, _18807_, _11261_);
  or _70582_ (_18812_, _18811_, _11052_);
  or _70583_ (_18813_, _18812_, _18810_);
  and _70584_ (_18814_, _18813_, _18644_);
  or _70585_ (_18815_, _18814_, _06613_);
  or _70586_ (_18816_, _10590_, _06614_);
  and _70587_ (_18817_, _18816_, _11071_);
  and _70588_ (_18818_, _18817_, _18815_);
  and _70589_ (_18819_, _11064_, _11344_);
  or _70590_ (_18820_, _18819_, _06502_);
  or _70591_ (_18821_, _18820_, _18818_);
  and _70592_ (_18822_, _18821_, _18643_);
  or _70593_ (_18823_, _18822_, _06615_);
  or _70594_ (_18824_, _18641_, _07337_);
  and _70595_ (_18825_, _17857_, _17855_);
  and _70596_ (_18826_, _18825_, _18824_);
  and _70597_ (_18827_, _18826_, _18823_);
  nor _70598_ (_18828_, _18825_, _11259_);
  or _70599_ (_18829_, _18828_, _17863_);
  or _70600_ (_18830_, _18829_, _18827_);
  or _70601_ (_18831_, _17869_, _11258_);
  and _70602_ (_18832_, _18831_, _10611_);
  and _70603_ (_18833_, _18832_, _18830_);
  and _70604_ (_18834_, _11300_, _06976_);
  or _70605_ (_18835_, _18834_, _06608_);
  or _70606_ (_18836_, _18835_, _18833_);
  and _70607_ (_18837_, _18836_, _18639_);
  and _70608_ (_18838_, _11089_, _11341_);
  or _70609_ (_18839_, _18838_, _18837_);
  and _70610_ (_18840_, _18839_, _07339_);
  nand _70611_ (_18841_, _18798_, _06507_);
  nor _70612_ (_18842_, _18841_, _10589_);
  or _70613_ (_18843_, _18842_, _10609_);
  or _70614_ (_18844_, _18843_, _18840_);
  and _70615_ (_18845_, _18844_, _18637_);
  or _70616_ (_18846_, _18845_, _11102_);
  and _70617_ (_18847_, _11260_, _06985_);
  or _70618_ (_18848_, _18847_, _11104_);
  and _70619_ (_18849_, _18848_, _18846_);
  and _70620_ (_18850_, _11260_, _06984_);
  or _70621_ (_18851_, _18850_, _06987_);
  or _70622_ (_18852_, _18851_, _18849_);
  not _70623_ (_18853_, _06987_);
  or _70624_ (_18854_, _11302_, _18853_);
  and _70625_ (_18855_, _18854_, _06605_);
  and _70626_ (_18856_, _18855_, _18852_);
  nand _70627_ (_18857_, _17625_, _10589_);
  and _70628_ (_18858_, _18857_, _12315_);
  or _70629_ (_18859_, _18858_, _18856_);
  and _70630_ (_18860_, _18859_, _18636_);
  or _70631_ (_18861_, _18860_, _06509_);
  and _70632_ (_18862_, _15342_, _08017_);
  or _70633_ (_18863_, _18641_, _09107_);
  or _70634_ (_18864_, _18863_, _18862_);
  and _70635_ (_18865_, _18864_, _11127_);
  and _70636_ (_18866_, _18865_, _18861_);
  or _70637_ (_18867_, _18866_, _18635_);
  and _70638_ (_18868_, _18867_, _18231_);
  or _70639_ (_18869_, _11173_, _10881_);
  and _70640_ (_18870_, _18869_, _11174_);
  and _70641_ (_18871_, _18870_, _17922_);
  or _70642_ (_18872_, _18871_, _07002_);
  or _70643_ (_18873_, _18872_, _18868_);
  or _70644_ (_18874_, _18870_, _18237_);
  and _70645_ (_18875_, _18874_, _06601_);
  and _70646_ (_18876_, _18875_, _18873_);
  or _70647_ (_18877_, _11203_, _10651_);
  and _70648_ (_18878_, _18877_, _11204_);
  or _70649_ (_18879_, _18878_, _11186_);
  and _70650_ (_18880_, _18879_, _11188_);
  or _70651_ (_18881_, _18880_, _18876_);
  or _70652_ (_18882_, _11232_, _11222_);
  and _70653_ (_18883_, _18882_, _11233_);
  or _70654_ (_18884_, _18883_, _11218_);
  and _70655_ (_18885_, _18884_, _18881_);
  or _70656_ (_18886_, _18885_, _11216_);
  nand _70657_ (_18887_, _11216_, _10334_);
  and _70658_ (_18888_, _18887_, _11248_);
  and _70659_ (_18889_, _18888_, _18886_);
  nor _70660_ (_18890_, _11277_, _11261_);
  nor _70661_ (_18891_, _18890_, _11278_);
  and _70662_ (_18892_, _18891_, _18254_);
  or _70663_ (_18893_, _18892_, _17690_);
  or _70664_ (_18894_, _18893_, _18889_);
  and _70665_ (_18895_, _18894_, _18632_);
  or _70666_ (_18896_, _18895_, _07019_);
  or _70667_ (_18897_, _18631_, _07020_);
  and _70668_ (_18898_, _18897_, _06364_);
  and _70669_ (_18899_, _18898_, _18896_);
  or _70670_ (_18900_, _18899_, _18629_);
  and _70671_ (_18901_, _18900_, _10567_);
  or _70672_ (_18902_, _11362_, _11344_);
  and _70673_ (_18903_, _18902_, _11363_);
  and _70674_ (_18904_, _18903_, _10566_);
  or _70675_ (_18905_, _18904_, _18901_);
  and _70676_ (_18906_, _18905_, _13049_);
  and _70677_ (_18907_, _10564_, \oc8051_golden_model_1.ACC [3]);
  or _70678_ (_18908_, _18907_, _06639_);
  or _70679_ (_18909_, _18908_, _18906_);
  or _70680_ (_18910_, _18712_, _07048_);
  and _70681_ (_18911_, _18910_, _11378_);
  and _70682_ (_18912_, _18911_, _18909_);
  nor _70683_ (_18913_, _11384_, _10204_);
  or _70684_ (_18914_, _18913_, _11385_);
  and _70685_ (_18915_, _18914_, _11377_);
  or _70686_ (_18916_, _18915_, _11382_);
  or _70687_ (_18917_, _18916_, _18912_);
  nand _70688_ (_18918_, _11382_, _10237_);
  and _70689_ (_18919_, _18918_, _05990_);
  and _70690_ (_18920_, _18919_, _18917_);
  and _70691_ (_18921_, _18737_, _05989_);
  or _70692_ (_18922_, _18921_, _06646_);
  or _70693_ (_18923_, _18922_, _18920_);
  and _70694_ (_18924_, _15524_, _08017_);
  or _70695_ (_18925_, _18641_, _06651_);
  or _70696_ (_18926_, _18925_, _18924_);
  and _70697_ (_18927_, _18926_, _11401_);
  and _70698_ (_18928_, _18927_, _18923_);
  nor _70699_ (_18929_, _11410_, \oc8051_golden_model_1.ACC [4]);
  nor _70700_ (_18930_, _18929_, _11411_);
  and _70701_ (_18931_, _18930_, _11400_);
  or _70702_ (_18932_, _18931_, _11407_);
  or _70703_ (_18933_, _18932_, _18928_);
  nand _70704_ (_18934_, _11407_, _10237_);
  and _70705_ (_18935_, _18934_, _01442_);
  and _70706_ (_18936_, _18935_, _18933_);
  or _70707_ (_18937_, _18936_, _18626_);
  and _70708_ (_44128_, _18937_, _43634_);
  nor _70709_ (_18938_, _01442_, _10237_);
  and _70710_ (_18939_, _11147_, _10813_);
  nor _70711_ (_18940_, _18939_, _11148_);
  or _70712_ (_18941_, _18940_, _11127_);
  nor _70713_ (_18942_, _11256_, _06984_);
  or _70714_ (_18943_, _18942_, _11104_);
  and _70715_ (_18944_, _11255_, _10617_);
  and _70716_ (_18945_, _15664_, _08017_);
  nor _70717_ (_18946_, _08017_, _10237_);
  or _70718_ (_18947_, _18946_, _07334_);
  or _70719_ (_18948_, _18947_, _18945_);
  or _70720_ (_18949_, _12626_, _06614_);
  and _70721_ (_18950_, _18949_, _11071_);
  nor _70722_ (_18951_, _18807_, _11046_);
  not _70723_ (_18952_, _18951_);
  and _70724_ (_18953_, _18952_, _11257_);
  not _70725_ (_18954_, _06803_);
  and _70726_ (_18955_, _11257_, _06964_);
  nand _70727_ (_18956_, _06685_, _06031_);
  nor _70728_ (_18957_, _08305_, _10619_);
  or _70729_ (_18958_, _18957_, _18946_);
  or _70730_ (_18959_, _18958_, _06327_);
  and _70731_ (_18960_, _07093_, \oc8051_golden_model_1.ACC [4]);
  nor _70732_ (_18961_, _18655_, _18960_);
  nor _70733_ (_18962_, _12644_, _18961_);
  and _70734_ (_18963_, _12644_, _18961_);
  nor _70735_ (_18964_, _18963_, _18962_);
  and _70736_ (_18965_, _18964_, \oc8051_golden_model_1.PSW [7]);
  nor _70737_ (_18966_, _18964_, \oc8051_golden_model_1.PSW [7]);
  nor _70738_ (_18967_, _18966_, _18965_);
  nor _70739_ (_18968_, _18661_, _18658_);
  not _70740_ (_18969_, _18968_);
  and _70741_ (_18970_, _18969_, _18967_);
  nor _70742_ (_18971_, _18969_, _18967_);
  nor _70743_ (_18972_, _18971_, _18970_);
  or _70744_ (_18973_, _18972_, _10624_);
  nand _70745_ (_18974_, _10696_, _08305_);
  and _70746_ (_18975_, _10703_, _09218_);
  nor _70747_ (_18976_, _10712_, _08305_);
  nor _70748_ (_18977_, _06855_, _10237_);
  and _70749_ (_18978_, _06855_, _10237_);
  or _70750_ (_18979_, _18978_, _18977_);
  and _70751_ (_18980_, _18979_, _10714_);
  or _70752_ (_18981_, _18980_, _18976_);
  or _70753_ (_18982_, _18981_, _18975_);
  and _70754_ (_18983_, _18982_, _10722_);
  and _70755_ (_18984_, _15550_, _08017_);
  or _70756_ (_18985_, _18984_, _18946_);
  and _70757_ (_18986_, _18985_, _06474_);
  or _70758_ (_18987_, _18986_, _10729_);
  or _70759_ (_18988_, _18987_, _18983_);
  nor _70760_ (_18989_, _10750_, _10742_);
  nand _70761_ (_18990_, _10750_, _10742_);
  nand _70762_ (_18991_, _18990_, _10729_);
  or _70763_ (_18992_, _18991_, _18989_);
  and _70764_ (_18993_, _18992_, _06418_);
  and _70765_ (_18994_, _18993_, _18988_);
  nor _70766_ (_18995_, _08645_, _10237_);
  and _70767_ (_18996_, _15566_, _08645_);
  or _70768_ (_18997_, _18996_, _18995_);
  and _70769_ (_18998_, _18997_, _06356_);
  and _70770_ (_18999_, _18958_, _06410_);
  or _70771_ (_19000_, _18999_, _10696_);
  or _70772_ (_19001_, _19000_, _18998_);
  or _70773_ (_19002_, _19001_, _18994_);
  and _70774_ (_19003_, _19002_, _18974_);
  or _70775_ (_19004_, _19003_, _07289_);
  or _70776_ (_19005_, _09218_, _07290_);
  and _70777_ (_19006_, _19005_, _06426_);
  and _70778_ (_19007_, _19006_, _19004_);
  nor _70779_ (_19008_, _08307_, _06426_);
  or _70780_ (_19009_, _19008_, _10694_);
  or _70781_ (_19010_, _19009_, _19007_);
  nand _70782_ (_19011_, _10694_, _06097_);
  and _70783_ (_19012_, _19011_, _19010_);
  or _70784_ (_19013_, _19012_, _06352_);
  and _70785_ (_19014_, _15544_, _08645_);
  or _70786_ (_19015_, _19014_, _18995_);
  or _70787_ (_19016_, _19015_, _06353_);
  and _70788_ (_19017_, _19016_, _06346_);
  and _70789_ (_19018_, _19017_, _19013_);
  or _70790_ (_19019_, _18995_, _15581_);
  and _70791_ (_19020_, _18997_, _06345_);
  and _70792_ (_19021_, _19020_, _19019_);
  or _70793_ (_19022_, _19021_, _19018_);
  and _70794_ (_19023_, _19022_, _09612_);
  or _70795_ (_19024_, _10106_, _10104_);
  nor _70796_ (_19025_, _10107_, _09612_);
  and _70797_ (_19026_, _19025_, _19024_);
  or _70798_ (_19027_, _19026_, _12338_);
  or _70799_ (_19028_, _19027_, _19023_);
  and _70800_ (_19029_, _08596_, \oc8051_golden_model_1.ACC [4]);
  nor _70801_ (_19030_, _18685_, _19029_);
  nor _70802_ (_19031_, _11257_, _19030_);
  and _70803_ (_19032_, _11257_, _19030_);
  nor _70804_ (_19033_, _19032_, _19031_);
  and _70805_ (_19034_, _19033_, \oc8051_golden_model_1.PSW [7]);
  nor _70806_ (_19035_, _19033_, \oc8051_golden_model_1.PSW [7]);
  nor _70807_ (_19036_, _19035_, _19034_);
  nor _70808_ (_19037_, _18692_, _18688_);
  not _70809_ (_19038_, _19037_);
  and _70810_ (_19039_, _19038_, _19036_);
  nor _70811_ (_19040_, _19038_, _19036_);
  nor _70812_ (_19041_, _19040_, _19039_);
  or _70813_ (_19042_, _19041_, _10784_);
  and _70814_ (_19043_, _19042_, _19028_);
  or _70815_ (_19044_, _19043_, _10853_);
  nor _70816_ (_19045_, _09264_, _10204_);
  nor _70817_ (_19046_, _18670_, _19045_);
  nor _70818_ (_19047_, _11299_, _19046_);
  and _70819_ (_19048_, _11299_, _19046_);
  nor _70820_ (_19049_, _19048_, _19047_);
  nor _70821_ (_19050_, _19049_, _10967_);
  and _70822_ (_19051_, _19049_, _10967_);
  nor _70823_ (_19052_, _19051_, _19050_);
  nor _70824_ (_19053_, _18677_, _18673_);
  not _70825_ (_19054_, _19053_);
  and _70826_ (_19055_, _19054_, _19052_);
  nor _70827_ (_19056_, _19054_, _19052_);
  nor _70828_ (_19057_, _19056_, _19055_);
  or _70829_ (_19058_, _19057_, _10854_);
  and _70830_ (_19059_, _19058_, _06458_);
  and _70831_ (_19060_, _19059_, _19044_);
  and _70832_ (_19061_, _08598_, \oc8051_golden_model_1.ACC [4]);
  nor _70833_ (_19062_, _18758_, _19061_);
  nor _70834_ (_19063_, _19062_, _12626_);
  and _70835_ (_19064_, _19062_, _12626_);
  nor _70836_ (_19065_, _19064_, _19063_);
  and _70837_ (_19066_, _19065_, \oc8051_golden_model_1.PSW [7]);
  nor _70838_ (_19067_, _19065_, \oc8051_golden_model_1.PSW [7]);
  nor _70839_ (_19068_, _19067_, _19066_);
  nor _70840_ (_19069_, _18765_, _18761_);
  not _70841_ (_19070_, _19069_);
  and _70842_ (_19071_, _19070_, _19068_);
  nor _70843_ (_19072_, _19070_, _19068_);
  nor _70844_ (_19073_, _19072_, _19071_);
  or _70845_ (_19074_, _19073_, _10623_);
  and _70846_ (_19075_, _19074_, _12337_);
  or _70847_ (_19076_, _19075_, _19060_);
  and _70848_ (_19077_, _19076_, _18973_);
  or _70849_ (_19078_, _19077_, _06042_);
  nand _70850_ (_19079_, _06685_, _06042_);
  and _70851_ (_19080_, _19079_, _06340_);
  and _70852_ (_19081_, _19080_, _19078_);
  and _70853_ (_19082_, _15546_, _08645_);
  or _70854_ (_19083_, _19082_, _18995_);
  and _70855_ (_19084_, _19083_, _06339_);
  or _70856_ (_19085_, _19084_, _10153_);
  or _70857_ (_19086_, _19085_, _19081_);
  and _70858_ (_19087_, _19086_, _18959_);
  or _70859_ (_19088_, _19087_, _09572_);
  and _70860_ (_19089_, _09218_, _08017_);
  or _70861_ (_19090_, _18946_, _06333_);
  or _70862_ (_19091_, _19090_, _19089_);
  and _70863_ (_19092_, _19091_, _06313_);
  and _70864_ (_19093_, _19092_, _19088_);
  and _70865_ (_19094_, _15649_, _08017_);
  or _70866_ (_19095_, _19094_, _18946_);
  and _70867_ (_19096_, _19095_, _06037_);
  or _70868_ (_19097_, _19096_, _10166_);
  or _70869_ (_19098_, _19097_, _19093_);
  or _70870_ (_19099_, _10222_, _10172_);
  and _70871_ (_19100_, _19099_, _19098_);
  or _70872_ (_19101_, _19100_, _06031_);
  and _70873_ (_19102_, _19101_, _18956_);
  or _70874_ (_19103_, _19102_, _06277_);
  and _70875_ (_19104_, _08954_, _08017_);
  or _70876_ (_19105_, _19104_, _18946_);
  or _70877_ (_19106_, _19105_, _06278_);
  and _70878_ (_19107_, _19106_, _11029_);
  and _70879_ (_19108_, _19107_, _19103_);
  nor _70880_ (_19109_, _11029_, _06685_);
  or _70881_ (_19110_, _19109_, _18318_);
  or _70882_ (_19111_, _19110_, _19108_);
  or _70883_ (_19112_, _11257_, _18319_);
  and _70884_ (_19113_, _19112_, _06965_);
  and _70885_ (_19114_, _19113_, _19111_);
  or _70886_ (_19115_, _19114_, _18955_);
  and _70887_ (_19116_, _19115_, _18954_);
  and _70888_ (_19117_, _11257_, _06803_);
  or _70889_ (_19118_, _19117_, _06802_);
  or _70890_ (_19119_, _19118_, _19116_);
  or _70891_ (_19120_, _11257_, _11044_);
  and _70892_ (_19121_, _19120_, _18951_);
  and _70893_ (_19122_, _19121_, _19119_);
  or _70894_ (_19123_, _19122_, _18953_);
  and _70895_ (_19124_, _19123_, _11060_);
  nor _70896_ (_19125_, _11060_, _11299_);
  or _70897_ (_19126_, _19125_, _06613_);
  or _70898_ (_19127_, _19126_, _19124_);
  and _70899_ (_19128_, _19127_, _18950_);
  and _70900_ (_19129_, _11064_, _12644_);
  or _70901_ (_19130_, _19129_, _06502_);
  or _70902_ (_19131_, _19130_, _19128_);
  and _70903_ (_19132_, _19131_, _18948_);
  or _70904_ (_19133_, _19132_, _06615_);
  or _70905_ (_19134_, _18946_, _07337_);
  and _70906_ (_19135_, _19134_, _10616_);
  and _70907_ (_19136_, _19135_, _19133_);
  or _70908_ (_19137_, _19136_, _18944_);
  and _70909_ (_19138_, _19137_, _06973_);
  and _70910_ (_19139_, _11255_, _06972_);
  or _70911_ (_19140_, _19139_, _19138_);
  and _70912_ (_19141_, _19140_, _10611_);
  and _70913_ (_19142_, _11297_, _06976_);
  or _70914_ (_19143_, _19142_, _06608_);
  or _70915_ (_19144_, _19143_, _19141_);
  or _70916_ (_19145_, _10569_, _06609_);
  and _70917_ (_19146_, _19145_, _11090_);
  and _70918_ (_19147_, _19146_, _19144_);
  and _70919_ (_19148_, _11089_, _11339_);
  or _70920_ (_19149_, _19148_, _19147_);
  and _70921_ (_19150_, _19149_, _07339_);
  nand _70922_ (_19151_, _19105_, _06507_);
  nor _70923_ (_19152_, _19151_, _10570_);
  or _70924_ (_19153_, _19152_, _19150_);
  and _70925_ (_19154_, _19153_, _17452_);
  nor _70926_ (_19155_, _11256_, _17452_);
  or _70927_ (_19156_, _19155_, _11102_);
  or _70928_ (_19157_, _19156_, _19154_);
  and _70929_ (_19158_, _19157_, _18943_);
  nor _70930_ (_19159_, _11256_, _06985_);
  or _70931_ (_19160_, _19159_, _06987_);
  or _70932_ (_19161_, _19160_, _19158_);
  nand _70933_ (_19162_, _06987_, _10237_);
  or _70934_ (_19163_, _19162_, _09218_);
  and _70935_ (_19164_, _19163_, _06605_);
  and _70936_ (_19165_, _19164_, _19161_);
  nor _70937_ (_19166_, _10570_, _06605_);
  or _70938_ (_19167_, _19166_, _11114_);
  or _70939_ (_19168_, _19167_, _19165_);
  nand _70940_ (_19169_, _11114_, _11340_);
  and _70941_ (_19170_, _19169_, _09107_);
  and _70942_ (_19171_, _19170_, _19168_);
  and _70943_ (_19172_, _15663_, _08017_);
  or _70944_ (_19173_, _19172_, _18946_);
  and _70945_ (_19174_, _19173_, _06509_);
  or _70946_ (_19175_, _19174_, _11130_);
  or _70947_ (_19176_, _19175_, _19171_);
  and _70948_ (_19177_, _19176_, _18941_);
  or _70949_ (_19178_, _19177_, _11129_);
  and _70950_ (_19179_, _11175_, _10874_);
  nor _70951_ (_19180_, _19179_, _11176_);
  or _70952_ (_19181_, _19180_, _11158_);
  and _70953_ (_19182_, _19181_, _06601_);
  and _70954_ (_19183_, _19182_, _19178_);
  nand _70955_ (_19184_, _11205_, _10648_);
  nor _70956_ (_19185_, _11206_, _06601_);
  and _70957_ (_19186_, _19185_, _19184_);
  or _70958_ (_19187_, _19186_, _11186_);
  or _70959_ (_19188_, _19187_, _19183_);
  and _70960_ (_19189_, _11234_, _10950_);
  nor _70961_ (_19190_, _19189_, _11235_);
  or _70962_ (_19191_, _19190_, _11218_);
  and _70963_ (_19192_, _19191_, _11217_);
  and _70964_ (_19193_, _19192_, _19188_);
  and _70965_ (_19194_, _07577_, _06360_);
  and _70966_ (_19195_, _11216_, \oc8051_golden_model_1.ACC [4]);
  or _70967_ (_19196_, _19195_, _19194_);
  or _70968_ (_19197_, _19196_, _19193_);
  and _70969_ (_19198_, _06315_, _06360_);
  not _70970_ (_19199_, _19194_);
  nor _70971_ (_19200_, _11280_, _11257_);
  nor _70972_ (_19201_, _19200_, _11281_);
  nor _70973_ (_19202_, _19201_, _19199_);
  nor _70974_ (_19203_, _19202_, _19198_);
  and _70975_ (_19204_, _19203_, _19197_);
  and _70976_ (_19205_, _19201_, _19198_);
  or _70977_ (_19206_, _19205_, _11290_);
  or _70978_ (_19207_, _19206_, _19204_);
  and _70979_ (_19208_, _11322_, _11299_);
  nor _70980_ (_19209_, _19208_, _11323_);
  or _70981_ (_19210_, _19209_, _11292_);
  and _70982_ (_19211_, _19210_, _06364_);
  and _70983_ (_19212_, _19211_, _19207_);
  and _70984_ (_19213_, _12626_, _10592_);
  nor _70985_ (_19214_, _12626_, _10592_);
  or _70986_ (_19215_, _19214_, _19213_);
  and _70987_ (_19216_, _19215_, _06363_);
  or _70988_ (_19217_, _19216_, _10566_);
  or _70989_ (_19218_, _19217_, _19212_);
  and _70990_ (_19219_, _11364_, _12644_);
  nor _70991_ (_19220_, _11364_, _12644_);
  or _70992_ (_19221_, _19220_, _19219_);
  or _70993_ (_19222_, _19221_, _10567_);
  and _70994_ (_19223_, _19222_, _13049_);
  and _70995_ (_19224_, _19223_, _19218_);
  and _70996_ (_19225_, _10564_, \oc8051_golden_model_1.ACC [4]);
  or _70997_ (_19226_, _19225_, _06639_);
  or _70998_ (_19227_, _19226_, _19224_);
  or _70999_ (_19228_, _18985_, _07048_);
  and _71000_ (_19229_, _19228_, _11378_);
  and _71001_ (_19230_, _19229_, _19227_);
  nor _71002_ (_19231_, _11385_, _10237_);
  or _71003_ (_19232_, _19231_, _11386_);
  and _71004_ (_19233_, _19232_, _11377_);
  or _71005_ (_19234_, _19233_, _11382_);
  or _71006_ (_19235_, _19234_, _19230_);
  nand _71007_ (_19236_, _11382_, _10193_);
  and _71008_ (_19237_, _19236_, _05990_);
  and _71009_ (_19238_, _19237_, _19235_);
  and _71010_ (_19239_, _19015_, _05989_);
  or _71011_ (_19240_, _19239_, _06646_);
  or _71012_ (_19241_, _19240_, _19238_);
  and _71013_ (_19242_, _15721_, _08017_);
  or _71014_ (_19243_, _18946_, _06651_);
  or _71015_ (_19244_, _19243_, _19242_);
  and _71016_ (_19245_, _19244_, _11401_);
  and _71017_ (_19246_, _19245_, _19241_);
  nor _71018_ (_19247_, _11411_, \oc8051_golden_model_1.ACC [5]);
  nor _71019_ (_19248_, _19247_, _11412_);
  and _71020_ (_19249_, _19248_, _11400_);
  or _71021_ (_19250_, _19249_, _11407_);
  or _71022_ (_19251_, _19250_, _19246_);
  nand _71023_ (_19252_, _11407_, _10193_);
  and _71024_ (_19253_, _19252_, _01442_);
  and _71025_ (_19254_, _19253_, _19251_);
  or _71026_ (_19255_, _19254_, _18938_);
  and _71027_ (_44129_, _19255_, _43634_);
  nor _71028_ (_19256_, _01442_, _10193_);
  or _71029_ (_19257_, _11236_, _10991_);
  and _71030_ (_19258_, _19257_, _11237_);
  or _71031_ (_19259_, _19258_, _11218_);
  nand _71032_ (_19260_, _11114_, _11337_);
  and _71033_ (_19261_, _15862_, _08017_);
  nor _71034_ (_19262_, _08017_, _10193_);
  or _71035_ (_19263_, _19262_, _07334_);
  or _71036_ (_19264_, _19263_, _19261_);
  or _71037_ (_19265_, _10596_, _06614_);
  and _71038_ (_19266_, _19265_, _11071_);
  and _71039_ (_19267_, _15846_, _08017_);
  or _71040_ (_19268_, _19267_, _19262_);
  and _71041_ (_19269_, _19268_, _06037_);
  nor _71042_ (_19270_, _08209_, _10619_);
  or _71043_ (_19271_, _19270_, _19262_);
  or _71044_ (_19272_, _19271_, _06327_);
  or _71045_ (_19273_, _09218_, _10237_);
  and _71046_ (_19274_, _09218_, _10237_);
  or _71047_ (_19275_, _19046_, _19274_);
  and _71048_ (_19276_, _19275_, _19273_);
  nor _71049_ (_19277_, _19276_, _11296_);
  and _71050_ (_19278_, _19276_, _11296_);
  nor _71051_ (_19279_, _19278_, _19277_);
  not _71052_ (_19280_, _19279_);
  or _71053_ (_19281_, _19055_, _19050_);
  or _71054_ (_19282_, _19281_, _10967_);
  nand _71055_ (_19283_, _19282_, _19280_);
  or _71056_ (_19284_, _19282_, _19280_);
  and _71057_ (_19285_, _19284_, _19283_);
  or _71058_ (_19286_, _19285_, _10854_);
  nand _71059_ (_19287_, _10696_, _08209_);
  and _71060_ (_19288_, _10703_, _09172_);
  nor _71061_ (_19289_, _06855_, _10193_);
  and _71062_ (_19290_, _06855_, _10193_);
  or _71063_ (_19291_, _19290_, _19289_);
  and _71064_ (_19292_, _19291_, _10714_);
  nor _71065_ (_19293_, _10712_, _08209_);
  or _71066_ (_19294_, _19293_, _19292_);
  or _71067_ (_19295_, _19294_, _19288_);
  and _71068_ (_19296_, _19295_, _10722_);
  and _71069_ (_19297_, _15759_, _08017_);
  or _71070_ (_19298_, _19297_, _19262_);
  and _71071_ (_19299_, _19298_, _06474_);
  or _71072_ (_19300_, _19299_, _10729_);
  or _71073_ (_19301_, _19300_, _19296_);
  or _71074_ (_19302_, _18989_, _10744_);
  nand _71075_ (_19303_, _18989_, _10744_);
  and _71076_ (_19304_, _19303_, _19302_);
  or _71077_ (_19305_, _19304_, _10730_);
  and _71078_ (_19306_, _19305_, _06418_);
  and _71079_ (_19307_, _19306_, _19301_);
  nor _71080_ (_19308_, _08645_, _10193_);
  and _71081_ (_19309_, _15763_, _08645_);
  or _71082_ (_19310_, _19309_, _19308_);
  and _71083_ (_19311_, _19310_, _06356_);
  and _71084_ (_19312_, _19271_, _06410_);
  or _71085_ (_19313_, _19312_, _10696_);
  or _71086_ (_19314_, _19313_, _19311_);
  or _71087_ (_19315_, _19314_, _19307_);
  and _71088_ (_19316_, _19315_, _19287_);
  or _71089_ (_19317_, _19316_, _07289_);
  or _71090_ (_19318_, _09172_, _07290_);
  and _71091_ (_19319_, _19318_, _06426_);
  and _71092_ (_19320_, _19319_, _19317_);
  nor _71093_ (_19321_, _08211_, _06426_);
  or _71094_ (_19322_, _19321_, _10694_);
  or _71095_ (_19323_, _19322_, _19320_);
  nand _71096_ (_19324_, _10694_, _10280_);
  and _71097_ (_19325_, _19324_, _19323_);
  or _71098_ (_19326_, _19325_, _06352_);
  and _71099_ (_19327_, _15743_, _08645_);
  or _71100_ (_19328_, _19327_, _19308_);
  or _71101_ (_19329_, _19328_, _06353_);
  and _71102_ (_19330_, _19329_, _06346_);
  and _71103_ (_19331_, _19330_, _19326_);
  or _71104_ (_19332_, _19308_, _15778_);
  and _71105_ (_19333_, _19310_, _06345_);
  and _71106_ (_19334_, _19333_, _19332_);
  or _71107_ (_19335_, _19334_, _09606_);
  or _71108_ (_19336_, _19335_, _19331_);
  nor _71109_ (_19337_, _10109_, _10107_);
  nor _71110_ (_19338_, _19337_, _10110_);
  or _71111_ (_19339_, _19338_, _09612_);
  and _71112_ (_19340_, _19339_, _10784_);
  and _71113_ (_19341_, _19340_, _19336_);
  nand _71114_ (_19342_, _08305_, \oc8051_golden_model_1.ACC [5]);
  nor _71115_ (_19343_, _08305_, \oc8051_golden_model_1.ACC [5]);
  or _71116_ (_19344_, _19030_, _19343_);
  and _71117_ (_19345_, _19344_, _19342_);
  nor _71118_ (_19346_, _19345_, _11254_);
  and _71119_ (_19347_, _19345_, _11254_);
  nor _71120_ (_19348_, _19347_, _19346_);
  nor _71121_ (_19349_, _19039_, _19034_);
  and _71122_ (_19350_, _19349_, \oc8051_golden_model_1.PSW [7]);
  nand _71123_ (_19351_, _19350_, _19348_);
  or _71124_ (_19352_, _19350_, _19348_);
  and _71125_ (_19353_, _19352_, _12338_);
  and _71126_ (_19354_, _19353_, _19351_);
  or _71127_ (_19355_, _19354_, _10853_);
  or _71128_ (_19356_, _19355_, _19341_);
  and _71129_ (_19357_, _19356_, _12336_);
  and _71130_ (_19358_, _19357_, _19286_);
  or _71131_ (_19359_, _19062_, _14333_);
  and _71132_ (_19360_, _19359_, _14331_);
  nor _71133_ (_19361_, _19360_, _10596_);
  and _71134_ (_19362_, _19360_, _10596_);
  nor _71135_ (_19363_, _19362_, _19361_);
  nor _71136_ (_19364_, _19071_, _19066_);
  and _71137_ (_19365_, _19364_, \oc8051_golden_model_1.PSW [7]);
  or _71138_ (_19366_, _19365_, _19363_);
  nand _71139_ (_19367_, _19365_, _19363_);
  and _71140_ (_19368_, _19367_, _06453_);
  and _71141_ (_19369_, _19368_, _19366_);
  or _71142_ (_19370_, _18961_, _14352_);
  and _71143_ (_19371_, _19370_, _14351_);
  nor _71144_ (_19372_, _19371_, _11338_);
  and _71145_ (_19373_, _19371_, _11338_);
  nor _71146_ (_19374_, _19373_, _19372_);
  nor _71147_ (_19375_, _18970_, _18965_);
  and _71148_ (_19376_, _19375_, \oc8051_golden_model_1.PSW [7]);
  or _71149_ (_19377_, _19376_, _19374_);
  nand _71150_ (_19378_, _19376_, _19374_);
  and _71151_ (_19379_, _19378_, _10623_);
  and _71152_ (_19380_, _19379_, _19377_);
  or _71153_ (_19381_, _19380_, _06042_);
  or _71154_ (_19382_, _19381_, _19369_);
  or _71155_ (_19383_, _19382_, _19358_);
  nand _71156_ (_19384_, _06397_, _06042_);
  and _71157_ (_19385_, _19384_, _06340_);
  and _71158_ (_19386_, _19385_, _19383_);
  and _71159_ (_19387_, _15745_, _08645_);
  or _71160_ (_19388_, _19387_, _19308_);
  and _71161_ (_19389_, _19388_, _06339_);
  or _71162_ (_19390_, _19389_, _10153_);
  or _71163_ (_19391_, _19390_, _19386_);
  and _71164_ (_19392_, _19391_, _19272_);
  or _71165_ (_19393_, _19392_, _09572_);
  and _71166_ (_19394_, _09172_, _08017_);
  or _71167_ (_19395_, _19262_, _06333_);
  or _71168_ (_19396_, _19395_, _19394_);
  and _71169_ (_19397_, _19396_, _06313_);
  and _71170_ (_19398_, _19397_, _19393_);
  or _71171_ (_19399_, _19398_, _19269_);
  and _71172_ (_19400_, _19399_, _12694_);
  nor _71173_ (_19401_, _06397_, _06032_);
  nand _71174_ (_19402_, _10189_, _10185_);
  nor _71175_ (_19403_, _19402_, _06030_);
  and _71176_ (_19404_, _19403_, _10166_);
  or _71177_ (_19405_, _19404_, _19401_);
  or _71178_ (_19406_, _19405_, _19400_);
  and _71179_ (_19407_, _19406_, _06278_);
  and _71180_ (_19408_, _15853_, _08017_);
  or _71181_ (_19409_, _19408_, _19262_);
  and _71182_ (_19410_, _19409_, _06277_);
  or _71183_ (_19411_, _19410_, _11028_);
  or _71184_ (_19412_, _19411_, _19407_);
  nand _71185_ (_19413_, _11028_, _06397_);
  and _71186_ (_19414_, _19413_, _18319_);
  and _71187_ (_19415_, _19414_, _19412_);
  and _71188_ (_19416_, _11254_, _18318_);
  or _71189_ (_19417_, _19416_, _19415_);
  or _71190_ (_19418_, _19417_, _06964_);
  or _71191_ (_19419_, _11254_, _06965_);
  or _71192_ (_19420_, _17573_, _11045_);
  nand _71193_ (_19421_, _18645_, _18954_);
  nor _71194_ (_19422_, _19421_, _19420_);
  and _71195_ (_19423_, _19422_, _19419_);
  and _71196_ (_19424_, _19423_, _19418_);
  not _71197_ (_19425_, _19422_);
  and _71198_ (_19426_, _19425_, _11254_);
  or _71199_ (_19427_, _19426_, _06966_);
  or _71200_ (_19428_, _19427_, _19424_);
  or _71201_ (_19429_, _11254_, _17570_);
  and _71202_ (_19430_, _19429_, _11060_);
  and _71203_ (_19431_, _19430_, _19428_);
  and _71204_ (_19432_, _11052_, _11296_);
  or _71205_ (_19433_, _19432_, _06613_);
  or _71206_ (_19434_, _19433_, _19431_);
  and _71207_ (_19435_, _19434_, _19266_);
  and _71208_ (_19436_, _11064_, _11338_);
  or _71209_ (_19437_, _19436_, _06502_);
  or _71210_ (_19438_, _19437_, _19435_);
  and _71211_ (_19439_, _19438_, _19264_);
  or _71212_ (_19440_, _19439_, _06615_);
  or _71213_ (_19441_, _19262_, _07337_);
  and _71214_ (_19442_, _19441_, _17595_);
  and _71215_ (_19443_, _19442_, _19440_);
  and _71216_ (_19444_, _17598_, _11251_);
  or _71217_ (_19445_, _19444_, _06976_);
  or _71218_ (_19446_, _19445_, _19443_);
  or _71219_ (_19447_, _11293_, _10611_);
  and _71220_ (_19449_, _19447_, _06609_);
  and _71221_ (_19450_, _19449_, _19446_);
  and _71222_ (_19451_, _10568_, _06608_);
  or _71223_ (_19452_, _19451_, _11089_);
  or _71224_ (_19453_, _19452_, _19450_);
  or _71225_ (_19454_, _11090_, _11335_);
  and _71226_ (_19455_, _19454_, _07339_);
  and _71227_ (_19456_, _19455_, _19453_);
  nand _71228_ (_19457_, _19409_, _06507_);
  nor _71229_ (_19458_, _19457_, _10595_);
  or _71230_ (_19460_, _19458_, _19456_);
  and _71231_ (_19461_, _19460_, _17452_);
  and _71232_ (_19462_, _11253_, _10609_);
  or _71233_ (_19463_, _19462_, _11102_);
  or _71234_ (_19464_, _19463_, _19461_);
  and _71235_ (_19465_, _11253_, _06985_);
  or _71236_ (_19466_, _19465_, _11104_);
  and _71237_ (_19467_, _19466_, _19464_);
  and _71238_ (_19468_, _11253_, _06984_);
  or _71239_ (_19469_, _19468_, _06987_);
  or _71240_ (_19471_, _19469_, _19467_);
  or _71241_ (_19472_, _11294_, _18853_);
  and _71242_ (_19473_, _19472_, _06605_);
  and _71243_ (_19474_, _19473_, _19471_);
  nand _71244_ (_19475_, _17625_, _10595_);
  and _71245_ (_19476_, _19475_, _12315_);
  or _71246_ (_19477_, _19476_, _19474_);
  and _71247_ (_19478_, _19477_, _19260_);
  or _71248_ (_19479_, _19478_, _06509_);
  and _71249_ (_19480_, _15859_, _08017_);
  or _71250_ (_19482_, _19262_, _09107_);
  or _71251_ (_19483_, _19482_, _19480_);
  and _71252_ (_19484_, _19483_, _11127_);
  and _71253_ (_19485_, _19484_, _19479_);
  nor _71254_ (_19486_, _11149_, _10846_);
  nor _71255_ (_19487_, _19486_, _11150_);
  and _71256_ (_19488_, _19487_, _11130_);
  or _71257_ (_19489_, _19488_, _17922_);
  or _71258_ (_19490_, _19489_, _19485_);
  or _71259_ (_19491_, _11177_, _10917_);
  and _71260_ (_19493_, _19491_, _11178_);
  or _71261_ (_19494_, _19493_, _18231_);
  and _71262_ (_19495_, _19494_, _19490_);
  or _71263_ (_19496_, _19495_, _07002_);
  or _71264_ (_19497_, _19493_, _18237_);
  and _71265_ (_19498_, _19497_, _06601_);
  and _71266_ (_19499_, _19498_, _19496_);
  or _71267_ (_19500_, _11207_, _10685_);
  and _71268_ (_19501_, _11208_, _06600_);
  and _71269_ (_19502_, _19501_, _19500_);
  or _71270_ (_19504_, _19502_, _11186_);
  or _71271_ (_19505_, _19504_, _19499_);
  and _71272_ (_19506_, _19505_, _19259_);
  or _71273_ (_19507_, _19506_, _11216_);
  nand _71274_ (_19508_, _11216_, _10237_);
  and _71275_ (_19509_, _19508_, _11248_);
  and _71276_ (_19510_, _19509_, _19507_);
  nor _71277_ (_19511_, _11282_, _11254_);
  nor _71278_ (_19512_, _19511_, _11283_);
  and _71279_ (_19513_, _19512_, _18254_);
  or _71280_ (_19515_, _19513_, _17690_);
  or _71281_ (_19516_, _19515_, _19510_);
  nor _71282_ (_19517_, _11324_, _11296_);
  nor _71283_ (_19518_, _19517_, _11325_);
  or _71284_ (_19519_, _19518_, _17691_);
  and _71285_ (_19520_, _19519_, _19516_);
  or _71286_ (_19521_, _19520_, _07019_);
  or _71287_ (_19522_, _19518_, _07020_);
  and _71288_ (_19523_, _19522_, _06364_);
  and _71289_ (_19524_, _19523_, _19521_);
  nor _71290_ (_19526_, _10596_, _10594_);
  nor _71291_ (_19527_, _19526_, _10597_);
  or _71292_ (_19528_, _19527_, _10566_);
  and _71293_ (_19529_, _19528_, _13047_);
  or _71294_ (_19530_, _19529_, _19524_);
  or _71295_ (_19531_, _11366_, _11338_);
  and _71296_ (_19532_, _19531_, _11367_);
  or _71297_ (_19533_, _19532_, _10567_);
  and _71298_ (_19534_, _19533_, _13049_);
  and _71299_ (_19535_, _19534_, _19530_);
  and _71300_ (_19537_, _10564_, \oc8051_golden_model_1.ACC [5]);
  or _71301_ (_19538_, _19537_, _06639_);
  or _71302_ (_19539_, _19538_, _19535_);
  or _71303_ (_19540_, _19298_, _07048_);
  and _71304_ (_19541_, _19540_, _11378_);
  and _71305_ (_19542_, _19541_, _19539_);
  nor _71306_ (_19543_, _11386_, _10193_);
  or _71307_ (_19544_, _19543_, _11387_);
  and _71308_ (_19545_, _19544_, _11377_);
  or _71309_ (_19546_, _19545_, _11382_);
  or _71310_ (_19548_, _19546_, _19542_);
  nand _71311_ (_19549_, _11382_, _08688_);
  and _71312_ (_19550_, _19549_, _05990_);
  and _71313_ (_19551_, _19550_, _19548_);
  and _71314_ (_19552_, _19328_, _05989_);
  or _71315_ (_19553_, _19552_, _06646_);
  or _71316_ (_19554_, _19553_, _19551_);
  and _71317_ (_19555_, _15921_, _08017_);
  or _71318_ (_19556_, _19262_, _06651_);
  or _71319_ (_19557_, _19556_, _19555_);
  and _71320_ (_19559_, _19557_, _11401_);
  and _71321_ (_19560_, _19559_, _19554_);
  nor _71322_ (_19561_, _11412_, \oc8051_golden_model_1.ACC [6]);
  nor _71323_ (_19562_, _19561_, _11413_);
  and _71324_ (_19563_, _19562_, _11400_);
  or _71325_ (_19564_, _19563_, _11407_);
  or _71326_ (_19565_, _19564_, _19560_);
  nand _71327_ (_19566_, _11407_, _08688_);
  and _71328_ (_19567_, _19566_, _01442_);
  and _71329_ (_19568_, _19567_, _19565_);
  or _71330_ (_19570_, _19568_, _19256_);
  and _71331_ (_44130_, _19570_, _43634_);
  not _71332_ (_19571_, \oc8051_golden_model_1.PCON [0]);
  nor _71333_ (_19572_, _01442_, _19571_);
  nor _71334_ (_19573_, _08042_, _19571_);
  nor _71335_ (_19574_, _12622_, _11424_);
  or _71336_ (_19575_, _19574_, _19573_);
  and _71337_ (_19576_, _10577_, _08042_);
  nor _71338_ (_19577_, _19576_, _07337_);
  and _71339_ (_19578_, _19577_, _19575_);
  and _71340_ (_19580_, _08042_, \oc8051_golden_model_1.ACC [0]);
  or _71341_ (_19581_, _19580_, _19573_);
  and _71342_ (_19582_, _19581_, _06417_);
  or _71343_ (_19583_, _19582_, _10153_);
  nor _71344_ (_19584_, _08453_, _11424_);
  or _71345_ (_19585_, _19584_, _19573_);
  and _71346_ (_19586_, _19585_, _06474_);
  nor _71347_ (_19587_, _07259_, _19571_);
  and _71348_ (_19588_, _19581_, _07259_);
  or _71349_ (_19589_, _19588_, _19587_);
  and _71350_ (_19591_, _19589_, _07275_);
  or _71351_ (_19592_, _19591_, _06410_);
  or _71352_ (_19593_, _19592_, _19586_);
  and _71353_ (_19594_, _19593_, _06426_);
  or _71354_ (_19595_, _19594_, _19583_);
  and _71355_ (_19596_, _08042_, _07250_);
  and _71356_ (_19597_, _06327_, _06772_);
  or _71357_ (_19598_, _19597_, _19573_);
  or _71358_ (_19599_, _19598_, _19596_);
  and _71359_ (_19600_, _19599_, _19595_);
  or _71360_ (_19602_, _19600_, _09572_);
  and _71361_ (_19603_, _09447_, _08042_);
  or _71362_ (_19604_, _19573_, _06333_);
  or _71363_ (_19605_, _19604_, _19603_);
  and _71364_ (_19606_, _19605_, _19602_);
  or _71365_ (_19607_, _19606_, _06037_);
  and _71366_ (_19608_, _14666_, _08042_);
  or _71367_ (_19609_, _19573_, _06313_);
  or _71368_ (_19610_, _19609_, _19608_);
  and _71369_ (_19611_, _19610_, _06278_);
  and _71370_ (_19613_, _19611_, _19607_);
  and _71371_ (_19614_, _08042_, _09008_);
  or _71372_ (_19615_, _19614_, _19573_);
  and _71373_ (_19616_, _19615_, _06277_);
  or _71374_ (_19617_, _19616_, _06502_);
  or _71375_ (_19618_, _19617_, _19613_);
  and _71376_ (_19619_, _14566_, _08042_);
  or _71377_ (_19620_, _19573_, _07334_);
  or _71378_ (_19621_, _19620_, _19619_);
  and _71379_ (_19622_, _19621_, _07337_);
  and _71380_ (_19623_, _19622_, _19618_);
  or _71381_ (_19624_, _19623_, _19578_);
  and _71382_ (_19625_, _19624_, _07339_);
  nand _71383_ (_19626_, _19615_, _06507_);
  nor _71384_ (_19627_, _19626_, _19584_);
  or _71385_ (_19628_, _19627_, _06610_);
  or _71386_ (_19629_, _19628_, _19625_);
  or _71387_ (_19630_, _19576_, _19573_);
  or _71388_ (_19631_, _19630_, _07331_);
  and _71389_ (_19632_, _19631_, _19629_);
  or _71390_ (_19634_, _19632_, _06509_);
  and _71391_ (_19635_, _14563_, _08042_);
  or _71392_ (_19636_, _19573_, _09107_);
  or _71393_ (_19637_, _19636_, _19635_);
  and _71394_ (_19638_, _19637_, _09112_);
  and _71395_ (_19639_, _19638_, _19634_);
  and _71396_ (_19640_, _19575_, _06602_);
  nor _71397_ (_19641_, _06646_, _06639_);
  not _71398_ (_19642_, _19641_);
  or _71399_ (_19643_, _19642_, _19640_);
  or _71400_ (_19645_, _19643_, _19639_);
  or _71401_ (_19646_, _19641_, _19585_);
  and _71402_ (_19647_, _19646_, _01442_);
  and _71403_ (_19648_, _19647_, _19645_);
  or _71404_ (_19649_, _19648_, _19572_);
  and _71405_ (_44132_, _19649_, _43634_);
  not _71406_ (_19650_, \oc8051_golden_model_1.PCON [1]);
  nor _71407_ (_19651_, _01442_, _19650_);
  or _71408_ (_19652_, _08042_, \oc8051_golden_model_1.PCON [1]);
  and _71409_ (_19653_, _14744_, _08042_);
  not _71410_ (_19655_, _19653_);
  and _71411_ (_19656_, _19655_, _19652_);
  or _71412_ (_19657_, _19656_, _07275_);
  nor _71413_ (_19658_, _08042_, _19650_);
  and _71414_ (_19659_, _08042_, \oc8051_golden_model_1.ACC [1]);
  or _71415_ (_19660_, _19659_, _19658_);
  and _71416_ (_19661_, _19660_, _07259_);
  nor _71417_ (_19662_, _07259_, _19650_);
  or _71418_ (_19663_, _19662_, _06474_);
  or _71419_ (_19664_, _19663_, _19661_);
  and _71420_ (_19666_, _19664_, _06772_);
  and _71421_ (_19667_, _19666_, _19657_);
  nor _71422_ (_19668_, _11424_, _07448_);
  or _71423_ (_19669_, _19668_, _19658_);
  and _71424_ (_19670_, _19669_, _06410_);
  or _71425_ (_19671_, _19670_, _19667_);
  and _71426_ (_19672_, _19671_, _06426_);
  and _71427_ (_19673_, _19660_, _06417_);
  or _71428_ (_19674_, _19673_, _10153_);
  or _71429_ (_19675_, _19674_, _19672_);
  or _71430_ (_19677_, _19669_, _06327_);
  and _71431_ (_19678_, _19677_, _16672_);
  and _71432_ (_19679_, _19678_, _19675_);
  or _71433_ (_19680_, _09402_, _11424_);
  and _71434_ (_19681_, _19652_, _14025_);
  and _71435_ (_19682_, _19681_, _19680_);
  or _71436_ (_19683_, _19682_, _19679_);
  and _71437_ (_19684_, _19683_, _06313_);
  or _71438_ (_19685_, _14851_, _11424_);
  and _71439_ (_19686_, _19652_, _06037_);
  and _71440_ (_19688_, _19686_, _19685_);
  or _71441_ (_19689_, _19688_, _19684_);
  and _71442_ (_19690_, _19689_, _06278_);
  nand _71443_ (_19691_, _08042_, _07160_);
  and _71444_ (_19692_, _19652_, _06277_);
  and _71445_ (_19693_, _19692_, _19691_);
  or _71446_ (_19694_, _19693_, _19690_);
  and _71447_ (_19695_, _19694_, _07334_);
  or _71448_ (_19696_, _14749_, _11424_);
  and _71449_ (_19697_, _19652_, _06502_);
  and _71450_ (_19699_, _19697_, _19696_);
  or _71451_ (_19700_, _19699_, _06615_);
  or _71452_ (_19701_, _19700_, _19695_);
  and _71453_ (_19702_, _10579_, _08042_);
  or _71454_ (_19703_, _19702_, _19658_);
  or _71455_ (_19704_, _19703_, _07337_);
  and _71456_ (_19705_, _19704_, _07339_);
  and _71457_ (_19706_, _19705_, _19701_);
  or _71458_ (_19707_, _14747_, _11424_);
  and _71459_ (_19708_, _19652_, _06507_);
  and _71460_ (_19710_, _19708_, _19707_);
  or _71461_ (_19711_, _19710_, _06610_);
  or _71462_ (_19712_, _19711_, _19706_);
  and _71463_ (_19713_, _19659_, _08404_);
  or _71464_ (_19714_, _19658_, _07331_);
  or _71465_ (_19715_, _19714_, _19713_);
  and _71466_ (_19716_, _19715_, _09107_);
  and _71467_ (_19717_, _19716_, _19712_);
  or _71468_ (_19718_, _19691_, _08404_);
  and _71469_ (_19719_, _19652_, _06509_);
  and _71470_ (_19722_, _19719_, _19718_);
  or _71471_ (_19723_, _19722_, _06602_);
  or _71472_ (_19724_, _19723_, _19717_);
  nor _71473_ (_19725_, _10578_, _11424_);
  or _71474_ (_19726_, _19725_, _19658_);
  or _71475_ (_19727_, _19726_, _09112_);
  and _71476_ (_19728_, _19727_, _07048_);
  and _71477_ (_19729_, _19728_, _19724_);
  and _71478_ (_19730_, _19656_, _06639_);
  or _71479_ (_19731_, _19730_, _06646_);
  or _71480_ (_19734_, _19731_, _19729_);
  or _71481_ (_19735_, _19658_, _06651_);
  or _71482_ (_19736_, _19735_, _19653_);
  and _71483_ (_19737_, _19736_, _01442_);
  and _71484_ (_19738_, _19737_, _19734_);
  or _71485_ (_19739_, _19738_, _19651_);
  and _71486_ (_44133_, _19739_, _43634_);
  not _71487_ (_19740_, \oc8051_golden_model_1.PCON [2]);
  nor _71488_ (_19741_, _01442_, _19740_);
  nor _71489_ (_19742_, _08042_, _19740_);
  or _71490_ (_19745_, _19742_, _08503_);
  and _71491_ (_19746_, _08042_, _09057_);
  or _71492_ (_19747_, _19746_, _19742_);
  and _71493_ (_19748_, _19747_, _06507_);
  and _71494_ (_19749_, _19748_, _19745_);
  nor _71495_ (_19750_, _10582_, _11424_);
  or _71496_ (_19751_, _19750_, _19742_);
  and _71497_ (_19752_, _08042_, \oc8051_golden_model_1.ACC [2]);
  nand _71498_ (_19753_, _19752_, _08503_);
  and _71499_ (_19754_, _19753_, _06615_);
  and _71500_ (_19757_, _19754_, _19751_);
  and _71501_ (_19758_, _09356_, _08042_);
  or _71502_ (_19759_, _19758_, _19742_);
  and _71503_ (_19760_, _19759_, _14025_);
  and _71504_ (_19761_, _14959_, _08042_);
  or _71505_ (_19762_, _19761_, _19742_);
  or _71506_ (_19763_, _19762_, _07275_);
  or _71507_ (_19764_, _19752_, _19742_);
  and _71508_ (_19765_, _19764_, _07259_);
  nor _71509_ (_19766_, _07259_, _19740_);
  or _71510_ (_19769_, _19766_, _06474_);
  or _71511_ (_19770_, _19769_, _19765_);
  and _71512_ (_19771_, _19770_, _06772_);
  and _71513_ (_19772_, _19771_, _19763_);
  nor _71514_ (_19773_, _11424_, _07854_);
  or _71515_ (_19774_, _19773_, _19742_);
  and _71516_ (_19775_, _19774_, _06410_);
  or _71517_ (_19776_, _19775_, _19772_);
  and _71518_ (_19777_, _19776_, _06426_);
  and _71519_ (_19778_, _19764_, _06417_);
  or _71520_ (_19781_, _19778_, _10153_);
  or _71521_ (_19782_, _19781_, _19777_);
  or _71522_ (_19783_, _19774_, _06327_);
  and _71523_ (_19784_, _19783_, _16672_);
  and _71524_ (_19785_, _19784_, _19782_);
  or _71525_ (_19786_, _19785_, _06037_);
  or _71526_ (_19787_, _19786_, _19760_);
  and _71527_ (_19788_, _15056_, _08042_);
  or _71528_ (_19789_, _19742_, _06313_);
  or _71529_ (_19790_, _19789_, _19788_);
  and _71530_ (_19793_, _19790_, _06278_);
  and _71531_ (_19794_, _19793_, _19787_);
  and _71532_ (_19795_, _19747_, _06277_);
  or _71533_ (_19796_, _19795_, _06502_);
  or _71534_ (_19797_, _19796_, _19794_);
  and _71535_ (_19798_, _14948_, _08042_);
  or _71536_ (_19799_, _19742_, _07334_);
  or _71537_ (_19800_, _19799_, _19798_);
  and _71538_ (_19801_, _19800_, _07337_);
  and _71539_ (_19802_, _19801_, _19797_);
  or _71540_ (_19804_, _19802_, _19757_);
  and _71541_ (_19805_, _19804_, _07339_);
  or _71542_ (_19806_, _19805_, _19749_);
  and _71543_ (_19807_, _19806_, _07331_);
  and _71544_ (_19808_, _19764_, _06610_);
  and _71545_ (_19809_, _19808_, _19745_);
  or _71546_ (_19810_, _19809_, _06509_);
  or _71547_ (_19811_, _19810_, _19807_);
  and _71548_ (_19812_, _14945_, _08042_);
  or _71549_ (_19813_, _19742_, _09107_);
  or _71550_ (_19815_, _19813_, _19812_);
  and _71551_ (_19816_, _19815_, _09112_);
  and _71552_ (_19817_, _19816_, _19811_);
  and _71553_ (_19818_, _19751_, _06602_);
  or _71554_ (_19819_, _19818_, _19817_);
  and _71555_ (_19820_, _19819_, _07048_);
  and _71556_ (_19821_, _19762_, _06639_);
  or _71557_ (_19822_, _19821_, _06646_);
  or _71558_ (_19823_, _19822_, _19820_);
  and _71559_ (_19824_, _15129_, _08042_);
  or _71560_ (_19826_, _19742_, _06651_);
  or _71561_ (_19827_, _19826_, _19824_);
  and _71562_ (_19828_, _19827_, _01442_);
  and _71563_ (_19829_, _19828_, _19823_);
  or _71564_ (_19830_, _19829_, _19741_);
  and _71565_ (_44134_, _19830_, _43634_);
  and _71566_ (_19831_, _11424_, \oc8051_golden_model_1.PCON [3]);
  nor _71567_ (_19832_, _10574_, _11424_);
  or _71568_ (_19833_, _19832_, _19831_);
  and _71569_ (_19834_, _08042_, \oc8051_golden_model_1.ACC [3]);
  nand _71570_ (_19836_, _19834_, _08359_);
  and _71571_ (_19837_, _19836_, _06615_);
  and _71572_ (_19838_, _19837_, _19833_);
  and _71573_ (_19839_, _15153_, _08042_);
  or _71574_ (_19840_, _19839_, _19831_);
  or _71575_ (_19841_, _19840_, _07275_);
  or _71576_ (_19842_, _19834_, _19831_);
  and _71577_ (_19843_, _19842_, _07259_);
  and _71578_ (_19844_, _07260_, \oc8051_golden_model_1.PCON [3]);
  or _71579_ (_19845_, _19844_, _06474_);
  or _71580_ (_19847_, _19845_, _19843_);
  and _71581_ (_19848_, _19847_, _06772_);
  and _71582_ (_19849_, _19848_, _19841_);
  nor _71583_ (_19850_, _11424_, _07680_);
  or _71584_ (_19851_, _19850_, _19831_);
  and _71585_ (_19852_, _19851_, _06410_);
  or _71586_ (_19853_, _19852_, _19849_);
  and _71587_ (_19854_, _19853_, _06426_);
  and _71588_ (_19855_, _19842_, _06417_);
  or _71589_ (_19856_, _19855_, _10153_);
  or _71590_ (_19858_, _19856_, _19854_);
  or _71591_ (_19859_, _19851_, _06327_);
  and _71592_ (_19860_, _19859_, _16672_);
  and _71593_ (_19861_, _19860_, _19858_);
  and _71594_ (_19862_, _09310_, _08042_);
  or _71595_ (_19863_, _19862_, _19831_);
  and _71596_ (_19864_, _19863_, _14025_);
  or _71597_ (_19865_, _19864_, _06037_);
  or _71598_ (_19866_, _19865_, _19861_);
  and _71599_ (_19867_, _15251_, _08042_);
  or _71600_ (_19869_, _19831_, _06313_);
  or _71601_ (_19870_, _19869_, _19867_);
  and _71602_ (_19871_, _19870_, _06278_);
  and _71603_ (_19872_, _19871_, _19866_);
  and _71604_ (_19873_, _08042_, _09014_);
  or _71605_ (_19874_, _19873_, _19831_);
  and _71606_ (_19875_, _19874_, _06277_);
  or _71607_ (_19876_, _19875_, _06502_);
  or _71608_ (_19877_, _19876_, _19872_);
  and _71609_ (_19878_, _15266_, _08042_);
  or _71610_ (_19880_, _19831_, _07334_);
  or _71611_ (_19881_, _19880_, _19878_);
  and _71612_ (_19882_, _19881_, _07337_);
  and _71613_ (_19883_, _19882_, _19877_);
  or _71614_ (_19884_, _19883_, _19838_);
  and _71615_ (_19885_, _19884_, _07339_);
  or _71616_ (_19886_, _19831_, _08359_);
  and _71617_ (_19887_, _19874_, _06507_);
  and _71618_ (_19888_, _19887_, _19886_);
  or _71619_ (_19889_, _19888_, _19885_);
  and _71620_ (_19891_, _19889_, _07331_);
  and _71621_ (_19892_, _19842_, _06610_);
  and _71622_ (_19893_, _19892_, _19886_);
  or _71623_ (_19894_, _19893_, _06509_);
  or _71624_ (_19895_, _19894_, _19891_);
  and _71625_ (_19896_, _15263_, _08042_);
  or _71626_ (_19897_, _19831_, _09107_);
  or _71627_ (_19898_, _19897_, _19896_);
  and _71628_ (_19899_, _19898_, _09112_);
  and _71629_ (_19900_, _19899_, _19895_);
  and _71630_ (_19902_, _19833_, _06602_);
  or _71631_ (_19903_, _19902_, _06639_);
  or _71632_ (_19904_, _19903_, _19900_);
  or _71633_ (_19905_, _19840_, _07048_);
  and _71634_ (_19906_, _19905_, _06651_);
  and _71635_ (_19907_, _19906_, _19904_);
  and _71636_ (_19908_, _15321_, _08042_);
  or _71637_ (_19909_, _19908_, _19831_);
  and _71638_ (_19910_, _19909_, _06646_);
  or _71639_ (_19911_, _19910_, _01446_);
  or _71640_ (_19913_, _19911_, _19907_);
  or _71641_ (_19914_, _01442_, \oc8051_golden_model_1.PCON [3]);
  and _71642_ (_19915_, _19914_, _43634_);
  and _71643_ (_44135_, _19915_, _19913_);
  and _71644_ (_19916_, _11424_, \oc8051_golden_model_1.PCON [4]);
  or _71645_ (_19917_, _19916_, _08599_);
  and _71646_ (_19918_, _08995_, _08042_);
  or _71647_ (_19919_, _19918_, _19916_);
  and _71648_ (_19920_, _19919_, _06507_);
  and _71649_ (_19921_, _19920_, _19917_);
  nor _71650_ (_19923_, _10589_, _11424_);
  or _71651_ (_19924_, _19923_, _19916_);
  and _71652_ (_19925_, _08042_, \oc8051_golden_model_1.ACC [4]);
  nand _71653_ (_19926_, _19925_, _08599_);
  and _71654_ (_19927_, _19926_, _06615_);
  and _71655_ (_19928_, _19927_, _19924_);
  nor _71656_ (_19929_, _08596_, _11424_);
  or _71657_ (_19930_, _19929_, _19916_);
  or _71658_ (_19931_, _19930_, _06327_);
  and _71659_ (_19932_, _15367_, _08042_);
  or _71660_ (_19934_, _19932_, _19916_);
  or _71661_ (_19935_, _19934_, _07275_);
  or _71662_ (_19936_, _19925_, _19916_);
  and _71663_ (_19937_, _19936_, _07259_);
  and _71664_ (_19938_, _07260_, \oc8051_golden_model_1.PCON [4]);
  or _71665_ (_19939_, _19938_, _06474_);
  or _71666_ (_19940_, _19939_, _19937_);
  and _71667_ (_19941_, _19940_, _06772_);
  and _71668_ (_19942_, _19941_, _19935_);
  and _71669_ (_19943_, _19930_, _06410_);
  or _71670_ (_19945_, _19943_, _19942_);
  and _71671_ (_19946_, _19945_, _06426_);
  and _71672_ (_19947_, _19936_, _06417_);
  or _71673_ (_19948_, _19947_, _10153_);
  or _71674_ (_19949_, _19948_, _19946_);
  and _71675_ (_19950_, _19949_, _19931_);
  or _71676_ (_19951_, _19950_, _09572_);
  and _71677_ (_19952_, _09264_, _08042_);
  or _71678_ (_19953_, _19916_, _16672_);
  or _71679_ (_19954_, _19953_, _19952_);
  and _71680_ (_19956_, _19954_, _19951_);
  or _71681_ (_19957_, _19956_, _06037_);
  and _71682_ (_19958_, _15452_, _08042_);
  or _71683_ (_19959_, _19916_, _06313_);
  or _71684_ (_19960_, _19959_, _19958_);
  and _71685_ (_19961_, _19960_, _06278_);
  and _71686_ (_19962_, _19961_, _19957_);
  and _71687_ (_19963_, _19919_, _06277_);
  or _71688_ (_19964_, _19963_, _06502_);
  or _71689_ (_19965_, _19964_, _19962_);
  and _71690_ (_19967_, _15345_, _08042_);
  or _71691_ (_19968_, _19916_, _07334_);
  or _71692_ (_19969_, _19968_, _19967_);
  and _71693_ (_19970_, _19969_, _07337_);
  and _71694_ (_19971_, _19970_, _19965_);
  or _71695_ (_19972_, _19971_, _19928_);
  and _71696_ (_19973_, _19972_, _07339_);
  or _71697_ (_19974_, _19973_, _19921_);
  and _71698_ (_19975_, _19974_, _07331_);
  and _71699_ (_19976_, _19936_, _06610_);
  and _71700_ (_19978_, _19976_, _19917_);
  or _71701_ (_19979_, _19978_, _06509_);
  or _71702_ (_19980_, _19979_, _19975_);
  and _71703_ (_19981_, _15342_, _08042_);
  or _71704_ (_19982_, _19916_, _09107_);
  or _71705_ (_19983_, _19982_, _19981_);
  and _71706_ (_19984_, _19983_, _09112_);
  and _71707_ (_19985_, _19984_, _19980_);
  and _71708_ (_19986_, _19924_, _06602_);
  or _71709_ (_19987_, _19986_, _06639_);
  or _71710_ (_19989_, _19987_, _19985_);
  or _71711_ (_19990_, _19934_, _07048_);
  and _71712_ (_19991_, _19990_, _06651_);
  and _71713_ (_19992_, _19991_, _19989_);
  and _71714_ (_19993_, _15524_, _08042_);
  or _71715_ (_19994_, _19993_, _19916_);
  and _71716_ (_19995_, _19994_, _06646_);
  or _71717_ (_19996_, _19995_, _01446_);
  or _71718_ (_19997_, _19996_, _19992_);
  or _71719_ (_19998_, _01442_, \oc8051_golden_model_1.PCON [4]);
  and _71720_ (_20000_, _19998_, _43634_);
  and _71721_ (_44136_, _20000_, _19997_);
  and _71722_ (_20001_, _11424_, \oc8051_golden_model_1.PCON [5]);
  nor _71723_ (_20002_, _08305_, _11424_);
  or _71724_ (_20003_, _20002_, _20001_);
  or _71725_ (_20004_, _20003_, _06327_);
  and _71726_ (_20005_, _15550_, _08042_);
  or _71727_ (_20006_, _20005_, _20001_);
  or _71728_ (_20007_, _20006_, _07275_);
  and _71729_ (_20008_, _08042_, \oc8051_golden_model_1.ACC [5]);
  or _71730_ (_20010_, _20008_, _20001_);
  and _71731_ (_20011_, _20010_, _07259_);
  and _71732_ (_20012_, _07260_, \oc8051_golden_model_1.PCON [5]);
  or _71733_ (_20013_, _20012_, _06474_);
  or _71734_ (_20014_, _20013_, _20011_);
  and _71735_ (_20015_, _20014_, _06772_);
  and _71736_ (_20016_, _20015_, _20007_);
  and _71737_ (_20017_, _20003_, _06410_);
  or _71738_ (_20018_, _20017_, _20016_);
  and _71739_ (_20019_, _20018_, _06426_);
  and _71740_ (_20021_, _20010_, _06417_);
  or _71741_ (_20022_, _20021_, _10153_);
  or _71742_ (_20023_, _20022_, _20019_);
  and _71743_ (_20024_, _20023_, _20004_);
  or _71744_ (_20025_, _20024_, _09572_);
  and _71745_ (_20026_, _09218_, _08042_);
  or _71746_ (_20027_, _20001_, _06333_);
  or _71747_ (_20028_, _20027_, _20026_);
  and _71748_ (_20029_, _20028_, _06313_);
  and _71749_ (_20030_, _20029_, _20025_);
  and _71750_ (_20032_, _15649_, _08042_);
  or _71751_ (_20033_, _20032_, _20001_);
  and _71752_ (_20034_, _20033_, _06037_);
  or _71753_ (_20035_, _20034_, _06277_);
  or _71754_ (_20036_, _20035_, _20030_);
  and _71755_ (_20037_, _08954_, _08042_);
  or _71756_ (_20038_, _20037_, _20001_);
  or _71757_ (_20039_, _20038_, _06278_);
  and _71758_ (_20040_, _20039_, _20036_);
  or _71759_ (_20041_, _20040_, _06502_);
  and _71760_ (_20043_, _15664_, _08042_);
  or _71761_ (_20044_, _20001_, _07334_);
  or _71762_ (_20045_, _20044_, _20043_);
  and _71763_ (_20046_, _20045_, _07337_);
  and _71764_ (_20047_, _20046_, _20041_);
  and _71765_ (_20048_, _12626_, _08042_);
  or _71766_ (_20049_, _20048_, _20001_);
  and _71767_ (_20050_, _20049_, _06615_);
  or _71768_ (_20051_, _20050_, _20047_);
  and _71769_ (_20052_, _20051_, _07339_);
  or _71770_ (_20054_, _20001_, _08308_);
  and _71771_ (_20055_, _20038_, _06507_);
  and _71772_ (_20056_, _20055_, _20054_);
  or _71773_ (_20057_, _20056_, _20052_);
  and _71774_ (_20058_, _20057_, _07331_);
  and _71775_ (_20059_, _20010_, _06610_);
  and _71776_ (_20060_, _20059_, _20054_);
  or _71777_ (_20061_, _20060_, _06509_);
  or _71778_ (_20062_, _20061_, _20058_);
  and _71779_ (_20063_, _15663_, _08042_);
  or _71780_ (_20065_, _20001_, _09107_);
  or _71781_ (_20066_, _20065_, _20063_);
  and _71782_ (_20067_, _20066_, _09112_);
  and _71783_ (_20068_, _20067_, _20062_);
  nor _71784_ (_20069_, _10570_, _11424_);
  or _71785_ (_20070_, _20069_, _20001_);
  and _71786_ (_20071_, _20070_, _06602_);
  or _71787_ (_20072_, _20071_, _06639_);
  or _71788_ (_20073_, _20072_, _20068_);
  or _71789_ (_20074_, _20006_, _07048_);
  and _71790_ (_20076_, _20074_, _06651_);
  and _71791_ (_20077_, _20076_, _20073_);
  and _71792_ (_20078_, _15721_, _08042_);
  or _71793_ (_20079_, _20078_, _20001_);
  and _71794_ (_20080_, _20079_, _06646_);
  or _71795_ (_20081_, _20080_, _01446_);
  or _71796_ (_20082_, _20081_, _20077_);
  or _71797_ (_20083_, _01442_, \oc8051_golden_model_1.PCON [5]);
  and _71798_ (_20084_, _20083_, _43634_);
  and _71799_ (_44137_, _20084_, _20082_);
  and _71800_ (_20086_, _11424_, \oc8051_golden_model_1.PCON [6]);
  nor _71801_ (_20087_, _10595_, _11424_);
  or _71802_ (_20088_, _20087_, _20086_);
  and _71803_ (_20089_, _08042_, \oc8051_golden_model_1.ACC [6]);
  nand _71804_ (_20090_, _20089_, _08212_);
  and _71805_ (_20091_, _20090_, _06615_);
  and _71806_ (_20092_, _20091_, _20088_);
  and _71807_ (_20093_, _15759_, _08042_);
  or _71808_ (_20094_, _20093_, _20086_);
  or _71809_ (_20095_, _20094_, _07275_);
  or _71810_ (_20097_, _20089_, _20086_);
  and _71811_ (_20098_, _20097_, _07259_);
  and _71812_ (_20099_, _07260_, \oc8051_golden_model_1.PCON [6]);
  or _71813_ (_20100_, _20099_, _06474_);
  or _71814_ (_20101_, _20100_, _20098_);
  and _71815_ (_20102_, _20101_, _06772_);
  and _71816_ (_20103_, _20102_, _20095_);
  nor _71817_ (_20104_, _08209_, _11424_);
  or _71818_ (_20105_, _20104_, _20086_);
  and _71819_ (_20106_, _20105_, _06410_);
  or _71820_ (_20108_, _20106_, _20103_);
  and _71821_ (_20109_, _20108_, _06426_);
  and _71822_ (_20110_, _20097_, _06417_);
  or _71823_ (_20111_, _20110_, _10153_);
  or _71824_ (_20112_, _20111_, _20109_);
  or _71825_ (_20113_, _20105_, _06327_);
  and _71826_ (_20114_, _20113_, _20112_);
  or _71827_ (_20115_, _20114_, _09572_);
  and _71828_ (_20116_, _09172_, _08042_);
  or _71829_ (_20117_, _20086_, _06333_);
  or _71830_ (_20119_, _20117_, _20116_);
  and _71831_ (_20120_, _20119_, _06313_);
  and _71832_ (_20121_, _20120_, _20115_);
  and _71833_ (_20122_, _15846_, _08042_);
  or _71834_ (_20123_, _20122_, _20086_);
  and _71835_ (_20124_, _20123_, _06037_);
  or _71836_ (_20125_, _20124_, _06277_);
  or _71837_ (_20126_, _20125_, _20121_);
  and _71838_ (_20127_, _15853_, _08042_);
  or _71839_ (_20128_, _20127_, _20086_);
  or _71840_ (_20130_, _20128_, _06278_);
  and _71841_ (_20131_, _20130_, _20126_);
  or _71842_ (_20132_, _20131_, _06502_);
  and _71843_ (_20133_, _15862_, _08042_);
  or _71844_ (_20134_, _20086_, _07334_);
  or _71845_ (_20135_, _20134_, _20133_);
  and _71846_ (_20136_, _20135_, _07337_);
  and _71847_ (_20137_, _20136_, _20132_);
  or _71848_ (_20138_, _20137_, _20092_);
  and _71849_ (_20139_, _20138_, _07339_);
  or _71850_ (_20141_, _20086_, _08212_);
  and _71851_ (_20142_, _20128_, _06507_);
  and _71852_ (_20143_, _20142_, _20141_);
  or _71853_ (_20144_, _20143_, _20139_);
  and _71854_ (_20145_, _20144_, _07331_);
  and _71855_ (_20146_, _20097_, _06610_);
  and _71856_ (_20147_, _20146_, _20141_);
  or _71857_ (_20148_, _20147_, _06509_);
  or _71858_ (_20149_, _20148_, _20145_);
  and _71859_ (_20150_, _15859_, _08042_);
  or _71860_ (_20152_, _20086_, _09107_);
  or _71861_ (_20153_, _20152_, _20150_);
  and _71862_ (_20154_, _20153_, _09112_);
  and _71863_ (_20155_, _20154_, _20149_);
  and _71864_ (_20156_, _20088_, _06602_);
  or _71865_ (_20157_, _20156_, _06639_);
  or _71866_ (_20158_, _20157_, _20155_);
  or _71867_ (_20159_, _20094_, _07048_);
  and _71868_ (_20160_, _20159_, _06651_);
  and _71869_ (_20161_, _20160_, _20158_);
  and _71870_ (_20163_, _15921_, _08042_);
  or _71871_ (_20164_, _20163_, _20086_);
  and _71872_ (_20165_, _20164_, _06646_);
  or _71873_ (_20166_, _20165_, _01446_);
  or _71874_ (_20167_, _20166_, _20161_);
  or _71875_ (_20168_, _01442_, \oc8051_golden_model_1.PCON [6]);
  and _71876_ (_20169_, _20168_, _43634_);
  and _71877_ (_44138_, _20169_, _20167_);
  and _71878_ (_20170_, _01446_, \oc8051_golden_model_1.TMOD [0]);
  and _71879_ (_20171_, _11502_, \oc8051_golden_model_1.TMOD [0]);
  and _71880_ (_20173_, _07965_, _07250_);
  or _71881_ (_20174_, _20173_, _20171_);
  or _71882_ (_20175_, _20174_, _06327_);
  nor _71883_ (_20176_, _08453_, _11502_);
  or _71884_ (_20177_, _20176_, _20171_);
  or _71885_ (_20178_, _20177_, _07275_);
  and _71886_ (_20179_, _07965_, \oc8051_golden_model_1.ACC [0]);
  or _71887_ (_20180_, _20179_, _20171_);
  and _71888_ (_20181_, _20180_, _07259_);
  and _71889_ (_20182_, _07260_, \oc8051_golden_model_1.TMOD [0]);
  or _71890_ (_20184_, _20182_, _06474_);
  or _71891_ (_20185_, _20184_, _20181_);
  and _71892_ (_20186_, _20185_, _06772_);
  and _71893_ (_20187_, _20186_, _20178_);
  and _71894_ (_20188_, _20174_, _06410_);
  or _71895_ (_20189_, _20188_, _20187_);
  and _71896_ (_20190_, _20189_, _06426_);
  and _71897_ (_20191_, _20180_, _06417_);
  or _71898_ (_20192_, _20191_, _10153_);
  or _71899_ (_20193_, _20192_, _20190_);
  and _71900_ (_20195_, _20193_, _20175_);
  or _71901_ (_20196_, _20195_, _09572_);
  and _71902_ (_20197_, _09447_, _07965_);
  or _71903_ (_20198_, _20171_, _06333_);
  or _71904_ (_20199_, _20198_, _20197_);
  and _71905_ (_20200_, _20199_, _20196_);
  or _71906_ (_20201_, _20200_, _06037_);
  and _71907_ (_20202_, _14666_, _07965_);
  or _71908_ (_20203_, _20171_, _06313_);
  or _71909_ (_20204_, _20203_, _20202_);
  and _71910_ (_20206_, _20204_, _06278_);
  and _71911_ (_20207_, _20206_, _20201_);
  and _71912_ (_20208_, _07965_, _09008_);
  or _71913_ (_20209_, _20208_, _20171_);
  and _71914_ (_20210_, _20209_, _06277_);
  or _71915_ (_20211_, _20210_, _06502_);
  or _71916_ (_20212_, _20211_, _20207_);
  and _71917_ (_20213_, _14566_, _07965_);
  or _71918_ (_20214_, _20171_, _07334_);
  or _71919_ (_20215_, _20214_, _20213_);
  and _71920_ (_20217_, _20215_, _07337_);
  and _71921_ (_20218_, _20217_, _20212_);
  nor _71922_ (_20219_, _12622_, _11502_);
  or _71923_ (_20220_, _20219_, _20171_);
  and _71924_ (_20221_, _10577_, _07965_);
  nor _71925_ (_20222_, _20221_, _07337_);
  and _71926_ (_20223_, _20222_, _20220_);
  or _71927_ (_20224_, _20223_, _20218_);
  and _71928_ (_20225_, _20224_, _07339_);
  nand _71929_ (_20226_, _20209_, _06507_);
  nor _71930_ (_20228_, _20226_, _20176_);
  or _71931_ (_20229_, _20228_, _06610_);
  or _71932_ (_20230_, _20229_, _20225_);
  or _71933_ (_20231_, _20221_, _20171_);
  or _71934_ (_20232_, _20231_, _07331_);
  and _71935_ (_20233_, _20232_, _20230_);
  or _71936_ (_20234_, _20233_, _06509_);
  and _71937_ (_20235_, _14563_, _07965_);
  or _71938_ (_20236_, _20171_, _09107_);
  or _71939_ (_20237_, _20236_, _20235_);
  and _71940_ (_20239_, _20237_, _09112_);
  and _71941_ (_20240_, _20239_, _20234_);
  and _71942_ (_20241_, _20220_, _06602_);
  or _71943_ (_20242_, _20241_, _19642_);
  or _71944_ (_20243_, _20242_, _20240_);
  or _71945_ (_20244_, _20177_, _19641_);
  and _71946_ (_20245_, _20244_, _01442_);
  and _71947_ (_20246_, _20245_, _20243_);
  or _71948_ (_20247_, _20246_, _20170_);
  and _71949_ (_44140_, _20247_, _43634_);
  not _71950_ (_20249_, \oc8051_golden_model_1.TMOD [1]);
  nor _71951_ (_20250_, _01442_, _20249_);
  or _71952_ (_20251_, _14851_, _11502_);
  or _71953_ (_20252_, _07965_, \oc8051_golden_model_1.TMOD [1]);
  and _71954_ (_20253_, _20252_, _06037_);
  and _71955_ (_20254_, _20253_, _20251_);
  and _71956_ (_20255_, _14744_, _07965_);
  not _71957_ (_20256_, _20255_);
  and _71958_ (_20257_, _20256_, _20252_);
  or _71959_ (_20258_, _20257_, _07275_);
  nor _71960_ (_20260_, _07965_, _20249_);
  and _71961_ (_20261_, _07965_, \oc8051_golden_model_1.ACC [1]);
  or _71962_ (_20262_, _20261_, _20260_);
  and _71963_ (_20263_, _20262_, _07259_);
  nor _71964_ (_20264_, _07259_, _20249_);
  or _71965_ (_20265_, _20264_, _06474_);
  or _71966_ (_20266_, _20265_, _20263_);
  and _71967_ (_20267_, _20266_, _06772_);
  and _71968_ (_20268_, _20267_, _20258_);
  nor _71969_ (_20269_, _11502_, _07448_);
  or _71970_ (_20271_, _20269_, _20260_);
  and _71971_ (_20272_, _20271_, _06410_);
  or _71972_ (_20273_, _20272_, _20268_);
  and _71973_ (_20274_, _20273_, _06426_);
  and _71974_ (_20275_, _20262_, _06417_);
  or _71975_ (_20276_, _20275_, _10153_);
  or _71976_ (_20277_, _20276_, _20274_);
  or _71977_ (_20278_, _20271_, _06327_);
  and _71978_ (_20279_, _20278_, _16672_);
  and _71979_ (_20280_, _20279_, _20277_);
  or _71980_ (_20282_, _09402_, _11502_);
  and _71981_ (_20283_, _20252_, _14025_);
  and _71982_ (_20284_, _20283_, _20282_);
  or _71983_ (_20285_, _20284_, _20280_);
  and _71984_ (_20286_, _20285_, _06313_);
  or _71985_ (_20287_, _20286_, _20254_);
  and _71986_ (_20288_, _20287_, _06278_);
  nand _71987_ (_20289_, _07965_, _07160_);
  and _71988_ (_20290_, _20252_, _06277_);
  and _71989_ (_20291_, _20290_, _20289_);
  or _71990_ (_20293_, _20291_, _20288_);
  and _71991_ (_20294_, _20293_, _07334_);
  or _71992_ (_20295_, _14749_, _11502_);
  and _71993_ (_20296_, _20252_, _06502_);
  and _71994_ (_20297_, _20296_, _20295_);
  or _71995_ (_20298_, _20297_, _06615_);
  or _71996_ (_20299_, _20298_, _20294_);
  nor _71997_ (_20300_, _10578_, _11502_);
  or _71998_ (_20301_, _20300_, _20260_);
  nand _71999_ (_20302_, _10576_, _07965_);
  and _72000_ (_20304_, _20302_, _20301_);
  or _72001_ (_20305_, _20304_, _07337_);
  and _72002_ (_20306_, _20305_, _07339_);
  and _72003_ (_20307_, _20306_, _20299_);
  or _72004_ (_20308_, _14747_, _11502_);
  and _72005_ (_20309_, _20252_, _06507_);
  and _72006_ (_20310_, _20309_, _20308_);
  or _72007_ (_20311_, _20310_, _06610_);
  or _72008_ (_20312_, _20311_, _20307_);
  nor _72009_ (_20313_, _20260_, _07331_);
  nand _72010_ (_20315_, _20313_, _20302_);
  and _72011_ (_20316_, _20315_, _09107_);
  and _72012_ (_20317_, _20316_, _20312_);
  or _72013_ (_20318_, _20289_, _08404_);
  and _72014_ (_20319_, _20252_, _06509_);
  and _72015_ (_20320_, _20319_, _20318_);
  or _72016_ (_20321_, _20320_, _06602_);
  or _72017_ (_20322_, _20321_, _20317_);
  or _72018_ (_20323_, _20301_, _09112_);
  and _72019_ (_20324_, _20323_, _07048_);
  and _72020_ (_20326_, _20324_, _20322_);
  and _72021_ (_20327_, _20257_, _06639_);
  or _72022_ (_20328_, _20327_, _06646_);
  or _72023_ (_20329_, _20328_, _20326_);
  or _72024_ (_20330_, _20260_, _06651_);
  or _72025_ (_20331_, _20330_, _20255_);
  and _72026_ (_20332_, _20331_, _01442_);
  and _72027_ (_20333_, _20332_, _20329_);
  or _72028_ (_20334_, _20333_, _20250_);
  and _72029_ (_44141_, _20334_, _43634_);
  and _72030_ (_20336_, _01446_, \oc8051_golden_model_1.TMOD [2]);
  and _72031_ (_20337_, _11502_, \oc8051_golden_model_1.TMOD [2]);
  and _72032_ (_20338_, _09356_, _07965_);
  or _72033_ (_20339_, _20338_, _20337_);
  and _72034_ (_20340_, _20339_, _14025_);
  and _72035_ (_20341_, _14959_, _07965_);
  or _72036_ (_20342_, _20341_, _20337_);
  or _72037_ (_20343_, _20342_, _07275_);
  and _72038_ (_20344_, _07965_, \oc8051_golden_model_1.ACC [2]);
  or _72039_ (_20345_, _20344_, _20337_);
  and _72040_ (_20347_, _20345_, _07259_);
  and _72041_ (_20348_, _07260_, \oc8051_golden_model_1.TMOD [2]);
  or _72042_ (_20349_, _20348_, _06474_);
  or _72043_ (_20350_, _20349_, _20347_);
  and _72044_ (_20351_, _20350_, _06772_);
  and _72045_ (_20352_, _20351_, _20343_);
  nor _72046_ (_20353_, _11502_, _07854_);
  or _72047_ (_20354_, _20353_, _20337_);
  and _72048_ (_20355_, _20354_, _06410_);
  or _72049_ (_20356_, _20355_, _20352_);
  and _72050_ (_20358_, _20356_, _06426_);
  and _72051_ (_20359_, _20345_, _06417_);
  or _72052_ (_20360_, _20359_, _10153_);
  or _72053_ (_20361_, _20360_, _20358_);
  or _72054_ (_20362_, _20354_, _06327_);
  and _72055_ (_20363_, _20362_, _16672_);
  and _72056_ (_20364_, _20363_, _20361_);
  or _72057_ (_20365_, _20364_, _06037_);
  or _72058_ (_20366_, _20365_, _20340_);
  and _72059_ (_20367_, _15056_, _07965_);
  or _72060_ (_20369_, _20337_, _06313_);
  or _72061_ (_20370_, _20369_, _20367_);
  and _72062_ (_20371_, _20370_, _06278_);
  and _72063_ (_20372_, _20371_, _20366_);
  and _72064_ (_20373_, _07965_, _09057_);
  or _72065_ (_20374_, _20373_, _20337_);
  and _72066_ (_20375_, _20374_, _06277_);
  or _72067_ (_20376_, _20375_, _06502_);
  or _72068_ (_20377_, _20376_, _20372_);
  and _72069_ (_20378_, _14948_, _07965_);
  or _72070_ (_20380_, _20337_, _07334_);
  or _72071_ (_20381_, _20380_, _20378_);
  and _72072_ (_20382_, _20381_, _07337_);
  and _72073_ (_20383_, _20382_, _20377_);
  and _72074_ (_20384_, _10583_, _07965_);
  or _72075_ (_20385_, _20384_, _20337_);
  and _72076_ (_20386_, _20385_, _06615_);
  or _72077_ (_20387_, _20386_, _20383_);
  and _72078_ (_20388_, _20387_, _07339_);
  or _72079_ (_20389_, _20337_, _08503_);
  and _72080_ (_20391_, _20374_, _06507_);
  and _72081_ (_20392_, _20391_, _20389_);
  or _72082_ (_20393_, _20392_, _20388_);
  and _72083_ (_20394_, _20393_, _07331_);
  and _72084_ (_20395_, _20345_, _06610_);
  and _72085_ (_20396_, _20395_, _20389_);
  or _72086_ (_20397_, _20396_, _06509_);
  or _72087_ (_20398_, _20397_, _20394_);
  and _72088_ (_20399_, _14945_, _07965_);
  or _72089_ (_20400_, _20337_, _09107_);
  or _72090_ (_20402_, _20400_, _20399_);
  and _72091_ (_20403_, _20402_, _09112_);
  and _72092_ (_20404_, _20403_, _20398_);
  nor _72093_ (_20405_, _10582_, _11502_);
  or _72094_ (_20406_, _20405_, _20337_);
  and _72095_ (_20407_, _20406_, _06602_);
  or _72096_ (_20408_, _20407_, _20404_);
  and _72097_ (_20409_, _20408_, _07048_);
  and _72098_ (_20410_, _20342_, _06639_);
  or _72099_ (_20411_, _20410_, _06646_);
  or _72100_ (_20413_, _20411_, _20409_);
  and _72101_ (_20414_, _15129_, _07965_);
  or _72102_ (_20415_, _20337_, _06651_);
  or _72103_ (_20416_, _20415_, _20414_);
  and _72104_ (_20417_, _20416_, _01442_);
  and _72105_ (_20418_, _20417_, _20413_);
  or _72106_ (_20419_, _20418_, _20336_);
  and _72107_ (_44142_, _20419_, _43634_);
  and _72108_ (_20420_, _11502_, \oc8051_golden_model_1.TMOD [3]);
  or _72109_ (_20421_, _20420_, _08359_);
  and _72110_ (_20423_, _07965_, _09014_);
  or _72111_ (_20424_, _20423_, _20420_);
  and _72112_ (_20425_, _20424_, _06507_);
  and _72113_ (_20426_, _20425_, _20421_);
  and _72114_ (_20427_, _15153_, _07965_);
  or _72115_ (_20428_, _20427_, _20420_);
  or _72116_ (_20429_, _20428_, _07275_);
  and _72117_ (_20430_, _07965_, \oc8051_golden_model_1.ACC [3]);
  or _72118_ (_20431_, _20430_, _20420_);
  and _72119_ (_20432_, _20431_, _07259_);
  and _72120_ (_20434_, _07260_, \oc8051_golden_model_1.TMOD [3]);
  or _72121_ (_20435_, _20434_, _06474_);
  or _72122_ (_20436_, _20435_, _20432_);
  and _72123_ (_20437_, _20436_, _06772_);
  and _72124_ (_20438_, _20437_, _20429_);
  nor _72125_ (_20439_, _11502_, _07680_);
  or _72126_ (_20440_, _20439_, _20420_);
  and _72127_ (_20441_, _20440_, _06410_);
  or _72128_ (_20442_, _20441_, _20438_);
  and _72129_ (_20443_, _20442_, _06426_);
  and _72130_ (_20445_, _20431_, _06417_);
  or _72131_ (_20446_, _20445_, _10153_);
  or _72132_ (_20447_, _20446_, _20443_);
  or _72133_ (_20448_, _20440_, _06327_);
  and _72134_ (_20449_, _20448_, _20447_);
  or _72135_ (_20450_, _20449_, _09572_);
  and _72136_ (_20451_, _09310_, _07965_);
  or _72137_ (_20452_, _20420_, _06333_);
  or _72138_ (_20453_, _20452_, _20451_);
  and _72139_ (_20454_, _20453_, _06313_);
  and _72140_ (_20456_, _20454_, _20450_);
  and _72141_ (_20457_, _15251_, _07965_);
  or _72142_ (_20458_, _20457_, _20420_);
  and _72143_ (_20459_, _20458_, _06037_);
  or _72144_ (_20460_, _20459_, _06277_);
  or _72145_ (_20461_, _20460_, _20456_);
  or _72146_ (_20462_, _20424_, _06278_);
  and _72147_ (_20463_, _20462_, _20461_);
  or _72148_ (_20464_, _20463_, _06502_);
  and _72149_ (_20465_, _15266_, _07965_);
  or _72150_ (_20467_, _20420_, _07334_);
  or _72151_ (_20468_, _20467_, _20465_);
  and _72152_ (_20469_, _20468_, _07337_);
  and _72153_ (_20470_, _20469_, _20464_);
  and _72154_ (_20471_, _12619_, _07965_);
  or _72155_ (_20472_, _20471_, _20420_);
  and _72156_ (_20473_, _20472_, _06615_);
  or _72157_ (_20474_, _20473_, _20470_);
  and _72158_ (_20475_, _20474_, _07339_);
  or _72159_ (_20476_, _20475_, _20426_);
  and _72160_ (_20478_, _20476_, _07331_);
  and _72161_ (_20479_, _20431_, _06610_);
  and _72162_ (_20480_, _20479_, _20421_);
  or _72163_ (_20481_, _20480_, _06509_);
  or _72164_ (_20482_, _20481_, _20478_);
  and _72165_ (_20483_, _15263_, _07965_);
  or _72166_ (_20484_, _20420_, _09107_);
  or _72167_ (_20485_, _20484_, _20483_);
  and _72168_ (_20486_, _20485_, _09112_);
  and _72169_ (_20487_, _20486_, _20482_);
  nor _72170_ (_20489_, _10574_, _11502_);
  or _72171_ (_20490_, _20489_, _20420_);
  and _72172_ (_20491_, _20490_, _06602_);
  or _72173_ (_20492_, _20491_, _06639_);
  or _72174_ (_20493_, _20492_, _20487_);
  or _72175_ (_20494_, _20428_, _07048_);
  and _72176_ (_20495_, _20494_, _06651_);
  and _72177_ (_20496_, _20495_, _20493_);
  and _72178_ (_20497_, _15321_, _07965_);
  or _72179_ (_20498_, _20497_, _20420_);
  and _72180_ (_20500_, _20498_, _06646_);
  or _72181_ (_20501_, _20500_, _01446_);
  or _72182_ (_20502_, _20501_, _20496_);
  or _72183_ (_20503_, _01442_, \oc8051_golden_model_1.TMOD [3]);
  and _72184_ (_20504_, _20503_, _43634_);
  and _72185_ (_44144_, _20504_, _20502_);
  and _72186_ (_20505_, _11502_, \oc8051_golden_model_1.TMOD [4]);
  or _72187_ (_20506_, _20505_, _08599_);
  and _72188_ (_20507_, _08995_, _07965_);
  or _72189_ (_20508_, _20507_, _20505_);
  and _72190_ (_20510_, _20508_, _06507_);
  and _72191_ (_20511_, _20510_, _20506_);
  nor _72192_ (_20512_, _10589_, _11502_);
  or _72193_ (_20513_, _20512_, _20505_);
  and _72194_ (_20514_, _07965_, \oc8051_golden_model_1.ACC [4]);
  nand _72195_ (_20515_, _20514_, _08599_);
  and _72196_ (_20516_, _20515_, _06615_);
  and _72197_ (_20517_, _20516_, _20513_);
  nor _72198_ (_20518_, _08596_, _11502_);
  or _72199_ (_20519_, _20518_, _20505_);
  or _72200_ (_20521_, _20519_, _06327_);
  and _72201_ (_20522_, _15367_, _07965_);
  or _72202_ (_20523_, _20522_, _20505_);
  or _72203_ (_20524_, _20523_, _07275_);
  or _72204_ (_20525_, _20514_, _20505_);
  and _72205_ (_20526_, _20525_, _07259_);
  and _72206_ (_20527_, _07260_, \oc8051_golden_model_1.TMOD [4]);
  or _72207_ (_20528_, _20527_, _06474_);
  or _72208_ (_20529_, _20528_, _20526_);
  and _72209_ (_20530_, _20529_, _06772_);
  and _72210_ (_20532_, _20530_, _20524_);
  and _72211_ (_20533_, _20519_, _06410_);
  or _72212_ (_20534_, _20533_, _20532_);
  and _72213_ (_20535_, _20534_, _06426_);
  and _72214_ (_20536_, _20525_, _06417_);
  or _72215_ (_20537_, _20536_, _10153_);
  or _72216_ (_20538_, _20537_, _20535_);
  and _72217_ (_20539_, _20538_, _20521_);
  or _72218_ (_20540_, _20539_, _09572_);
  and _72219_ (_20541_, _09264_, _07965_);
  or _72220_ (_20543_, _20505_, _16672_);
  or _72221_ (_20544_, _20543_, _20541_);
  and _72222_ (_20545_, _20544_, _20540_);
  or _72223_ (_20546_, _20545_, _06037_);
  and _72224_ (_20547_, _15452_, _07965_);
  or _72225_ (_20548_, _20505_, _06313_);
  or _72226_ (_20549_, _20548_, _20547_);
  and _72227_ (_20550_, _20549_, _06278_);
  and _72228_ (_20551_, _20550_, _20546_);
  and _72229_ (_20552_, _20508_, _06277_);
  or _72230_ (_20554_, _20552_, _06502_);
  or _72231_ (_20555_, _20554_, _20551_);
  and _72232_ (_20556_, _15345_, _07965_);
  or _72233_ (_20557_, _20505_, _07334_);
  or _72234_ (_20558_, _20557_, _20556_);
  and _72235_ (_20559_, _20558_, _07337_);
  and _72236_ (_20560_, _20559_, _20555_);
  or _72237_ (_20561_, _20560_, _20517_);
  and _72238_ (_20562_, _20561_, _07339_);
  or _72239_ (_20563_, _20562_, _20511_);
  and _72240_ (_20565_, _20563_, _07331_);
  and _72241_ (_20566_, _20525_, _06610_);
  and _72242_ (_20567_, _20566_, _20506_);
  or _72243_ (_20568_, _20567_, _06509_);
  or _72244_ (_20569_, _20568_, _20565_);
  and _72245_ (_20570_, _15342_, _07965_);
  or _72246_ (_20571_, _20505_, _09107_);
  or _72247_ (_20572_, _20571_, _20570_);
  and _72248_ (_20573_, _20572_, _09112_);
  and _72249_ (_20574_, _20573_, _20569_);
  and _72250_ (_20576_, _20513_, _06602_);
  or _72251_ (_20577_, _20576_, _06639_);
  or _72252_ (_20578_, _20577_, _20574_);
  or _72253_ (_20579_, _20523_, _07048_);
  and _72254_ (_20580_, _20579_, _06651_);
  and _72255_ (_20581_, _20580_, _20578_);
  and _72256_ (_20582_, _15524_, _07965_);
  or _72257_ (_20583_, _20582_, _20505_);
  and _72258_ (_20584_, _20583_, _06646_);
  or _72259_ (_20585_, _20584_, _01446_);
  or _72260_ (_20587_, _20585_, _20581_);
  or _72261_ (_20588_, _01442_, \oc8051_golden_model_1.TMOD [4]);
  and _72262_ (_20589_, _20588_, _43634_);
  and _72263_ (_44145_, _20589_, _20587_);
  and _72264_ (_20590_, _11502_, \oc8051_golden_model_1.TMOD [5]);
  nor _72265_ (_20591_, _10570_, _11502_);
  or _72266_ (_20592_, _20591_, _20590_);
  and _72267_ (_20593_, _07965_, \oc8051_golden_model_1.ACC [5]);
  nand _72268_ (_20594_, _20593_, _08308_);
  and _72269_ (_20595_, _20594_, _06615_);
  and _72270_ (_20597_, _20595_, _20592_);
  nor _72271_ (_20598_, _08305_, _11502_);
  or _72272_ (_20599_, _20598_, _20590_);
  or _72273_ (_20600_, _20599_, _06327_);
  and _72274_ (_20601_, _15550_, _07965_);
  or _72275_ (_20602_, _20601_, _20590_);
  or _72276_ (_20603_, _20602_, _07275_);
  or _72277_ (_20604_, _20593_, _20590_);
  and _72278_ (_20605_, _20604_, _07259_);
  and _72279_ (_20606_, _07260_, \oc8051_golden_model_1.TMOD [5]);
  or _72280_ (_20608_, _20606_, _06474_);
  or _72281_ (_20609_, _20608_, _20605_);
  and _72282_ (_20610_, _20609_, _06772_);
  and _72283_ (_20611_, _20610_, _20603_);
  and _72284_ (_20612_, _20599_, _06410_);
  or _72285_ (_20613_, _20612_, _20611_);
  and _72286_ (_20614_, _20613_, _06426_);
  and _72287_ (_20615_, _20604_, _06417_);
  or _72288_ (_20616_, _20615_, _10153_);
  or _72289_ (_20617_, _20616_, _20614_);
  and _72290_ (_20619_, _20617_, _20600_);
  or _72291_ (_20620_, _20619_, _09572_);
  and _72292_ (_20621_, _09218_, _07965_);
  or _72293_ (_20622_, _20590_, _06333_);
  or _72294_ (_20623_, _20622_, _20621_);
  and _72295_ (_20624_, _20623_, _06313_);
  and _72296_ (_20625_, _20624_, _20620_);
  and _72297_ (_20626_, _15649_, _07965_);
  or _72298_ (_20627_, _20626_, _20590_);
  and _72299_ (_20628_, _20627_, _06037_);
  or _72300_ (_20629_, _20628_, _06277_);
  or _72301_ (_20630_, _20629_, _20625_);
  and _72302_ (_20631_, _08954_, _07965_);
  or _72303_ (_20632_, _20631_, _20590_);
  or _72304_ (_20633_, _20632_, _06278_);
  and _72305_ (_20634_, _20633_, _20630_);
  or _72306_ (_20635_, _20634_, _06502_);
  and _72307_ (_20636_, _15664_, _07965_);
  or _72308_ (_20637_, _20590_, _07334_);
  or _72309_ (_20638_, _20637_, _20636_);
  and _72310_ (_20641_, _20638_, _07337_);
  and _72311_ (_20642_, _20641_, _20635_);
  or _72312_ (_20643_, _20642_, _20597_);
  and _72313_ (_20644_, _20643_, _07339_);
  or _72314_ (_20645_, _20590_, _08308_);
  and _72315_ (_20646_, _20632_, _06507_);
  and _72316_ (_20647_, _20646_, _20645_);
  or _72317_ (_20648_, _20647_, _20644_);
  and _72318_ (_20649_, _20648_, _07331_);
  and _72319_ (_20650_, _20604_, _06610_);
  and _72320_ (_20652_, _20650_, _20645_);
  or _72321_ (_20653_, _20652_, _06509_);
  or _72322_ (_20654_, _20653_, _20649_);
  and _72323_ (_20655_, _15663_, _07965_);
  or _72324_ (_20656_, _20590_, _09107_);
  or _72325_ (_20657_, _20656_, _20655_);
  and _72326_ (_20658_, _20657_, _09112_);
  and _72327_ (_20659_, _20658_, _20654_);
  and _72328_ (_20660_, _20592_, _06602_);
  or _72329_ (_20661_, _20660_, _06639_);
  or _72330_ (_20663_, _20661_, _20659_);
  or _72331_ (_20664_, _20602_, _07048_);
  and _72332_ (_20665_, _20664_, _06651_);
  and _72333_ (_20666_, _20665_, _20663_);
  and _72334_ (_20667_, _15721_, _07965_);
  or _72335_ (_20668_, _20667_, _20590_);
  and _72336_ (_20669_, _20668_, _06646_);
  or _72337_ (_20670_, _20669_, _01446_);
  or _72338_ (_20671_, _20670_, _20666_);
  or _72339_ (_20672_, _01442_, \oc8051_golden_model_1.TMOD [5]);
  and _72340_ (_20673_, _20672_, _43634_);
  and _72341_ (_44146_, _20673_, _20671_);
  and _72342_ (_20674_, _11502_, \oc8051_golden_model_1.TMOD [6]);
  and _72343_ (_20675_, _15759_, _07965_);
  or _72344_ (_20676_, _20675_, _20674_);
  or _72345_ (_20677_, _20676_, _07275_);
  and _72346_ (_20678_, _07965_, \oc8051_golden_model_1.ACC [6]);
  or _72347_ (_20679_, _20678_, _20674_);
  and _72348_ (_20680_, _20679_, _07259_);
  and _72349_ (_20681_, _07260_, \oc8051_golden_model_1.TMOD [6]);
  or _72350_ (_20684_, _20681_, _06474_);
  or _72351_ (_20685_, _20684_, _20680_);
  and _72352_ (_20686_, _20685_, _06772_);
  and _72353_ (_20687_, _20686_, _20677_);
  nor _72354_ (_20688_, _08209_, _11502_);
  or _72355_ (_20689_, _20688_, _20674_);
  and _72356_ (_20690_, _20689_, _06410_);
  or _72357_ (_20691_, _20690_, _20687_);
  and _72358_ (_20692_, _20691_, _06426_);
  and _72359_ (_20693_, _20679_, _06417_);
  or _72360_ (_20695_, _20693_, _10153_);
  or _72361_ (_20696_, _20695_, _20692_);
  or _72362_ (_20697_, _20689_, _06327_);
  and _72363_ (_20698_, _20697_, _20696_);
  or _72364_ (_20699_, _20698_, _09572_);
  and _72365_ (_20700_, _09172_, _07965_);
  or _72366_ (_20701_, _20674_, _06333_);
  or _72367_ (_20702_, _20701_, _20700_);
  and _72368_ (_20703_, _20702_, _06313_);
  and _72369_ (_20704_, _20703_, _20699_);
  and _72370_ (_20705_, _15846_, _07965_);
  or _72371_ (_20706_, _20705_, _20674_);
  and _72372_ (_20707_, _20706_, _06037_);
  or _72373_ (_20708_, _20707_, _06277_);
  or _72374_ (_20709_, _20708_, _20704_);
  and _72375_ (_20710_, _15853_, _07965_);
  or _72376_ (_20711_, _20710_, _20674_);
  or _72377_ (_20712_, _20711_, _06278_);
  and _72378_ (_20713_, _20712_, _20709_);
  or _72379_ (_20714_, _20713_, _06502_);
  and _72380_ (_20717_, _15862_, _07965_);
  or _72381_ (_20718_, _20674_, _07334_);
  or _72382_ (_20719_, _20718_, _20717_);
  and _72383_ (_20720_, _20719_, _07337_);
  and _72384_ (_20721_, _20720_, _20714_);
  and _72385_ (_20722_, _10596_, _07965_);
  or _72386_ (_20723_, _20722_, _20674_);
  and _72387_ (_20724_, _20723_, _06615_);
  or _72388_ (_20725_, _20724_, _20721_);
  and _72389_ (_20726_, _20725_, _07339_);
  or _72390_ (_20728_, _20674_, _08212_);
  and _72391_ (_20729_, _20711_, _06507_);
  and _72392_ (_20730_, _20729_, _20728_);
  or _72393_ (_20731_, _20730_, _20726_);
  and _72394_ (_20732_, _20731_, _07331_);
  and _72395_ (_20733_, _20679_, _06610_);
  and _72396_ (_20734_, _20733_, _20728_);
  or _72397_ (_20735_, _20734_, _06509_);
  or _72398_ (_20736_, _20735_, _20732_);
  and _72399_ (_20737_, _15859_, _07965_);
  or _72400_ (_20739_, _20674_, _09107_);
  or _72401_ (_20740_, _20739_, _20737_);
  and _72402_ (_20741_, _20740_, _09112_);
  and _72403_ (_20742_, _20741_, _20736_);
  nor _72404_ (_20743_, _10595_, _11502_);
  or _72405_ (_20744_, _20743_, _20674_);
  and _72406_ (_20745_, _20744_, _06602_);
  or _72407_ (_20746_, _20745_, _06639_);
  or _72408_ (_20747_, _20746_, _20742_);
  or _72409_ (_20748_, _20676_, _07048_);
  and _72410_ (_20750_, _20748_, _06651_);
  and _72411_ (_20751_, _20750_, _20747_);
  and _72412_ (_20752_, _15921_, _07965_);
  or _72413_ (_20753_, _20752_, _20674_);
  and _72414_ (_20754_, _20753_, _06646_);
  or _72415_ (_20755_, _20754_, _01446_);
  or _72416_ (_20756_, _20755_, _20751_);
  or _72417_ (_20757_, _01442_, \oc8051_golden_model_1.TMOD [6]);
  and _72418_ (_20758_, _20757_, _43634_);
  and _72419_ (_44147_, _20758_, _20756_);
  not _72420_ (_20759_, \oc8051_golden_model_1.DPL [0]);
  nor _72421_ (_20760_, _01442_, _20759_);
  nor _72422_ (_20761_, _08001_, _20759_);
  and _72423_ (_20762_, _08001_, _07250_);
  or _72424_ (_20763_, _20762_, _20761_);
  or _72425_ (_20764_, _20763_, _06327_);
  and _72426_ (_20765_, _08158_, \oc8051_golden_model_1.ACC [0]);
  or _72427_ (_20766_, _20765_, _20761_);
  or _72428_ (_20767_, _20766_, _06426_);
  nor _72429_ (_20768_, _08453_, _11585_);
  or _72430_ (_20771_, _20768_, _20761_);
  or _72431_ (_20772_, _20771_, _07275_);
  and _72432_ (_20773_, _20766_, _07259_);
  nor _72433_ (_20774_, _07259_, _20759_);
  or _72434_ (_20775_, _20774_, _06474_);
  or _72435_ (_20776_, _20775_, _20773_);
  and _72436_ (_20777_, _20776_, _06772_);
  and _72437_ (_20778_, _20777_, _20772_);
  and _72438_ (_20779_, _20763_, _06410_);
  or _72439_ (_20780_, _20779_, _06417_);
  or _72440_ (_20782_, _20780_, _20778_);
  and _72441_ (_20783_, _20782_, _20767_);
  or _72442_ (_20784_, _20783_, _11603_);
  nand _72443_ (_20785_, _11603_, \oc8051_golden_model_1.DPL [0]);
  and _72444_ (_20786_, _20785_, _06487_);
  and _72445_ (_20787_, _20786_, _20784_);
  nor _72446_ (_20788_, _06950_, _06487_);
  or _72447_ (_20789_, _20788_, _10153_);
  or _72448_ (_20790_, _20789_, _20787_);
  and _72449_ (_20791_, _20790_, _20764_);
  or _72450_ (_20793_, _20791_, _09572_);
  and _72451_ (_20794_, _09447_, _08158_);
  or _72452_ (_20795_, _20761_, _06333_);
  or _72453_ (_20796_, _20795_, _20794_);
  and _72454_ (_20797_, _20796_, _20793_);
  or _72455_ (_20798_, _20797_, _06037_);
  and _72456_ (_20799_, _14666_, _08001_);
  or _72457_ (_20800_, _20761_, _06313_);
  or _72458_ (_20801_, _20800_, _20799_);
  and _72459_ (_20802_, _20801_, _06278_);
  and _72460_ (_20804_, _20802_, _20798_);
  and _72461_ (_20805_, _08158_, _09008_);
  or _72462_ (_20806_, _20805_, _20761_);
  and _72463_ (_20807_, _20806_, _06277_);
  or _72464_ (_20808_, _20807_, _06502_);
  or _72465_ (_20809_, _20808_, _20804_);
  and _72466_ (_20810_, _14566_, _08001_);
  or _72467_ (_20811_, _20761_, _07334_);
  or _72468_ (_20812_, _20811_, _20810_);
  and _72469_ (_20813_, _20812_, _07337_);
  and _72470_ (_20815_, _20813_, _20809_);
  nor _72471_ (_20816_, _12622_, _11585_);
  or _72472_ (_20817_, _20816_, _20761_);
  and _72473_ (_20818_, _20765_, _08453_);
  nor _72474_ (_20819_, _20818_, _07337_);
  and _72475_ (_20820_, _20819_, _20817_);
  or _72476_ (_20821_, _20820_, _20815_);
  and _72477_ (_20822_, _20821_, _07339_);
  nand _72478_ (_20823_, _20806_, _06507_);
  nor _72479_ (_20824_, _20823_, _20768_);
  or _72480_ (_20826_, _20824_, _06610_);
  or _72481_ (_20827_, _20826_, _20822_);
  or _72482_ (_20828_, _20818_, _20761_);
  or _72483_ (_20829_, _20828_, _07331_);
  and _72484_ (_20830_, _20829_, _20827_);
  or _72485_ (_20831_, _20830_, _06509_);
  and _72486_ (_20832_, _14563_, _08001_);
  or _72487_ (_20833_, _20761_, _09107_);
  or _72488_ (_20834_, _20833_, _20832_);
  and _72489_ (_20835_, _20834_, _09112_);
  and _72490_ (_20837_, _20835_, _20831_);
  and _72491_ (_20838_, _20817_, _06602_);
  or _72492_ (_20839_, _20838_, _19642_);
  or _72493_ (_20840_, _20839_, _20837_);
  or _72494_ (_20841_, _20771_, _19641_);
  and _72495_ (_20842_, _20841_, _01442_);
  and _72496_ (_20843_, _20842_, _20840_);
  or _72497_ (_20844_, _20843_, _20760_);
  and _72498_ (_44149_, _20844_, _43634_);
  and _72499_ (_20845_, _01446_, \oc8051_golden_model_1.DPL [1]);
  or _72500_ (_20847_, _09402_, _11585_);
  or _72501_ (_20848_, _08001_, \oc8051_golden_model_1.DPL [1]);
  and _72502_ (_20849_, _20848_, _14025_);
  and _72503_ (_20850_, _20849_, _20847_);
  nor _72504_ (_20851_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _72505_ (_20852_, _20851_, _11608_);
  and _72506_ (_20853_, _20852_, _11603_);
  nand _72507_ (_20854_, _14744_, _08001_);
  and _72508_ (_20855_, _20854_, _20848_);
  or _72509_ (_20856_, _20855_, _07275_);
  and _72510_ (_20858_, _11585_, \oc8051_golden_model_1.DPL [1]);
  and _72511_ (_20859_, _08158_, \oc8051_golden_model_1.ACC [1]);
  or _72512_ (_20860_, _20859_, _20858_);
  and _72513_ (_20861_, _20860_, _07259_);
  and _72514_ (_20862_, _07260_, \oc8051_golden_model_1.DPL [1]);
  or _72515_ (_20863_, _20862_, _06474_);
  or _72516_ (_20864_, _20863_, _20861_);
  and _72517_ (_20865_, _20864_, _06772_);
  and _72518_ (_20866_, _20865_, _20856_);
  nor _72519_ (_20867_, _11585_, _07448_);
  or _72520_ (_20869_, _20867_, _20858_);
  and _72521_ (_20870_, _20869_, _06410_);
  or _72522_ (_20871_, _20870_, _06417_);
  or _72523_ (_20872_, _20871_, _20866_);
  or _72524_ (_20873_, _20860_, _06426_);
  and _72525_ (_20874_, _20873_, _11604_);
  and _72526_ (_20875_, _20874_, _20872_);
  or _72527_ (_20876_, _20875_, _20853_);
  and _72528_ (_20877_, _20876_, _06487_);
  nor _72529_ (_20878_, _07160_, _06487_);
  or _72530_ (_20880_, _20878_, _10153_);
  or _72531_ (_20881_, _20880_, _20877_);
  or _72532_ (_20882_, _20869_, _06327_);
  and _72533_ (_20883_, _20882_, _16672_);
  and _72534_ (_20884_, _20883_, _20881_);
  or _72535_ (_20885_, _20884_, _20850_);
  and _72536_ (_20886_, _20885_, _06313_);
  and _72537_ (_20887_, _14851_, _08158_);
  or _72538_ (_20888_, _20887_, _20858_);
  and _72539_ (_20889_, _20888_, _06037_);
  or _72540_ (_20890_, _20889_, _20886_);
  and _72541_ (_20891_, _20890_, _06278_);
  and _72542_ (_20892_, _20848_, _06277_);
  nand _72543_ (_20893_, _08001_, _07160_);
  and _72544_ (_20894_, _20893_, _20892_);
  or _72545_ (_20895_, _20894_, _20891_);
  and _72546_ (_20896_, _20895_, _07334_);
  or _72547_ (_20897_, _14749_, _11585_);
  and _72548_ (_20898_, _20848_, _06502_);
  and _72549_ (_20899_, _20898_, _20897_);
  or _72550_ (_20902_, _20899_, _06615_);
  or _72551_ (_20903_, _20902_, _20896_);
  nor _72552_ (_20904_, _10578_, _11585_);
  or _72553_ (_20905_, _20904_, _20858_);
  nand _72554_ (_20906_, _10576_, _08001_);
  and _72555_ (_20907_, _20906_, _20905_);
  or _72556_ (_20908_, _20907_, _07337_);
  and _72557_ (_20909_, _20908_, _07339_);
  and _72558_ (_20910_, _20909_, _20903_);
  or _72559_ (_20911_, _14747_, _11585_);
  and _72560_ (_20913_, _20848_, _06507_);
  and _72561_ (_20914_, _20913_, _20911_);
  or _72562_ (_20915_, _20914_, _06610_);
  or _72563_ (_20916_, _20915_, _20910_);
  nor _72564_ (_20917_, _20858_, _07331_);
  nand _72565_ (_20918_, _20917_, _20906_);
  and _72566_ (_20919_, _20918_, _09107_);
  and _72567_ (_20920_, _20919_, _20916_);
  or _72568_ (_20921_, _20893_, _08404_);
  and _72569_ (_20922_, _20848_, _06509_);
  and _72570_ (_20924_, _20922_, _20921_);
  or _72571_ (_20925_, _20924_, _06602_);
  or _72572_ (_20926_, _20925_, _20920_);
  or _72573_ (_20927_, _20905_, _09112_);
  and _72574_ (_20928_, _20927_, _07048_);
  and _72575_ (_20929_, _20928_, _20926_);
  and _72576_ (_20930_, _20855_, _06639_);
  or _72577_ (_20931_, _20930_, _06646_);
  or _72578_ (_20932_, _20931_, _20929_);
  nor _72579_ (_20933_, _20858_, _06651_);
  nand _72580_ (_20935_, _20933_, _20854_);
  and _72581_ (_20936_, _20935_, _01442_);
  and _72582_ (_20937_, _20936_, _20932_);
  or _72583_ (_20938_, _20937_, _20845_);
  and _72584_ (_44150_, _20938_, _43634_);
  and _72585_ (_20939_, _01446_, \oc8051_golden_model_1.DPL [2]);
  and _72586_ (_20940_, _11585_, \oc8051_golden_model_1.DPL [2]);
  nor _72587_ (_20941_, _11585_, _07854_);
  or _72588_ (_20942_, _20941_, _20940_);
  or _72589_ (_20943_, _20942_, _06327_);
  nor _72590_ (_20945_, _11608_, \oc8051_golden_model_1.DPL [2]);
  nor _72591_ (_20946_, _20945_, _11609_);
  and _72592_ (_20947_, _20946_, _11603_);
  or _72593_ (_20948_, _20942_, _06772_);
  and _72594_ (_20949_, _14959_, _08001_);
  or _72595_ (_20950_, _20949_, _20940_);
  and _72596_ (_20951_, _20950_, _06474_);
  and _72597_ (_20952_, _07260_, \oc8051_golden_model_1.DPL [2]);
  and _72598_ (_20953_, _08158_, \oc8051_golden_model_1.ACC [2]);
  or _72599_ (_20954_, _20953_, _20940_);
  and _72600_ (_20956_, _20954_, _07259_);
  or _72601_ (_20957_, _20956_, _20952_);
  and _72602_ (_20958_, _20957_, _07275_);
  or _72603_ (_20959_, _20958_, _06410_);
  or _72604_ (_20960_, _20959_, _20951_);
  and _72605_ (_20961_, _20960_, _20948_);
  or _72606_ (_20962_, _20961_, _06417_);
  or _72607_ (_20963_, _20954_, _06426_);
  and _72608_ (_20964_, _20963_, _11604_);
  and _72609_ (_20965_, _20964_, _20962_);
  or _72610_ (_20967_, _20965_, _20947_);
  and _72611_ (_20968_, _20967_, _06487_);
  nor _72612_ (_20969_, _06769_, _06487_);
  or _72613_ (_20970_, _20969_, _10153_);
  or _72614_ (_20971_, _20970_, _20968_);
  and _72615_ (_20972_, _20971_, _20943_);
  or _72616_ (_20973_, _20972_, _09572_);
  and _72617_ (_20974_, _09356_, _08158_);
  or _72618_ (_20975_, _20940_, _06333_);
  or _72619_ (_20976_, _20975_, _20974_);
  and _72620_ (_20978_, _20976_, _06313_);
  and _72621_ (_20979_, _20978_, _20973_);
  and _72622_ (_20980_, _15056_, _08158_);
  or _72623_ (_20981_, _20980_, _20940_);
  and _72624_ (_20982_, _20981_, _06037_);
  or _72625_ (_20983_, _20982_, _06277_);
  or _72626_ (_20984_, _20983_, _20979_);
  and _72627_ (_20985_, _08158_, _09057_);
  or _72628_ (_20986_, _20985_, _20940_);
  or _72629_ (_20987_, _20986_, _06278_);
  and _72630_ (_20989_, _20987_, _20984_);
  or _72631_ (_20990_, _20989_, _06502_);
  and _72632_ (_20991_, _14948_, _08001_);
  or _72633_ (_20992_, _20940_, _07334_);
  or _72634_ (_20993_, _20992_, _20991_);
  and _72635_ (_20994_, _20993_, _07337_);
  and _72636_ (_20995_, _20994_, _20990_);
  and _72637_ (_20996_, _10583_, _08158_);
  or _72638_ (_20997_, _20996_, _20940_);
  and _72639_ (_20998_, _20997_, _06615_);
  or _72640_ (_21000_, _20998_, _20995_);
  and _72641_ (_21001_, _21000_, _07339_);
  or _72642_ (_21002_, _20940_, _08503_);
  and _72643_ (_21003_, _20986_, _06507_);
  and _72644_ (_21004_, _21003_, _21002_);
  or _72645_ (_21005_, _21004_, _21001_);
  and _72646_ (_21006_, _21005_, _07331_);
  and _72647_ (_21007_, _20954_, _06610_);
  and _72648_ (_21008_, _21007_, _21002_);
  or _72649_ (_21009_, _21008_, _06509_);
  or _72650_ (_21011_, _21009_, _21006_);
  and _72651_ (_21012_, _14945_, _08001_);
  or _72652_ (_21013_, _20940_, _09107_);
  or _72653_ (_21014_, _21013_, _21012_);
  and _72654_ (_21015_, _21014_, _09112_);
  and _72655_ (_21016_, _21015_, _21011_);
  nor _72656_ (_21017_, _10582_, _11585_);
  or _72657_ (_21018_, _21017_, _20940_);
  and _72658_ (_21019_, _21018_, _06602_);
  or _72659_ (_21020_, _21019_, _21016_);
  and _72660_ (_21022_, _21020_, _07048_);
  and _72661_ (_21023_, _20950_, _06639_);
  or _72662_ (_21024_, _21023_, _06646_);
  or _72663_ (_21025_, _21024_, _21022_);
  and _72664_ (_21026_, _15129_, _08001_);
  or _72665_ (_21027_, _20940_, _06651_);
  or _72666_ (_21028_, _21027_, _21026_);
  and _72667_ (_21029_, _21028_, _01442_);
  and _72668_ (_21030_, _21029_, _21025_);
  or _72669_ (_21031_, _21030_, _20939_);
  and _72670_ (_44151_, _21031_, _43634_);
  and _72671_ (_21033_, _11585_, \oc8051_golden_model_1.DPL [3]);
  nor _72672_ (_21034_, _11585_, _07680_);
  or _72673_ (_21035_, _21034_, _21033_);
  or _72674_ (_21036_, _21035_, _06327_);
  and _72675_ (_21037_, _15153_, _08001_);
  or _72676_ (_21038_, _21037_, _21033_);
  or _72677_ (_21039_, _21038_, _07275_);
  and _72678_ (_21040_, _08158_, \oc8051_golden_model_1.ACC [3]);
  or _72679_ (_21041_, _21040_, _21033_);
  and _72680_ (_21043_, _21041_, _07259_);
  and _72681_ (_21044_, _07260_, \oc8051_golden_model_1.DPL [3]);
  or _72682_ (_21045_, _21044_, _06474_);
  or _72683_ (_21046_, _21045_, _21043_);
  and _72684_ (_21047_, _21046_, _06772_);
  and _72685_ (_21048_, _21047_, _21039_);
  and _72686_ (_21049_, _21035_, _06410_);
  or _72687_ (_21050_, _21049_, _06417_);
  or _72688_ (_21051_, _21050_, _21048_);
  or _72689_ (_21052_, _21041_, _06426_);
  and _72690_ (_21054_, _21052_, _11604_);
  and _72691_ (_21055_, _21054_, _21051_);
  nor _72692_ (_21056_, _11609_, \oc8051_golden_model_1.DPL [3]);
  nor _72693_ (_21057_, _21056_, _11610_);
  and _72694_ (_21058_, _21057_, _11603_);
  or _72695_ (_21059_, _21058_, _21055_);
  and _72696_ (_21060_, _21059_, _06487_);
  nor _72697_ (_21061_, _06595_, _06487_);
  or _72698_ (_21062_, _21061_, _10153_);
  or _72699_ (_21063_, _21062_, _21060_);
  and _72700_ (_21064_, _21063_, _21036_);
  or _72701_ (_21065_, _21064_, _09572_);
  and _72702_ (_21066_, _09310_, _08158_);
  or _72703_ (_21067_, _21033_, _06333_);
  or _72704_ (_21068_, _21067_, _21066_);
  and _72705_ (_21069_, _21068_, _06313_);
  and _72706_ (_21070_, _21069_, _21065_);
  and _72707_ (_21071_, _15251_, _08158_);
  or _72708_ (_21072_, _21071_, _21033_);
  and _72709_ (_21073_, _21072_, _06037_);
  or _72710_ (_21076_, _21073_, _06277_);
  or _72711_ (_21077_, _21076_, _21070_);
  and _72712_ (_21078_, _08158_, _09014_);
  or _72713_ (_21079_, _21078_, _21033_);
  or _72714_ (_21080_, _21079_, _06278_);
  and _72715_ (_21081_, _21080_, _21077_);
  or _72716_ (_21082_, _21081_, _06502_);
  and _72717_ (_21083_, _15266_, _08001_);
  or _72718_ (_21084_, _21033_, _07334_);
  or _72719_ (_21085_, _21084_, _21083_);
  and _72720_ (_21087_, _21085_, _07337_);
  and _72721_ (_21088_, _21087_, _21082_);
  and _72722_ (_21089_, _12619_, _08158_);
  or _72723_ (_21090_, _21089_, _21033_);
  and _72724_ (_21091_, _21090_, _06615_);
  or _72725_ (_21092_, _21091_, _21088_);
  and _72726_ (_21093_, _21092_, _07339_);
  or _72727_ (_21094_, _21033_, _08359_);
  and _72728_ (_21095_, _21079_, _06507_);
  and _72729_ (_21096_, _21095_, _21094_);
  or _72730_ (_21098_, _21096_, _21093_);
  and _72731_ (_21099_, _21098_, _07331_);
  and _72732_ (_21100_, _21041_, _06610_);
  and _72733_ (_21101_, _21100_, _21094_);
  or _72734_ (_21102_, _21101_, _06509_);
  or _72735_ (_21103_, _21102_, _21099_);
  and _72736_ (_21104_, _15263_, _08001_);
  or _72737_ (_21105_, _21033_, _09107_);
  or _72738_ (_21106_, _21105_, _21104_);
  and _72739_ (_21107_, _21106_, _09112_);
  and _72740_ (_21109_, _21107_, _21103_);
  nor _72741_ (_21110_, _10574_, _11585_);
  or _72742_ (_21111_, _21110_, _21033_);
  and _72743_ (_21112_, _21111_, _06602_);
  or _72744_ (_21113_, _21112_, _06639_);
  or _72745_ (_21114_, _21113_, _21109_);
  or _72746_ (_21115_, _21038_, _07048_);
  and _72747_ (_21116_, _21115_, _06651_);
  and _72748_ (_21117_, _21116_, _21114_);
  and _72749_ (_21118_, _15321_, _08001_);
  or _72750_ (_21120_, _21118_, _21033_);
  and _72751_ (_21121_, _21120_, _06646_);
  or _72752_ (_21122_, _21121_, _01446_);
  or _72753_ (_21123_, _21122_, _21117_);
  or _72754_ (_21124_, _01442_, \oc8051_golden_model_1.DPL [3]);
  and _72755_ (_21125_, _21124_, _43634_);
  and _72756_ (_44152_, _21125_, _21123_);
  and _72757_ (_21126_, _11585_, \oc8051_golden_model_1.DPL [4]);
  nor _72758_ (_21127_, _08596_, _11585_);
  or _72759_ (_21128_, _21127_, _21126_);
  or _72760_ (_21130_, _21128_, _06327_);
  and _72761_ (_21131_, _15367_, _08001_);
  or _72762_ (_21132_, _21131_, _21126_);
  or _72763_ (_21133_, _21132_, _07275_);
  and _72764_ (_21134_, _08158_, \oc8051_golden_model_1.ACC [4]);
  or _72765_ (_21135_, _21134_, _21126_);
  and _72766_ (_21136_, _21135_, _07259_);
  and _72767_ (_21137_, _07260_, \oc8051_golden_model_1.DPL [4]);
  or _72768_ (_21138_, _21137_, _06474_);
  or _72769_ (_21139_, _21138_, _21136_);
  and _72770_ (_21141_, _21139_, _06772_);
  and _72771_ (_21142_, _21141_, _21133_);
  and _72772_ (_21143_, _21128_, _06410_);
  or _72773_ (_21144_, _21143_, _06417_);
  or _72774_ (_21145_, _21144_, _21142_);
  or _72775_ (_21146_, _21135_, _06426_);
  and _72776_ (_21147_, _21146_, _11604_);
  and _72777_ (_21148_, _21147_, _21145_);
  nor _72778_ (_21149_, _11610_, \oc8051_golden_model_1.DPL [4]);
  nor _72779_ (_21150_, _21149_, _11611_);
  and _72780_ (_21152_, _21150_, _11603_);
  or _72781_ (_21153_, _21152_, _21148_);
  and _72782_ (_21154_, _21153_, _06487_);
  nor _72783_ (_21155_, _08986_, _06487_);
  or _72784_ (_21156_, _21155_, _10153_);
  or _72785_ (_21157_, _21156_, _21154_);
  and _72786_ (_21158_, _21157_, _21130_);
  or _72787_ (_21159_, _21158_, _09572_);
  and _72788_ (_21160_, _09264_, _08158_);
  or _72789_ (_21161_, _21126_, _06333_);
  or _72790_ (_21163_, _21161_, _21160_);
  and _72791_ (_21164_, _21163_, _06313_);
  and _72792_ (_21165_, _21164_, _21159_);
  and _72793_ (_21166_, _15452_, _08158_);
  or _72794_ (_21167_, _21166_, _21126_);
  and _72795_ (_21168_, _21167_, _06037_);
  or _72796_ (_21169_, _21168_, _06277_);
  or _72797_ (_21170_, _21169_, _21165_);
  and _72798_ (_21171_, _08995_, _08158_);
  or _72799_ (_21172_, _21171_, _21126_);
  or _72800_ (_21174_, _21172_, _06278_);
  and _72801_ (_21175_, _21174_, _21170_);
  or _72802_ (_21176_, _21175_, _06502_);
  and _72803_ (_21177_, _15345_, _08001_);
  or _72804_ (_21178_, _21126_, _07334_);
  or _72805_ (_21179_, _21178_, _21177_);
  and _72806_ (_21180_, _21179_, _07337_);
  and _72807_ (_21181_, _21180_, _21176_);
  and _72808_ (_21182_, _10590_, _08158_);
  or _72809_ (_21183_, _21182_, _21126_);
  and _72810_ (_21185_, _21183_, _06615_);
  or _72811_ (_21186_, _21185_, _21181_);
  and _72812_ (_21187_, _21186_, _07339_);
  or _72813_ (_21188_, _21126_, _08599_);
  and _72814_ (_21189_, _21172_, _06507_);
  and _72815_ (_21190_, _21189_, _21188_);
  or _72816_ (_21191_, _21190_, _21187_);
  and _72817_ (_21192_, _21191_, _07331_);
  and _72818_ (_21193_, _21135_, _06610_);
  and _72819_ (_21194_, _21193_, _21188_);
  or _72820_ (_21196_, _21194_, _06509_);
  or _72821_ (_21197_, _21196_, _21192_);
  and _72822_ (_21198_, _15342_, _08001_);
  or _72823_ (_21199_, _21126_, _09107_);
  or _72824_ (_21200_, _21199_, _21198_);
  and _72825_ (_21201_, _21200_, _09112_);
  and _72826_ (_21202_, _21201_, _21197_);
  nor _72827_ (_21203_, _10589_, _11585_);
  or _72828_ (_21204_, _21203_, _21126_);
  and _72829_ (_21205_, _21204_, _06602_);
  or _72830_ (_21207_, _21205_, _06639_);
  or _72831_ (_21208_, _21207_, _21202_);
  or _72832_ (_21209_, _21132_, _07048_);
  and _72833_ (_21210_, _21209_, _06651_);
  and _72834_ (_21211_, _21210_, _21208_);
  and _72835_ (_21212_, _15524_, _08001_);
  or _72836_ (_21213_, _21212_, _21126_);
  and _72837_ (_21214_, _21213_, _06646_);
  or _72838_ (_21215_, _21214_, _01446_);
  or _72839_ (_21216_, _21215_, _21211_);
  or _72840_ (_21218_, _01442_, \oc8051_golden_model_1.DPL [4]);
  and _72841_ (_21219_, _21218_, _43634_);
  and _72842_ (_44153_, _21219_, _21216_);
  and _72843_ (_21220_, _11585_, \oc8051_golden_model_1.DPL [5]);
  nor _72844_ (_21221_, _10570_, _11585_);
  or _72845_ (_21222_, _21221_, _21220_);
  and _72846_ (_21223_, _08158_, \oc8051_golden_model_1.ACC [5]);
  nand _72847_ (_21224_, _21223_, _08308_);
  and _72848_ (_21225_, _21224_, _06615_);
  and _72849_ (_21226_, _21225_, _21222_);
  nor _72850_ (_21228_, _08305_, _11585_);
  or _72851_ (_21229_, _21228_, _21220_);
  or _72852_ (_21230_, _21229_, _06327_);
  and _72853_ (_21231_, _15550_, _08001_);
  or _72854_ (_21232_, _21231_, _21220_);
  or _72855_ (_21233_, _21232_, _07275_);
  or _72856_ (_21234_, _21223_, _21220_);
  and _72857_ (_21235_, _21234_, _07259_);
  and _72858_ (_21236_, _07260_, \oc8051_golden_model_1.DPL [5]);
  or _72859_ (_21237_, _21236_, _06474_);
  or _72860_ (_21239_, _21237_, _21235_);
  and _72861_ (_21240_, _21239_, _06772_);
  and _72862_ (_21241_, _21240_, _21233_);
  and _72863_ (_21242_, _21229_, _06410_);
  or _72864_ (_21243_, _21242_, _06417_);
  or _72865_ (_21244_, _21243_, _21241_);
  or _72866_ (_21245_, _21234_, _06426_);
  and _72867_ (_21246_, _21245_, _11604_);
  and _72868_ (_21247_, _21246_, _21244_);
  nor _72869_ (_21248_, _11611_, \oc8051_golden_model_1.DPL [5]);
  nor _72870_ (_21250_, _21248_, _11612_);
  and _72871_ (_21251_, _21250_, _11603_);
  or _72872_ (_21252_, _21251_, _21247_);
  and _72873_ (_21253_, _21252_, _06487_);
  nor _72874_ (_21254_, _08953_, _06487_);
  or _72875_ (_21255_, _21254_, _10153_);
  or _72876_ (_21256_, _21255_, _21253_);
  and _72877_ (_21257_, _21256_, _21230_);
  or _72878_ (_21258_, _21257_, _09572_);
  and _72879_ (_21259_, _09218_, _08158_);
  or _72880_ (_21260_, _21220_, _06333_);
  or _72881_ (_21261_, _21260_, _21259_);
  and _72882_ (_21262_, _21261_, _06313_);
  and _72883_ (_21263_, _21262_, _21258_);
  and _72884_ (_21264_, _15649_, _08158_);
  or _72885_ (_21265_, _21264_, _21220_);
  and _72886_ (_21266_, _21265_, _06037_);
  or _72887_ (_21267_, _21266_, _06277_);
  or _72888_ (_21268_, _21267_, _21263_);
  and _72889_ (_21269_, _08954_, _08158_);
  or _72890_ (_21272_, _21269_, _21220_);
  or _72891_ (_21273_, _21272_, _06278_);
  and _72892_ (_21274_, _21273_, _21268_);
  or _72893_ (_21275_, _21274_, _06502_);
  and _72894_ (_21276_, _15664_, _08001_);
  or _72895_ (_21277_, _21220_, _07334_);
  or _72896_ (_21278_, _21277_, _21276_);
  and _72897_ (_21279_, _21278_, _07337_);
  and _72898_ (_21280_, _21279_, _21275_);
  or _72899_ (_21281_, _21280_, _21226_);
  and _72900_ (_21283_, _21281_, _07339_);
  or _72901_ (_21284_, _21220_, _08308_);
  and _72902_ (_21285_, _21272_, _06507_);
  and _72903_ (_21286_, _21285_, _21284_);
  or _72904_ (_21287_, _21286_, _21283_);
  and _72905_ (_21288_, _21287_, _07331_);
  and _72906_ (_21289_, _21234_, _06610_);
  and _72907_ (_21290_, _21289_, _21284_);
  or _72908_ (_21291_, _21290_, _06509_);
  or _72909_ (_21292_, _21291_, _21288_);
  and _72910_ (_21294_, _15663_, _08001_);
  or _72911_ (_21295_, _21220_, _09107_);
  or _72912_ (_21296_, _21295_, _21294_);
  and _72913_ (_21297_, _21296_, _09112_);
  and _72914_ (_21298_, _21297_, _21292_);
  and _72915_ (_21299_, _21222_, _06602_);
  or _72916_ (_21300_, _21299_, _06639_);
  or _72917_ (_21301_, _21300_, _21298_);
  or _72918_ (_21302_, _21232_, _07048_);
  and _72919_ (_21303_, _21302_, _06651_);
  and _72920_ (_21305_, _21303_, _21301_);
  and _72921_ (_21306_, _15721_, _08001_);
  or _72922_ (_21307_, _21306_, _21220_);
  and _72923_ (_21308_, _21307_, _06646_);
  or _72924_ (_21309_, _21308_, _01446_);
  or _72925_ (_21310_, _21309_, _21305_);
  or _72926_ (_21311_, _01442_, \oc8051_golden_model_1.DPL [5]);
  and _72927_ (_21312_, _21311_, _43634_);
  and _72928_ (_44154_, _21312_, _21310_);
  and _72929_ (_21313_, _11585_, \oc8051_golden_model_1.DPL [6]);
  nor _72930_ (_21315_, _10595_, _11585_);
  or _72931_ (_21316_, _21315_, _21313_);
  and _72932_ (_21317_, _08158_, \oc8051_golden_model_1.ACC [6]);
  nand _72933_ (_21318_, _21317_, _08212_);
  and _72934_ (_21319_, _21318_, _06615_);
  and _72935_ (_21320_, _21319_, _21316_);
  nor _72936_ (_21321_, _08209_, _11585_);
  or _72937_ (_21322_, _21321_, _21313_);
  or _72938_ (_21323_, _21322_, _06327_);
  and _72939_ (_21324_, _15759_, _08001_);
  or _72940_ (_21326_, _21324_, _21313_);
  or _72941_ (_21327_, _21326_, _07275_);
  or _72942_ (_21328_, _21317_, _21313_);
  and _72943_ (_21329_, _21328_, _07259_);
  and _72944_ (_21330_, _07260_, \oc8051_golden_model_1.DPL [6]);
  or _72945_ (_21331_, _21330_, _06474_);
  or _72946_ (_21332_, _21331_, _21329_);
  and _72947_ (_21333_, _21332_, _06772_);
  and _72948_ (_21334_, _21333_, _21327_);
  and _72949_ (_21335_, _21322_, _06410_);
  or _72950_ (_21337_, _21335_, _06417_);
  or _72951_ (_21338_, _21337_, _21334_);
  or _72952_ (_21339_, _21328_, _06426_);
  and _72953_ (_21340_, _21339_, _11604_);
  and _72954_ (_21341_, _21340_, _21338_);
  nor _72955_ (_21342_, _11612_, \oc8051_golden_model_1.DPL [6]);
  nor _72956_ (_21343_, _21342_, _11613_);
  and _72957_ (_21344_, _21343_, _11603_);
  or _72958_ (_21345_, _21344_, _21341_);
  and _72959_ (_21346_, _21345_, _06487_);
  nor _72960_ (_21348_, _08918_, _06487_);
  or _72961_ (_21349_, _21348_, _10153_);
  or _72962_ (_21350_, _21349_, _21346_);
  and _72963_ (_21351_, _21350_, _21323_);
  or _72964_ (_21352_, _21351_, _09572_);
  and _72965_ (_21353_, _09172_, _08158_);
  or _72966_ (_21354_, _21313_, _06333_);
  or _72967_ (_21355_, _21354_, _21353_);
  and _72968_ (_21356_, _21355_, _06313_);
  and _72969_ (_21357_, _21356_, _21352_);
  and _72970_ (_21359_, _15846_, _08158_);
  or _72971_ (_21360_, _21359_, _21313_);
  and _72972_ (_21361_, _21360_, _06037_);
  or _72973_ (_21362_, _21361_, _06277_);
  or _72974_ (_21363_, _21362_, _21357_);
  and _72975_ (_21364_, _15853_, _08158_);
  or _72976_ (_21365_, _21364_, _21313_);
  or _72977_ (_21366_, _21365_, _06278_);
  and _72978_ (_21367_, _21366_, _21363_);
  or _72979_ (_21368_, _21367_, _06502_);
  and _72980_ (_21370_, _15862_, _08001_);
  or _72981_ (_21371_, _21313_, _07334_);
  or _72982_ (_21372_, _21371_, _21370_);
  and _72983_ (_21373_, _21372_, _07337_);
  and _72984_ (_21374_, _21373_, _21368_);
  or _72985_ (_21375_, _21374_, _21320_);
  and _72986_ (_21376_, _21375_, _07339_);
  or _72987_ (_21377_, _21313_, _08212_);
  and _72988_ (_21378_, _21365_, _06507_);
  and _72989_ (_21379_, _21378_, _21377_);
  or _72990_ (_21381_, _21379_, _21376_);
  and _72991_ (_21382_, _21381_, _07331_);
  and _72992_ (_21383_, _21328_, _06610_);
  and _72993_ (_21384_, _21383_, _21377_);
  or _72994_ (_21385_, _21384_, _06509_);
  or _72995_ (_21386_, _21385_, _21382_);
  and _72996_ (_21387_, _15859_, _08001_);
  or _72997_ (_21388_, _21313_, _09107_);
  or _72998_ (_21389_, _21388_, _21387_);
  and _72999_ (_21390_, _21389_, _09112_);
  and _73000_ (_21392_, _21390_, _21386_);
  and _73001_ (_21393_, _21316_, _06602_);
  or _73002_ (_21394_, _21393_, _06639_);
  or _73003_ (_21395_, _21394_, _21392_);
  or _73004_ (_21396_, _21326_, _07048_);
  and _73005_ (_21397_, _21396_, _06651_);
  and _73006_ (_21398_, _21397_, _21395_);
  and _73007_ (_21399_, _15921_, _08001_);
  or _73008_ (_21400_, _21399_, _21313_);
  and _73009_ (_21401_, _21400_, _06646_);
  or _73010_ (_21403_, _21401_, _01446_);
  or _73011_ (_21404_, _21403_, _21398_);
  or _73012_ (_21405_, _01442_, \oc8051_golden_model_1.DPL [6]);
  and _73013_ (_21406_, _21405_, _43634_);
  and _73014_ (_44155_, _21406_, _21404_);
  nor _73015_ (_21407_, _01442_, _12726_);
  nor _73016_ (_21408_, _08153_, _12726_);
  nor _73017_ (_21409_, _12622_, _11681_);
  or _73018_ (_21410_, _21409_, _21408_);
  and _73019_ (_21411_, _08153_, \oc8051_golden_model_1.ACC [0]);
  and _73020_ (_21413_, _21411_, _08453_);
  nor _73021_ (_21414_, _21413_, _07337_);
  and _73022_ (_21415_, _21414_, _21410_);
  and _73023_ (_21416_, _09447_, _08153_);
  or _73024_ (_21417_, _21416_, _21408_);
  and _73025_ (_21418_, _21417_, _14025_);
  and _73026_ (_21419_, _07995_, _07250_);
  or _73027_ (_21420_, _21419_, _21408_);
  or _73028_ (_21421_, _21420_, _06772_);
  nor _73029_ (_21422_, _08453_, _11681_);
  or _73030_ (_21424_, _21422_, _21408_);
  and _73031_ (_21425_, _21424_, _06474_);
  nor _73032_ (_21426_, _07259_, _12726_);
  or _73033_ (_21427_, _21411_, _21408_);
  and _73034_ (_21428_, _21427_, _07259_);
  or _73035_ (_21429_, _21428_, _21426_);
  and _73036_ (_21430_, _21429_, _07275_);
  or _73037_ (_21431_, _21430_, _06410_);
  or _73038_ (_21432_, _21431_, _21425_);
  and _73039_ (_21433_, _21432_, _21421_);
  or _73040_ (_21435_, _21433_, _06417_);
  or _73041_ (_21436_, _21427_, _06426_);
  and _73042_ (_21437_, _21436_, _11604_);
  and _73043_ (_21438_, _21437_, _21435_);
  nor _73044_ (_21439_, _11615_, \oc8051_golden_model_1.DPH [0]);
  nor _73045_ (_21440_, _21439_, _11702_);
  and _73046_ (_21441_, _21440_, _11603_);
  or _73047_ (_21442_, _21441_, _21438_);
  and _73048_ (_21443_, _21442_, _06487_);
  nor _73049_ (_21444_, _06487_, _06310_);
  or _73050_ (_21446_, _21444_, _10153_);
  or _73051_ (_21447_, _21446_, _21443_);
  or _73052_ (_21448_, _21420_, _06327_);
  and _73053_ (_21449_, _21448_, _16672_);
  and _73054_ (_21450_, _21449_, _21447_);
  or _73055_ (_21451_, _21450_, _06037_);
  or _73056_ (_21452_, _21451_, _21418_);
  and _73057_ (_21453_, _14666_, _07995_);
  or _73058_ (_21454_, _21408_, _06313_);
  or _73059_ (_21455_, _21454_, _21453_);
  and _73060_ (_21457_, _21455_, _06278_);
  and _73061_ (_21458_, _21457_, _21452_);
  and _73062_ (_21459_, _08153_, _09008_);
  or _73063_ (_21460_, _21459_, _21408_);
  and _73064_ (_21461_, _21460_, _06277_);
  or _73065_ (_21462_, _21461_, _06502_);
  or _73066_ (_21463_, _21462_, _21458_);
  and _73067_ (_21464_, _14566_, _07995_);
  or _73068_ (_21465_, _21408_, _07334_);
  or _73069_ (_21466_, _21465_, _21464_);
  and _73070_ (_21468_, _21466_, _07337_);
  and _73071_ (_21469_, _21468_, _21463_);
  or _73072_ (_21470_, _21469_, _21415_);
  and _73073_ (_21471_, _21470_, _07339_);
  nand _73074_ (_21472_, _21460_, _06507_);
  nor _73075_ (_21473_, _21472_, _21422_);
  or _73076_ (_21474_, _21473_, _06610_);
  or _73077_ (_21475_, _21474_, _21471_);
  or _73078_ (_21476_, _21413_, _21408_);
  or _73079_ (_21477_, _21476_, _07331_);
  and _73080_ (_21479_, _21477_, _21475_);
  or _73081_ (_21480_, _21479_, _06509_);
  and _73082_ (_21481_, _14563_, _07995_);
  or _73083_ (_21482_, _21408_, _09107_);
  or _73084_ (_21483_, _21482_, _21481_);
  and _73085_ (_21484_, _21483_, _09112_);
  and _73086_ (_21485_, _21484_, _21480_);
  and _73087_ (_21486_, _21410_, _06602_);
  or _73088_ (_21487_, _21486_, _19642_);
  or _73089_ (_21488_, _21487_, _21485_);
  or _73090_ (_21490_, _21424_, _19641_);
  and _73091_ (_21491_, _21490_, _01442_);
  and _73092_ (_21492_, _21491_, _21488_);
  or _73093_ (_21493_, _21492_, _21407_);
  and _73094_ (_44157_, _21493_, _43634_);
  not _73095_ (_21494_, \oc8051_golden_model_1.DPH [1]);
  nor _73096_ (_21495_, _08153_, _21494_);
  nor _73097_ (_21496_, _10578_, _11681_);
  or _73098_ (_21497_, _21496_, _21495_);
  or _73099_ (_21498_, _21497_, _09112_);
  or _73100_ (_21500_, _08153_, \oc8051_golden_model_1.DPH [1]);
  and _73101_ (_21501_, _21500_, _06277_);
  nand _73102_ (_21502_, _07995_, _07160_);
  and _73103_ (_21503_, _21502_, _21501_);
  or _73104_ (_21504_, _09402_, _11681_);
  and _73105_ (_21505_, _21500_, _14025_);
  and _73106_ (_21506_, _21505_, _21504_);
  nor _73107_ (_21507_, _11702_, \oc8051_golden_model_1.DPH [1]);
  nor _73108_ (_21508_, _21507_, _11703_);
  and _73109_ (_21509_, _21508_, _11603_);
  and _73110_ (_21511_, _14744_, _07995_);
  not _73111_ (_21512_, _21511_);
  and _73112_ (_21513_, _21512_, _21500_);
  or _73113_ (_21514_, _21513_, _07275_);
  and _73114_ (_21515_, _08153_, \oc8051_golden_model_1.ACC [1]);
  or _73115_ (_21516_, _21515_, _21495_);
  and _73116_ (_21517_, _21516_, _07259_);
  nor _73117_ (_21518_, _07259_, _21494_);
  or _73118_ (_21519_, _21518_, _06474_);
  or _73119_ (_21520_, _21519_, _21517_);
  and _73120_ (_21522_, _21520_, _06772_);
  and _73121_ (_21523_, _21522_, _21514_);
  nor _73122_ (_21524_, _11681_, _07448_);
  or _73123_ (_21525_, _21524_, _21495_);
  and _73124_ (_21526_, _21525_, _06410_);
  or _73125_ (_21527_, _21526_, _06417_);
  or _73126_ (_21528_, _21527_, _21523_);
  or _73127_ (_21529_, _21516_, _06426_);
  and _73128_ (_21530_, _21529_, _11604_);
  and _73129_ (_21531_, _21530_, _21528_);
  or _73130_ (_21533_, _21531_, _21509_);
  and _73131_ (_21534_, _21533_, _06487_);
  nor _73132_ (_21535_, _07127_, _06487_);
  or _73133_ (_21536_, _21535_, _10153_);
  or _73134_ (_21537_, _21536_, _21534_);
  or _73135_ (_21538_, _21525_, _06327_);
  and _73136_ (_21539_, _21538_, _16672_);
  and _73137_ (_21540_, _21539_, _21537_);
  or _73138_ (_21541_, _21540_, _21506_);
  and _73139_ (_21542_, _21541_, _06313_);
  and _73140_ (_21544_, _14851_, _08153_);
  or _73141_ (_21545_, _21544_, _21495_);
  and _73142_ (_21546_, _21545_, _06037_);
  or _73143_ (_21547_, _21546_, _21542_);
  and _73144_ (_21548_, _21547_, _06278_);
  or _73145_ (_21549_, _21548_, _21503_);
  and _73146_ (_21550_, _21549_, _07334_);
  or _73147_ (_21551_, _14749_, _11681_);
  and _73148_ (_21552_, _21500_, _06502_);
  and _73149_ (_21553_, _21552_, _21551_);
  or _73150_ (_21555_, _21553_, _06615_);
  or _73151_ (_21556_, _21555_, _21550_);
  nand _73152_ (_21557_, _10576_, _07995_);
  and _73153_ (_21558_, _21557_, _21497_);
  or _73154_ (_21559_, _21558_, _07337_);
  and _73155_ (_21560_, _21559_, _07339_);
  and _73156_ (_21561_, _21560_, _21556_);
  or _73157_ (_21562_, _14747_, _11681_);
  and _73158_ (_21563_, _21500_, _06507_);
  and _73159_ (_21564_, _21563_, _21562_);
  or _73160_ (_21566_, _21564_, _06610_);
  or _73161_ (_21567_, _21566_, _21561_);
  nor _73162_ (_21568_, _21495_, _07331_);
  nand _73163_ (_21569_, _21568_, _21557_);
  and _73164_ (_21570_, _21569_, _09107_);
  and _73165_ (_21571_, _21570_, _21567_);
  or _73166_ (_21572_, _21502_, _08404_);
  and _73167_ (_21573_, _21500_, _06509_);
  and _73168_ (_21574_, _21573_, _21572_);
  or _73169_ (_21575_, _21574_, _06602_);
  or _73170_ (_21577_, _21575_, _21571_);
  and _73171_ (_21578_, _21577_, _21498_);
  or _73172_ (_21579_, _21578_, _06639_);
  or _73173_ (_21580_, _21513_, _07048_);
  and _73174_ (_21581_, _21580_, _06651_);
  and _73175_ (_21582_, _21581_, _21579_);
  or _73176_ (_21583_, _21511_, _21495_);
  and _73177_ (_21584_, _21583_, _06646_);
  or _73178_ (_21585_, _21584_, _01446_);
  or _73179_ (_21586_, _21585_, _21582_);
  or _73180_ (_21588_, _01442_, \oc8051_golden_model_1.DPH [1]);
  and _73181_ (_21589_, _21588_, _43634_);
  and _73182_ (_44158_, _21589_, _21586_);
  and _73183_ (_21590_, _01446_, \oc8051_golden_model_1.DPH [2]);
  and _73184_ (_21591_, _11681_, \oc8051_golden_model_1.DPH [2]);
  nor _73185_ (_21592_, _11681_, _07854_);
  or _73186_ (_21593_, _21592_, _21591_);
  or _73187_ (_21594_, _21593_, _06327_);
  or _73188_ (_21595_, _11703_, \oc8051_golden_model_1.DPH [2]);
  nor _73189_ (_21596_, _11704_, _11604_);
  and _73190_ (_21598_, _21596_, _21595_);
  and _73191_ (_21599_, _14959_, _07995_);
  or _73192_ (_21600_, _21599_, _21591_);
  or _73193_ (_21601_, _21600_, _07275_);
  and _73194_ (_21602_, _08153_, \oc8051_golden_model_1.ACC [2]);
  or _73195_ (_21603_, _21602_, _21591_);
  and _73196_ (_21604_, _21603_, _07259_);
  and _73197_ (_21605_, _07260_, \oc8051_golden_model_1.DPH [2]);
  or _73198_ (_21606_, _21605_, _06474_);
  or _73199_ (_21607_, _21606_, _21604_);
  and _73200_ (_21608_, _21607_, _06772_);
  and _73201_ (_21609_, _21608_, _21601_);
  and _73202_ (_21610_, _21593_, _06410_);
  or _73203_ (_21611_, _21610_, _06417_);
  or _73204_ (_21612_, _21611_, _21609_);
  or _73205_ (_21613_, _21603_, _06426_);
  and _73206_ (_21614_, _21613_, _11604_);
  and _73207_ (_21615_, _21614_, _21612_);
  or _73208_ (_21616_, _21615_, _21598_);
  and _73209_ (_21617_, _21616_, _06487_);
  nor _73210_ (_21620_, _06727_, _06487_);
  or _73211_ (_21621_, _21620_, _10153_);
  or _73212_ (_21622_, _21621_, _21617_);
  and _73213_ (_21623_, _21622_, _21594_);
  or _73214_ (_21624_, _21623_, _09572_);
  and _73215_ (_21625_, _09356_, _08153_);
  or _73216_ (_21626_, _21591_, _06333_);
  or _73217_ (_21627_, _21626_, _21625_);
  and _73218_ (_21628_, _21627_, _06313_);
  and _73219_ (_21629_, _21628_, _21624_);
  and _73220_ (_21631_, _15056_, _08153_);
  or _73221_ (_21632_, _21631_, _21591_);
  and _73222_ (_21633_, _21632_, _06037_);
  or _73223_ (_21634_, _21633_, _06277_);
  or _73224_ (_21635_, _21634_, _21629_);
  and _73225_ (_21636_, _08153_, _09057_);
  or _73226_ (_21637_, _21636_, _21591_);
  or _73227_ (_21638_, _21637_, _06278_);
  and _73228_ (_21639_, _21638_, _21635_);
  or _73229_ (_21640_, _21639_, _06502_);
  and _73230_ (_21642_, _14948_, _07995_);
  or _73231_ (_21643_, _21591_, _07334_);
  or _73232_ (_21644_, _21643_, _21642_);
  and _73233_ (_21645_, _21644_, _07337_);
  and _73234_ (_21646_, _21645_, _21640_);
  and _73235_ (_21647_, _10583_, _08153_);
  or _73236_ (_21648_, _21647_, _21591_);
  and _73237_ (_21649_, _21648_, _06615_);
  or _73238_ (_21650_, _21649_, _21646_);
  and _73239_ (_21651_, _21650_, _07339_);
  or _73240_ (_21653_, _21591_, _08503_);
  and _73241_ (_21654_, _21637_, _06507_);
  and _73242_ (_21655_, _21654_, _21653_);
  or _73243_ (_21656_, _21655_, _21651_);
  and _73244_ (_21657_, _21656_, _07331_);
  and _73245_ (_21658_, _21603_, _06610_);
  and _73246_ (_21659_, _21658_, _21653_);
  or _73247_ (_21660_, _21659_, _06509_);
  or _73248_ (_21661_, _21660_, _21657_);
  and _73249_ (_21662_, _14945_, _07995_);
  or _73250_ (_21664_, _21591_, _09107_);
  or _73251_ (_21665_, _21664_, _21662_);
  and _73252_ (_21666_, _21665_, _09112_);
  and _73253_ (_21667_, _21666_, _21661_);
  nor _73254_ (_21668_, _10582_, _11681_);
  or _73255_ (_21669_, _21668_, _21591_);
  and _73256_ (_21670_, _21669_, _06602_);
  or _73257_ (_21671_, _21670_, _21667_);
  and _73258_ (_21672_, _21671_, _07048_);
  and _73259_ (_21673_, _21600_, _06639_);
  or _73260_ (_21675_, _21673_, _06646_);
  or _73261_ (_21676_, _21675_, _21672_);
  and _73262_ (_21677_, _15129_, _07995_);
  or _73263_ (_21678_, _21591_, _06651_);
  or _73264_ (_21679_, _21678_, _21677_);
  and _73265_ (_21680_, _21679_, _01442_);
  and _73266_ (_21681_, _21680_, _21676_);
  or _73267_ (_21682_, _21681_, _21590_);
  and _73268_ (_44159_, _21682_, _43634_);
  and _73269_ (_21683_, _11681_, \oc8051_golden_model_1.DPH [3]);
  nor _73270_ (_21685_, _11681_, _07680_);
  or _73271_ (_21686_, _21685_, _21683_);
  or _73272_ (_21687_, _21686_, _06327_);
  and _73273_ (_21688_, _15153_, _07995_);
  or _73274_ (_21689_, _21688_, _21683_);
  or _73275_ (_21690_, _21689_, _07275_);
  and _73276_ (_21691_, _08153_, \oc8051_golden_model_1.ACC [3]);
  or _73277_ (_21692_, _21691_, _21683_);
  and _73278_ (_21693_, _21692_, _07259_);
  and _73279_ (_21694_, _07260_, \oc8051_golden_model_1.DPH [3]);
  or _73280_ (_21696_, _21694_, _06474_);
  or _73281_ (_21697_, _21696_, _21693_);
  and _73282_ (_21698_, _21697_, _06772_);
  and _73283_ (_21699_, _21698_, _21690_);
  and _73284_ (_21700_, _21686_, _06410_);
  or _73285_ (_21701_, _21700_, _06417_);
  or _73286_ (_21702_, _21701_, _21699_);
  or _73287_ (_21703_, _21692_, _06426_);
  and _73288_ (_21704_, _21703_, _11604_);
  and _73289_ (_21705_, _21704_, _21702_);
  or _73290_ (_21707_, _11704_, \oc8051_golden_model_1.DPH [3]);
  nor _73291_ (_21708_, _11705_, _11604_);
  and _73292_ (_21709_, _21708_, _21707_);
  or _73293_ (_21710_, _21709_, _21705_);
  and _73294_ (_21711_, _21710_, _06487_);
  nor _73295_ (_21712_, _06487_, _06269_);
  or _73296_ (_21713_, _21712_, _10153_);
  or _73297_ (_21714_, _21713_, _21711_);
  and _73298_ (_21715_, _21714_, _21687_);
  or _73299_ (_21716_, _21715_, _09572_);
  and _73300_ (_21717_, _09310_, _08153_);
  or _73301_ (_21718_, _21683_, _06333_);
  or _73302_ (_21719_, _21718_, _21717_);
  and _73303_ (_21720_, _21719_, _06313_);
  and _73304_ (_21721_, _21720_, _21716_);
  and _73305_ (_21722_, _15251_, _08153_);
  or _73306_ (_21723_, _21722_, _21683_);
  and _73307_ (_21724_, _21723_, _06037_);
  or _73308_ (_21725_, _21724_, _06277_);
  or _73309_ (_21726_, _21725_, _21721_);
  and _73310_ (_21729_, _08153_, _09014_);
  or _73311_ (_21730_, _21729_, _21683_);
  or _73312_ (_21731_, _21730_, _06278_);
  and _73313_ (_21732_, _21731_, _21726_);
  or _73314_ (_21733_, _21732_, _06502_);
  and _73315_ (_21734_, _15266_, _07995_);
  or _73316_ (_21735_, _21683_, _07334_);
  or _73317_ (_21736_, _21735_, _21734_);
  and _73318_ (_21737_, _21736_, _07337_);
  and _73319_ (_21738_, _21737_, _21733_);
  and _73320_ (_21740_, _12619_, _08153_);
  or _73321_ (_21741_, _21740_, _21683_);
  and _73322_ (_21742_, _21741_, _06615_);
  or _73323_ (_21743_, _21742_, _21738_);
  and _73324_ (_21744_, _21743_, _07339_);
  or _73325_ (_21745_, _21683_, _08359_);
  and _73326_ (_21746_, _21730_, _06507_);
  and _73327_ (_21747_, _21746_, _21745_);
  or _73328_ (_21748_, _21747_, _21744_);
  and _73329_ (_21749_, _21748_, _07331_);
  and _73330_ (_21751_, _21692_, _06610_);
  and _73331_ (_21752_, _21751_, _21745_);
  or _73332_ (_21753_, _21752_, _06509_);
  or _73333_ (_21754_, _21753_, _21749_);
  and _73334_ (_21755_, _15263_, _07995_);
  or _73335_ (_21756_, _21683_, _09107_);
  or _73336_ (_21757_, _21756_, _21755_);
  and _73337_ (_21758_, _21757_, _09112_);
  and _73338_ (_21759_, _21758_, _21754_);
  nor _73339_ (_21760_, _10574_, _11681_);
  or _73340_ (_21762_, _21760_, _21683_);
  and _73341_ (_21763_, _21762_, _06602_);
  or _73342_ (_21764_, _21763_, _06639_);
  or _73343_ (_21765_, _21764_, _21759_);
  or _73344_ (_21766_, _21689_, _07048_);
  and _73345_ (_21767_, _21766_, _06651_);
  and _73346_ (_21768_, _21767_, _21765_);
  and _73347_ (_21769_, _15321_, _07995_);
  or _73348_ (_21770_, _21769_, _21683_);
  and _73349_ (_21771_, _21770_, _06646_);
  or _73350_ (_21773_, _21771_, _01446_);
  or _73351_ (_21774_, _21773_, _21768_);
  or _73352_ (_21775_, _01442_, \oc8051_golden_model_1.DPH [3]);
  and _73353_ (_21776_, _21775_, _43634_);
  and _73354_ (_44160_, _21776_, _21774_);
  not _73355_ (_21777_, \oc8051_golden_model_1.DPH [4]);
  nor _73356_ (_21778_, _08153_, _21777_);
  nor _73357_ (_21779_, _08596_, _11681_);
  or _73358_ (_21780_, _21779_, _21778_);
  or _73359_ (_21781_, _21780_, _06327_);
  and _73360_ (_21783_, _15367_, _07995_);
  or _73361_ (_21784_, _21783_, _21778_);
  or _73362_ (_21785_, _21784_, _07275_);
  and _73363_ (_21786_, _08153_, \oc8051_golden_model_1.ACC [4]);
  or _73364_ (_21787_, _21786_, _21778_);
  and _73365_ (_21788_, _21787_, _07259_);
  nor _73366_ (_21789_, _07259_, _21777_);
  or _73367_ (_21790_, _21789_, _06474_);
  or _73368_ (_21791_, _21790_, _21788_);
  and _73369_ (_21792_, _21791_, _06772_);
  and _73370_ (_21794_, _21792_, _21785_);
  and _73371_ (_21795_, _21780_, _06410_);
  or _73372_ (_21796_, _21795_, _06417_);
  or _73373_ (_21797_, _21796_, _21794_);
  or _73374_ (_21798_, _21787_, _06426_);
  and _73375_ (_21799_, _21798_, _11604_);
  and _73376_ (_21800_, _21799_, _21797_);
  or _73377_ (_21801_, _11705_, \oc8051_golden_model_1.DPH [4]);
  nor _73378_ (_21802_, _11706_, _11604_);
  and _73379_ (_21803_, _21802_, _21801_);
  or _73380_ (_21805_, _21803_, _21800_);
  and _73381_ (_21806_, _21805_, _06487_);
  nor _73382_ (_21807_, _07093_, _06487_);
  or _73383_ (_21808_, _21807_, _10153_);
  or _73384_ (_21809_, _21808_, _21806_);
  and _73385_ (_21810_, _21809_, _21781_);
  or _73386_ (_21811_, _21810_, _09572_);
  and _73387_ (_21812_, _09264_, _08153_);
  or _73388_ (_21813_, _21778_, _06333_);
  or _73389_ (_21814_, _21813_, _21812_);
  and _73390_ (_21816_, _21814_, _06313_);
  and _73391_ (_21817_, _21816_, _21811_);
  and _73392_ (_21818_, _15452_, _08153_);
  or _73393_ (_21819_, _21818_, _21778_);
  and _73394_ (_21820_, _21819_, _06037_);
  or _73395_ (_21821_, _21820_, _06277_);
  or _73396_ (_21822_, _21821_, _21817_);
  and _73397_ (_21823_, _08995_, _08153_);
  or _73398_ (_21824_, _21823_, _21778_);
  or _73399_ (_21825_, _21824_, _06278_);
  and _73400_ (_21827_, _21825_, _21822_);
  or _73401_ (_21828_, _21827_, _06502_);
  and _73402_ (_21829_, _15345_, _07995_);
  or _73403_ (_21830_, _21778_, _07334_);
  or _73404_ (_21831_, _21830_, _21829_);
  and _73405_ (_21832_, _21831_, _07337_);
  and _73406_ (_21833_, _21832_, _21828_);
  and _73407_ (_21834_, _10590_, _08153_);
  or _73408_ (_21835_, _21834_, _21778_);
  and _73409_ (_21836_, _21835_, _06615_);
  or _73410_ (_21838_, _21836_, _21833_);
  and _73411_ (_21839_, _21838_, _07339_);
  or _73412_ (_21840_, _21778_, _08599_);
  and _73413_ (_21841_, _21824_, _06507_);
  and _73414_ (_21842_, _21841_, _21840_);
  or _73415_ (_21843_, _21842_, _21839_);
  and _73416_ (_21844_, _21843_, _07331_);
  and _73417_ (_21845_, _21787_, _06610_);
  and _73418_ (_21846_, _21845_, _21840_);
  or _73419_ (_21847_, _21846_, _06509_);
  or _73420_ (_21849_, _21847_, _21844_);
  and _73421_ (_21850_, _15342_, _07995_);
  or _73422_ (_21851_, _21778_, _09107_);
  or _73423_ (_21852_, _21851_, _21850_);
  and _73424_ (_21853_, _21852_, _09112_);
  and _73425_ (_21854_, _21853_, _21849_);
  nor _73426_ (_21855_, _10589_, _11681_);
  or _73427_ (_21856_, _21855_, _21778_);
  and _73428_ (_21857_, _21856_, _06602_);
  or _73429_ (_21858_, _21857_, _06639_);
  or _73430_ (_21860_, _21858_, _21854_);
  or _73431_ (_21861_, _21784_, _07048_);
  and _73432_ (_21862_, _21861_, _06651_);
  and _73433_ (_21863_, _21862_, _21860_);
  and _73434_ (_21864_, _15524_, _07995_);
  or _73435_ (_21865_, _21864_, _21778_);
  and _73436_ (_21866_, _21865_, _06646_);
  or _73437_ (_21867_, _21866_, _01446_);
  or _73438_ (_21868_, _21867_, _21863_);
  or _73439_ (_21869_, _01442_, \oc8051_golden_model_1.DPH [4]);
  and _73440_ (_21871_, _21869_, _43634_);
  and _73441_ (_44161_, _21871_, _21868_);
  and _73442_ (_21872_, _11681_, \oc8051_golden_model_1.DPH [5]);
  nor _73443_ (_21873_, _10570_, _11681_);
  or _73444_ (_21874_, _21873_, _21872_);
  and _73445_ (_21875_, _08153_, \oc8051_golden_model_1.ACC [5]);
  nand _73446_ (_21876_, _21875_, _08308_);
  and _73447_ (_21877_, _21876_, _06615_);
  and _73448_ (_21878_, _21877_, _21874_);
  nor _73449_ (_21879_, _08305_, _11681_);
  or _73450_ (_21881_, _21879_, _21872_);
  or _73451_ (_21882_, _21881_, _06327_);
  and _73452_ (_21883_, _15550_, _07995_);
  or _73453_ (_21884_, _21883_, _21872_);
  or _73454_ (_21885_, _21884_, _07275_);
  or _73455_ (_21886_, _21875_, _21872_);
  and _73456_ (_21887_, _21886_, _07259_);
  and _73457_ (_21888_, _07260_, \oc8051_golden_model_1.DPH [5]);
  or _73458_ (_21889_, _21888_, _06474_);
  or _73459_ (_21890_, _21889_, _21887_);
  and _73460_ (_21892_, _21890_, _06772_);
  and _73461_ (_21893_, _21892_, _21885_);
  and _73462_ (_21894_, _21881_, _06410_);
  or _73463_ (_21895_, _21894_, _06417_);
  or _73464_ (_21896_, _21895_, _21893_);
  or _73465_ (_21897_, _21886_, _06426_);
  and _73466_ (_21898_, _21897_, _11604_);
  and _73467_ (_21899_, _21898_, _21896_);
  or _73468_ (_21900_, _11706_, \oc8051_golden_model_1.DPH [5]);
  nor _73469_ (_21901_, _11707_, _11604_);
  and _73470_ (_21903_, _21901_, _21900_);
  or _73471_ (_21904_, _21903_, _21899_);
  and _73472_ (_21905_, _21904_, _06487_);
  nor _73473_ (_21906_, _06685_, _06487_);
  or _73474_ (_21907_, _21906_, _10153_);
  or _73475_ (_21908_, _21907_, _21905_);
  and _73476_ (_21909_, _21908_, _21882_);
  or _73477_ (_21910_, _21909_, _09572_);
  and _73478_ (_21911_, _09218_, _08153_);
  or _73479_ (_21912_, _21872_, _06333_);
  or _73480_ (_21914_, _21912_, _21911_);
  and _73481_ (_21915_, _21914_, _06313_);
  and _73482_ (_21916_, _21915_, _21910_);
  and _73483_ (_21917_, _15649_, _08153_);
  or _73484_ (_21918_, _21917_, _21872_);
  and _73485_ (_21919_, _21918_, _06037_);
  or _73486_ (_21920_, _21919_, _06277_);
  or _73487_ (_21921_, _21920_, _21916_);
  and _73488_ (_21922_, _08954_, _08153_);
  or _73489_ (_21923_, _21922_, _21872_);
  or _73490_ (_21925_, _21923_, _06278_);
  and _73491_ (_21926_, _21925_, _21921_);
  or _73492_ (_21927_, _21926_, _06502_);
  and _73493_ (_21928_, _15664_, _07995_);
  or _73494_ (_21929_, _21872_, _07334_);
  or _73495_ (_21930_, _21929_, _21928_);
  and _73496_ (_21931_, _21930_, _07337_);
  and _73497_ (_21932_, _21931_, _21927_);
  or _73498_ (_21933_, _21932_, _21878_);
  and _73499_ (_21934_, _21933_, _07339_);
  or _73500_ (_21936_, _21872_, _08308_);
  and _73501_ (_21937_, _21923_, _06507_);
  and _73502_ (_21938_, _21937_, _21936_);
  or _73503_ (_21939_, _21938_, _21934_);
  and _73504_ (_21940_, _21939_, _07331_);
  and _73505_ (_21941_, _21886_, _06610_);
  and _73506_ (_21942_, _21941_, _21936_);
  or _73507_ (_21943_, _21942_, _06509_);
  or _73508_ (_21944_, _21943_, _21940_);
  and _73509_ (_21945_, _15663_, _07995_);
  or _73510_ (_21947_, _21872_, _09107_);
  or _73511_ (_21948_, _21947_, _21945_);
  and _73512_ (_21949_, _21948_, _09112_);
  and _73513_ (_21950_, _21949_, _21944_);
  and _73514_ (_21951_, _21874_, _06602_);
  or _73515_ (_21952_, _21951_, _06639_);
  or _73516_ (_21953_, _21952_, _21950_);
  or _73517_ (_21954_, _21884_, _07048_);
  and _73518_ (_21955_, _21954_, _06651_);
  and _73519_ (_21956_, _21955_, _21953_);
  and _73520_ (_21958_, _15721_, _07995_);
  or _73521_ (_21959_, _21958_, _21872_);
  and _73522_ (_21960_, _21959_, _06646_);
  or _73523_ (_21961_, _21960_, _01446_);
  or _73524_ (_21962_, _21961_, _21956_);
  or _73525_ (_21963_, _01442_, \oc8051_golden_model_1.DPH [5]);
  and _73526_ (_21964_, _21963_, _43634_);
  and _73527_ (_44162_, _21964_, _21962_);
  and _73528_ (_21965_, _11681_, \oc8051_golden_model_1.DPH [6]);
  nor _73529_ (_21966_, _08209_, _11681_);
  or _73530_ (_21968_, _21966_, _21965_);
  or _73531_ (_21969_, _21968_, _06327_);
  and _73532_ (_21970_, _15759_, _07995_);
  or _73533_ (_21971_, _21970_, _21965_);
  or _73534_ (_21972_, _21971_, _07275_);
  and _73535_ (_21973_, _08153_, \oc8051_golden_model_1.ACC [6]);
  or _73536_ (_21974_, _21973_, _21965_);
  and _73537_ (_21975_, _21974_, _07259_);
  and _73538_ (_21976_, _07260_, \oc8051_golden_model_1.DPH [6]);
  or _73539_ (_21977_, _21976_, _06474_);
  or _73540_ (_21979_, _21977_, _21975_);
  and _73541_ (_21980_, _21979_, _06772_);
  and _73542_ (_21981_, _21980_, _21972_);
  and _73543_ (_21982_, _21968_, _06410_);
  or _73544_ (_21983_, _21982_, _06417_);
  or _73545_ (_21984_, _21983_, _21981_);
  or _73546_ (_21985_, _21974_, _06426_);
  and _73547_ (_21986_, _21985_, _11604_);
  and _73548_ (_21987_, _21986_, _21984_);
  or _73549_ (_21988_, _11707_, \oc8051_golden_model_1.DPH [6]);
  nor _73550_ (_21990_, _11708_, _11604_);
  and _73551_ (_21991_, _21990_, _21988_);
  or _73552_ (_21992_, _21991_, _21987_);
  and _73553_ (_21993_, _21992_, _06487_);
  nor _73554_ (_21994_, _06487_, _06397_);
  or _73555_ (_21995_, _21994_, _10153_);
  or _73556_ (_21996_, _21995_, _21993_);
  and _73557_ (_21997_, _21996_, _21969_);
  or _73558_ (_21998_, _21997_, _09572_);
  and _73559_ (_21999_, _09172_, _08153_);
  or _73560_ (_22001_, _21965_, _06333_);
  or _73561_ (_22002_, _22001_, _21999_);
  and _73562_ (_22003_, _22002_, _06313_);
  and _73563_ (_22004_, _22003_, _21998_);
  and _73564_ (_22005_, _15846_, _08153_);
  or _73565_ (_22006_, _22005_, _21965_);
  and _73566_ (_22007_, _22006_, _06037_);
  or _73567_ (_22008_, _22007_, _06277_);
  or _73568_ (_22009_, _22008_, _22004_);
  and _73569_ (_22010_, _15853_, _08153_);
  or _73570_ (_22012_, _22010_, _21965_);
  or _73571_ (_22013_, _22012_, _06278_);
  and _73572_ (_22014_, _22013_, _22009_);
  or _73573_ (_22015_, _22014_, _06502_);
  and _73574_ (_22016_, _15862_, _07995_);
  or _73575_ (_22017_, _21965_, _07334_);
  or _73576_ (_22018_, _22017_, _22016_);
  and _73577_ (_22019_, _22018_, _07337_);
  and _73578_ (_22020_, _22019_, _22015_);
  and _73579_ (_22021_, _10596_, _08153_);
  or _73580_ (_22023_, _22021_, _21965_);
  and _73581_ (_22024_, _22023_, _06615_);
  or _73582_ (_22025_, _22024_, _22020_);
  and _73583_ (_22026_, _22025_, _07339_);
  or _73584_ (_22027_, _21965_, _08212_);
  and _73585_ (_22028_, _22012_, _06507_);
  and _73586_ (_22029_, _22028_, _22027_);
  or _73587_ (_22030_, _22029_, _22026_);
  and _73588_ (_22031_, _22030_, _07331_);
  and _73589_ (_22032_, _21974_, _06610_);
  and _73590_ (_22034_, _22032_, _22027_);
  or _73591_ (_22035_, _22034_, _06509_);
  or _73592_ (_22036_, _22035_, _22031_);
  and _73593_ (_22037_, _15859_, _07995_);
  or _73594_ (_22038_, _21965_, _09107_);
  or _73595_ (_22039_, _22038_, _22037_);
  and _73596_ (_22040_, _22039_, _09112_);
  and _73597_ (_22041_, _22040_, _22036_);
  nor _73598_ (_22042_, _10595_, _11681_);
  or _73599_ (_22043_, _22042_, _21965_);
  and _73600_ (_22045_, _22043_, _06602_);
  or _73601_ (_22046_, _22045_, _06639_);
  or _73602_ (_22047_, _22046_, _22041_);
  or _73603_ (_22048_, _21971_, _07048_);
  and _73604_ (_22049_, _22048_, _06651_);
  and _73605_ (_22050_, _22049_, _22047_);
  and _73606_ (_22051_, _15921_, _07995_);
  or _73607_ (_22052_, _22051_, _21965_);
  and _73608_ (_22053_, _22052_, _06646_);
  or _73609_ (_22054_, _22053_, _01446_);
  or _73610_ (_22056_, _22054_, _22050_);
  or _73611_ (_22057_, _01442_, \oc8051_golden_model_1.DPH [6]);
  and _73612_ (_22058_, _22057_, _43634_);
  and _73613_ (_44163_, _22058_, _22056_);
  not _73614_ (_22059_, \oc8051_golden_model_1.TL1 [0]);
  nor _73615_ (_22060_, _01442_, _22059_);
  nor _73616_ (_22061_, _07991_, _22059_);
  and _73617_ (_22062_, _07991_, _07250_);
  or _73618_ (_22063_, _22062_, _22061_);
  or _73619_ (_22064_, _22063_, _06327_);
  nor _73620_ (_22066_, _08453_, _11771_);
  or _73621_ (_22067_, _22066_, _22061_);
  or _73622_ (_22068_, _22067_, _07275_);
  and _73623_ (_22069_, _07991_, \oc8051_golden_model_1.ACC [0]);
  or _73624_ (_22070_, _22069_, _22061_);
  and _73625_ (_22071_, _22070_, _07259_);
  nor _73626_ (_22072_, _07259_, _22059_);
  or _73627_ (_22073_, _22072_, _06474_);
  or _73628_ (_22074_, _22073_, _22071_);
  and _73629_ (_22075_, _22074_, _06772_);
  and _73630_ (_22078_, _22075_, _22068_);
  and _73631_ (_22079_, _22063_, _06410_);
  or _73632_ (_22080_, _22079_, _22078_);
  and _73633_ (_22081_, _22080_, _06426_);
  and _73634_ (_22082_, _22070_, _06417_);
  or _73635_ (_22083_, _22082_, _10153_);
  or _73636_ (_22084_, _22083_, _22081_);
  and _73637_ (_22085_, _22084_, _22064_);
  or _73638_ (_22086_, _22085_, _09572_);
  and _73639_ (_22087_, _09447_, _07991_);
  or _73640_ (_22089_, _22061_, _06333_);
  or _73641_ (_22090_, _22089_, _22087_);
  and _73642_ (_22091_, _22090_, _22086_);
  or _73643_ (_22092_, _22091_, _06037_);
  and _73644_ (_22093_, _14666_, _07991_);
  or _73645_ (_22094_, _22061_, _06313_);
  or _73646_ (_22095_, _22094_, _22093_);
  and _73647_ (_22096_, _22095_, _06278_);
  and _73648_ (_22097_, _22096_, _22092_);
  and _73649_ (_22098_, _07991_, _09008_);
  or _73650_ (_22100_, _22098_, _22061_);
  and _73651_ (_22101_, _22100_, _06277_);
  or _73652_ (_22102_, _22101_, _06502_);
  or _73653_ (_22103_, _22102_, _22097_);
  and _73654_ (_22104_, _14566_, _07991_);
  or _73655_ (_22105_, _22061_, _07334_);
  or _73656_ (_22106_, _22105_, _22104_);
  and _73657_ (_22107_, _22106_, _07337_);
  and _73658_ (_22108_, _22107_, _22103_);
  nor _73659_ (_22109_, _12622_, _11771_);
  or _73660_ (_22111_, _22109_, _22061_);
  and _73661_ (_22112_, _10577_, _07991_);
  nor _73662_ (_22113_, _22112_, _07337_);
  and _73663_ (_22114_, _22113_, _22111_);
  or _73664_ (_22115_, _22114_, _22108_);
  and _73665_ (_22116_, _22115_, _07339_);
  nand _73666_ (_22117_, _22100_, _06507_);
  nor _73667_ (_22118_, _22117_, _22066_);
  or _73668_ (_22119_, _22118_, _06610_);
  or _73669_ (_22120_, _22119_, _22116_);
  or _73670_ (_22122_, _22112_, _22061_);
  or _73671_ (_22123_, _22122_, _07331_);
  and _73672_ (_22124_, _22123_, _22120_);
  or _73673_ (_22125_, _22124_, _06509_);
  and _73674_ (_22126_, _14563_, _07991_);
  or _73675_ (_22127_, _22061_, _09107_);
  or _73676_ (_22128_, _22127_, _22126_);
  and _73677_ (_22129_, _22128_, _09112_);
  and _73678_ (_22130_, _22129_, _22125_);
  and _73679_ (_22131_, _22111_, _06602_);
  or _73680_ (_22133_, _22131_, _19642_);
  or _73681_ (_22134_, _22133_, _22130_);
  or _73682_ (_22135_, _22067_, _19641_);
  and _73683_ (_22136_, _22135_, _01442_);
  and _73684_ (_22137_, _22136_, _22134_);
  or _73685_ (_22138_, _22137_, _22060_);
  and _73686_ (_44164_, _22138_, _43634_);
  not _73687_ (_22139_, \oc8051_golden_model_1.TL1 [1]);
  nor _73688_ (_22140_, _01442_, _22139_);
  or _73689_ (_22141_, _14851_, _11771_);
  or _73690_ (_22143_, _07991_, \oc8051_golden_model_1.TL1 [1]);
  and _73691_ (_22144_, _22143_, _06037_);
  and _73692_ (_22145_, _22144_, _22141_);
  and _73693_ (_22146_, _14744_, _07991_);
  not _73694_ (_22147_, _22146_);
  and _73695_ (_22148_, _22147_, _22143_);
  or _73696_ (_22149_, _22148_, _07275_);
  nor _73697_ (_22150_, _07991_, _22139_);
  and _73698_ (_22151_, _07991_, \oc8051_golden_model_1.ACC [1]);
  or _73699_ (_22152_, _22151_, _22150_);
  and _73700_ (_22154_, _22152_, _07259_);
  nor _73701_ (_22155_, _07259_, _22139_);
  or _73702_ (_22156_, _22155_, _06474_);
  or _73703_ (_22157_, _22156_, _22154_);
  and _73704_ (_22158_, _22157_, _06772_);
  and _73705_ (_22159_, _22158_, _22149_);
  nor _73706_ (_22160_, _11771_, _07448_);
  or _73707_ (_22161_, _22160_, _22150_);
  and _73708_ (_22162_, _22161_, _06410_);
  or _73709_ (_22163_, _22162_, _22159_);
  and _73710_ (_22164_, _22163_, _06426_);
  and _73711_ (_22165_, _22152_, _06417_);
  or _73712_ (_22166_, _22165_, _10153_);
  or _73713_ (_22167_, _22166_, _22164_);
  or _73714_ (_22168_, _22161_, _06327_);
  and _73715_ (_22169_, _22168_, _16672_);
  and _73716_ (_22170_, _22169_, _22167_);
  or _73717_ (_22171_, _09402_, _11771_);
  and _73718_ (_22172_, _22143_, _14025_);
  and _73719_ (_22173_, _22172_, _22171_);
  or _73720_ (_22176_, _22173_, _22170_);
  and _73721_ (_22177_, _22176_, _06313_);
  or _73722_ (_22178_, _22177_, _22145_);
  and _73723_ (_22179_, _22178_, _06278_);
  nand _73724_ (_22180_, _07991_, _07160_);
  and _73725_ (_22181_, _22143_, _06277_);
  and _73726_ (_22182_, _22181_, _22180_);
  or _73727_ (_22183_, _22182_, _22179_);
  and _73728_ (_22184_, _22183_, _07334_);
  or _73729_ (_22185_, _14749_, _11771_);
  and _73730_ (_22187_, _22143_, _06502_);
  and _73731_ (_22188_, _22187_, _22185_);
  or _73732_ (_22189_, _22188_, _06615_);
  or _73733_ (_22190_, _22189_, _22184_);
  nor _73734_ (_22191_, _10578_, _11771_);
  or _73735_ (_22192_, _22191_, _22150_);
  nand _73736_ (_22193_, _10576_, _07991_);
  and _73737_ (_22194_, _22193_, _22192_);
  or _73738_ (_22195_, _22194_, _07337_);
  and _73739_ (_22196_, _22195_, _07339_);
  and _73740_ (_22198_, _22196_, _22190_);
  or _73741_ (_22199_, _14747_, _11771_);
  and _73742_ (_22200_, _22143_, _06507_);
  and _73743_ (_22201_, _22200_, _22199_);
  or _73744_ (_22202_, _22201_, _06610_);
  or _73745_ (_22203_, _22202_, _22198_);
  nor _73746_ (_22204_, _22150_, _07331_);
  nand _73747_ (_22205_, _22204_, _22193_);
  and _73748_ (_22206_, _22205_, _09107_);
  and _73749_ (_22207_, _22206_, _22203_);
  or _73750_ (_22209_, _22180_, _08404_);
  and _73751_ (_22210_, _22143_, _06509_);
  and _73752_ (_22211_, _22210_, _22209_);
  or _73753_ (_22212_, _22211_, _06602_);
  or _73754_ (_22213_, _22212_, _22207_);
  or _73755_ (_22214_, _22192_, _09112_);
  and _73756_ (_22215_, _22214_, _07048_);
  and _73757_ (_22216_, _22215_, _22213_);
  and _73758_ (_22217_, _22148_, _06639_);
  or _73759_ (_22218_, _22217_, _06646_);
  or _73760_ (_22220_, _22218_, _22216_);
  or _73761_ (_22221_, _22150_, _06651_);
  or _73762_ (_22222_, _22221_, _22146_);
  and _73763_ (_22223_, _22222_, _01442_);
  and _73764_ (_22224_, _22223_, _22220_);
  or _73765_ (_22225_, _22224_, _22140_);
  and _73766_ (_44166_, _22225_, _43634_);
  not _73767_ (_22226_, \oc8051_golden_model_1.TL1 [2]);
  nor _73768_ (_22227_, _01442_, _22226_);
  nor _73769_ (_22228_, _07991_, _22226_);
  or _73770_ (_22230_, _22228_, _08503_);
  and _73771_ (_22231_, _07991_, _09057_);
  or _73772_ (_22232_, _22231_, _22228_);
  and _73773_ (_22233_, _22232_, _06507_);
  and _73774_ (_22234_, _22233_, _22230_);
  nor _73775_ (_22235_, _10582_, _11771_);
  or _73776_ (_22236_, _22235_, _22228_);
  and _73777_ (_22237_, _07991_, \oc8051_golden_model_1.ACC [2]);
  nand _73778_ (_22238_, _22237_, _08503_);
  and _73779_ (_22239_, _22238_, _06615_);
  and _73780_ (_22241_, _22239_, _22236_);
  nor _73781_ (_22242_, _11771_, _07854_);
  or _73782_ (_22243_, _22242_, _22228_);
  or _73783_ (_22244_, _22243_, _06327_);
  and _73784_ (_22245_, _14959_, _07991_);
  or _73785_ (_22246_, _22245_, _22228_);
  and _73786_ (_22247_, _22246_, _06474_);
  nor _73787_ (_22248_, _07259_, _22226_);
  or _73788_ (_22249_, _22237_, _22228_);
  and _73789_ (_22250_, _22249_, _07259_);
  or _73790_ (_22252_, _22250_, _22248_);
  and _73791_ (_22253_, _22252_, _07275_);
  or _73792_ (_22254_, _22253_, _06410_);
  or _73793_ (_22255_, _22254_, _22247_);
  or _73794_ (_22256_, _22243_, _06772_);
  and _73795_ (_22257_, _22256_, _06426_);
  and _73796_ (_22258_, _22257_, _22255_);
  and _73797_ (_22259_, _22249_, _06417_);
  or _73798_ (_22260_, _22259_, _10153_);
  or _73799_ (_22261_, _22260_, _22258_);
  and _73800_ (_22263_, _22261_, _22244_);
  or _73801_ (_22264_, _22263_, _09572_);
  and _73802_ (_22265_, _09356_, _07991_);
  or _73803_ (_22266_, _22228_, _06333_);
  or _73804_ (_22267_, _22266_, _22265_);
  and _73805_ (_22268_, _22267_, _22264_);
  or _73806_ (_22269_, _22268_, _06037_);
  and _73807_ (_22270_, _15056_, _07991_);
  or _73808_ (_22271_, _22228_, _06313_);
  or _73809_ (_22272_, _22271_, _22270_);
  and _73810_ (_22274_, _22272_, _06278_);
  and _73811_ (_22275_, _22274_, _22269_);
  and _73812_ (_22276_, _22232_, _06277_);
  or _73813_ (_22277_, _22276_, _06502_);
  or _73814_ (_22278_, _22277_, _22275_);
  and _73815_ (_22279_, _14948_, _07991_);
  or _73816_ (_22280_, _22228_, _07334_);
  or _73817_ (_22281_, _22280_, _22279_);
  and _73818_ (_22282_, _22281_, _07337_);
  and _73819_ (_22283_, _22282_, _22278_);
  or _73820_ (_22285_, _22283_, _22241_);
  and _73821_ (_22286_, _22285_, _07339_);
  or _73822_ (_22287_, _22286_, _22234_);
  and _73823_ (_22288_, _22287_, _07331_);
  and _73824_ (_22289_, _22249_, _06610_);
  and _73825_ (_22290_, _22289_, _22230_);
  or _73826_ (_22291_, _22290_, _06509_);
  or _73827_ (_22292_, _22291_, _22288_);
  and _73828_ (_22293_, _14945_, _07991_);
  or _73829_ (_22294_, _22228_, _09107_);
  or _73830_ (_22296_, _22294_, _22293_);
  and _73831_ (_22297_, _22296_, _09112_);
  and _73832_ (_22298_, _22297_, _22292_);
  and _73833_ (_22299_, _22236_, _06602_);
  or _73834_ (_22300_, _22299_, _22298_);
  and _73835_ (_22301_, _22300_, _07048_);
  and _73836_ (_22302_, _22246_, _06639_);
  or _73837_ (_22303_, _22302_, _06646_);
  or _73838_ (_22304_, _22303_, _22301_);
  and _73839_ (_22305_, _15129_, _07991_);
  or _73840_ (_22307_, _22228_, _06651_);
  or _73841_ (_22308_, _22307_, _22305_);
  and _73842_ (_22309_, _22308_, _01442_);
  and _73843_ (_22310_, _22309_, _22304_);
  or _73844_ (_22311_, _22310_, _22227_);
  and _73845_ (_44167_, _22311_, _43634_);
  and _73846_ (_22312_, _11771_, \oc8051_golden_model_1.TL1 [3]);
  or _73847_ (_22313_, _22312_, _08359_);
  and _73848_ (_22314_, _07991_, _09014_);
  or _73849_ (_22315_, _22314_, _22312_);
  and _73850_ (_22317_, _22315_, _06507_);
  and _73851_ (_22318_, _22317_, _22313_);
  and _73852_ (_22319_, _15153_, _07991_);
  or _73853_ (_22320_, _22319_, _22312_);
  or _73854_ (_22321_, _22320_, _07275_);
  and _73855_ (_22322_, _07991_, \oc8051_golden_model_1.ACC [3]);
  or _73856_ (_22323_, _22322_, _22312_);
  and _73857_ (_22324_, _22323_, _07259_);
  and _73858_ (_22325_, _07260_, \oc8051_golden_model_1.TL1 [3]);
  or _73859_ (_22326_, _22325_, _06474_);
  or _73860_ (_22328_, _22326_, _22324_);
  and _73861_ (_22329_, _22328_, _06772_);
  and _73862_ (_22330_, _22329_, _22321_);
  nor _73863_ (_22331_, _11771_, _07680_);
  or _73864_ (_22332_, _22331_, _22312_);
  and _73865_ (_22333_, _22332_, _06410_);
  or _73866_ (_22334_, _22333_, _22330_);
  and _73867_ (_22335_, _22334_, _06426_);
  and _73868_ (_22336_, _22323_, _06417_);
  or _73869_ (_22337_, _22336_, _10153_);
  or _73870_ (_22339_, _22337_, _22335_);
  or _73871_ (_22340_, _22332_, _06327_);
  and _73872_ (_22341_, _22340_, _22339_);
  or _73873_ (_22342_, _22341_, _09572_);
  and _73874_ (_22343_, _09310_, _07991_);
  or _73875_ (_22344_, _22312_, _06333_);
  or _73876_ (_22345_, _22344_, _22343_);
  and _73877_ (_22346_, _22345_, _06313_);
  and _73878_ (_22347_, _22346_, _22342_);
  and _73879_ (_22348_, _15251_, _07991_);
  or _73880_ (_22350_, _22348_, _22312_);
  and _73881_ (_22351_, _22350_, _06037_);
  or _73882_ (_22352_, _22351_, _06277_);
  or _73883_ (_22353_, _22352_, _22347_);
  or _73884_ (_22354_, _22315_, _06278_);
  and _73885_ (_22355_, _22354_, _22353_);
  or _73886_ (_22356_, _22355_, _06502_);
  and _73887_ (_22357_, _15266_, _07991_);
  or _73888_ (_22358_, _22312_, _07334_);
  or _73889_ (_22359_, _22358_, _22357_);
  and _73890_ (_22361_, _22359_, _07337_);
  and _73891_ (_22362_, _22361_, _22356_);
  and _73892_ (_22363_, _12619_, _07991_);
  or _73893_ (_22364_, _22363_, _22312_);
  and _73894_ (_22365_, _22364_, _06615_);
  or _73895_ (_22366_, _22365_, _22362_);
  and _73896_ (_22367_, _22366_, _07339_);
  or _73897_ (_22368_, _22367_, _22318_);
  and _73898_ (_22369_, _22368_, _07331_);
  and _73899_ (_22370_, _22323_, _06610_);
  and _73900_ (_22372_, _22370_, _22313_);
  or _73901_ (_22373_, _22372_, _06509_);
  or _73902_ (_22374_, _22373_, _22369_);
  and _73903_ (_22375_, _15263_, _07991_);
  or _73904_ (_22376_, _22312_, _09107_);
  or _73905_ (_22377_, _22376_, _22375_);
  and _73906_ (_22378_, _22377_, _09112_);
  and _73907_ (_22379_, _22378_, _22374_);
  nor _73908_ (_22380_, _10574_, _11771_);
  or _73909_ (_22381_, _22380_, _22312_);
  and _73910_ (_22383_, _22381_, _06602_);
  or _73911_ (_22384_, _22383_, _06639_);
  or _73912_ (_22385_, _22384_, _22379_);
  or _73913_ (_22386_, _22320_, _07048_);
  and _73914_ (_22387_, _22386_, _06651_);
  and _73915_ (_22388_, _22387_, _22385_);
  and _73916_ (_22389_, _15321_, _07991_);
  or _73917_ (_22390_, _22389_, _22312_);
  and _73918_ (_22391_, _22390_, _06646_);
  or _73919_ (_22392_, _22391_, _01446_);
  or _73920_ (_22394_, _22392_, _22388_);
  or _73921_ (_22395_, _01442_, \oc8051_golden_model_1.TL1 [3]);
  and _73922_ (_22396_, _22395_, _43634_);
  and _73923_ (_44168_, _22396_, _22394_);
  and _73924_ (_22397_, _11771_, \oc8051_golden_model_1.TL1 [4]);
  or _73925_ (_22398_, _22397_, _08599_);
  and _73926_ (_22399_, _08995_, _07991_);
  or _73927_ (_22400_, _22399_, _22397_);
  and _73928_ (_22401_, _22400_, _06507_);
  and _73929_ (_22402_, _22401_, _22398_);
  and _73930_ (_22404_, _15367_, _07991_);
  or _73931_ (_22405_, _22404_, _22397_);
  or _73932_ (_22406_, _22405_, _07275_);
  and _73933_ (_22407_, _07991_, \oc8051_golden_model_1.ACC [4]);
  or _73934_ (_22408_, _22407_, _22397_);
  and _73935_ (_22409_, _22408_, _07259_);
  and _73936_ (_22410_, _07260_, \oc8051_golden_model_1.TL1 [4]);
  or _73937_ (_22411_, _22410_, _06474_);
  or _73938_ (_22412_, _22411_, _22409_);
  and _73939_ (_22413_, _22412_, _06772_);
  and _73940_ (_22415_, _22413_, _22406_);
  nor _73941_ (_22416_, _08596_, _11771_);
  or _73942_ (_22417_, _22416_, _22397_);
  and _73943_ (_22418_, _22417_, _06410_);
  or _73944_ (_22419_, _22418_, _22415_);
  and _73945_ (_22420_, _22419_, _06426_);
  and _73946_ (_22421_, _22408_, _06417_);
  or _73947_ (_22422_, _22421_, _10153_);
  or _73948_ (_22423_, _22422_, _22420_);
  or _73949_ (_22424_, _22417_, _06327_);
  and _73950_ (_22426_, _22424_, _22423_);
  or _73951_ (_22427_, _22426_, _09572_);
  and _73952_ (_22428_, _09264_, _07991_);
  or _73953_ (_22429_, _22397_, _16672_);
  or _73954_ (_22430_, _22429_, _22428_);
  and _73955_ (_22431_, _22430_, _22427_);
  or _73956_ (_22432_, _22431_, _06037_);
  and _73957_ (_22433_, _15452_, _07991_);
  or _73958_ (_22434_, _22397_, _06313_);
  or _73959_ (_22435_, _22434_, _22433_);
  and _73960_ (_22437_, _22435_, _06278_);
  and _73961_ (_22438_, _22437_, _22432_);
  and _73962_ (_22439_, _22400_, _06277_);
  or _73963_ (_22440_, _22439_, _06502_);
  or _73964_ (_22441_, _22440_, _22438_);
  and _73965_ (_22442_, _15345_, _07991_);
  or _73966_ (_22443_, _22397_, _07334_);
  or _73967_ (_22444_, _22443_, _22442_);
  and _73968_ (_22445_, _22444_, _07337_);
  and _73969_ (_22446_, _22445_, _22441_);
  and _73970_ (_22448_, _10590_, _07991_);
  or _73971_ (_22449_, _22448_, _22397_);
  and _73972_ (_22450_, _22449_, _06615_);
  or _73973_ (_22451_, _22450_, _22446_);
  and _73974_ (_22452_, _22451_, _07339_);
  or _73975_ (_22453_, _22452_, _22402_);
  and _73976_ (_22454_, _22453_, _07331_);
  and _73977_ (_22455_, _22408_, _06610_);
  and _73978_ (_22456_, _22455_, _22398_);
  or _73979_ (_22457_, _22456_, _06509_);
  or _73980_ (_22458_, _22457_, _22454_);
  and _73981_ (_22459_, _15342_, _07991_);
  or _73982_ (_22460_, _22397_, _09107_);
  or _73983_ (_22461_, _22460_, _22459_);
  and _73984_ (_22462_, _22461_, _09112_);
  and _73985_ (_22463_, _22462_, _22458_);
  nor _73986_ (_22464_, _10589_, _11771_);
  or _73987_ (_22465_, _22464_, _22397_);
  and _73988_ (_22466_, _22465_, _06602_);
  or _73989_ (_22467_, _22466_, _06639_);
  or _73990_ (_22470_, _22467_, _22463_);
  or _73991_ (_22471_, _22405_, _07048_);
  and _73992_ (_22472_, _22471_, _06651_);
  and _73993_ (_22473_, _22472_, _22470_);
  and _73994_ (_22474_, _15524_, _07991_);
  or _73995_ (_22475_, _22474_, _22397_);
  and _73996_ (_22476_, _22475_, _06646_);
  or _73997_ (_22477_, _22476_, _01446_);
  or _73998_ (_22478_, _22477_, _22473_);
  or _73999_ (_22479_, _01442_, \oc8051_golden_model_1.TL1 [4]);
  and _74000_ (_22481_, _22479_, _43634_);
  and _74001_ (_44169_, _22481_, _22478_);
  and _74002_ (_22482_, _11771_, \oc8051_golden_model_1.TL1 [5]);
  and _74003_ (_22483_, _15550_, _07991_);
  or _74004_ (_22484_, _22483_, _22482_);
  or _74005_ (_22485_, _22484_, _07275_);
  and _74006_ (_22486_, _07991_, \oc8051_golden_model_1.ACC [5]);
  or _74007_ (_22487_, _22486_, _22482_);
  and _74008_ (_22488_, _22487_, _07259_);
  and _74009_ (_22489_, _07260_, \oc8051_golden_model_1.TL1 [5]);
  or _74010_ (_22491_, _22489_, _06474_);
  or _74011_ (_22492_, _22491_, _22488_);
  and _74012_ (_22493_, _22492_, _06772_);
  and _74013_ (_22494_, _22493_, _22485_);
  nor _74014_ (_22495_, _08305_, _11771_);
  or _74015_ (_22496_, _22495_, _22482_);
  and _74016_ (_22497_, _22496_, _06410_);
  or _74017_ (_22498_, _22497_, _22494_);
  and _74018_ (_22499_, _22498_, _06426_);
  and _74019_ (_22500_, _22487_, _06417_);
  or _74020_ (_22502_, _22500_, _10153_);
  or _74021_ (_22503_, _22502_, _22499_);
  or _74022_ (_22504_, _22496_, _06327_);
  and _74023_ (_22505_, _22504_, _22503_);
  or _74024_ (_22506_, _22505_, _09572_);
  and _74025_ (_22507_, _09218_, _07991_);
  or _74026_ (_22508_, _22482_, _06333_);
  or _74027_ (_22509_, _22508_, _22507_);
  and _74028_ (_22510_, _22509_, _06313_);
  and _74029_ (_22511_, _22510_, _22506_);
  and _74030_ (_22513_, _15649_, _07991_);
  or _74031_ (_22514_, _22513_, _22482_);
  and _74032_ (_22515_, _22514_, _06037_);
  or _74033_ (_22516_, _22515_, _06277_);
  or _74034_ (_22517_, _22516_, _22511_);
  and _74035_ (_22518_, _08954_, _07991_);
  or _74036_ (_22519_, _22518_, _22482_);
  or _74037_ (_22520_, _22519_, _06278_);
  and _74038_ (_22521_, _22520_, _22517_);
  or _74039_ (_22522_, _22521_, _06502_);
  and _74040_ (_22524_, _15664_, _07991_);
  or _74041_ (_22525_, _22482_, _07334_);
  or _74042_ (_22526_, _22525_, _22524_);
  and _74043_ (_22527_, _22526_, _07337_);
  and _74044_ (_22528_, _22527_, _22522_);
  and _74045_ (_22529_, _12626_, _07991_);
  or _74046_ (_22530_, _22529_, _22482_);
  and _74047_ (_22531_, _22530_, _06615_);
  or _74048_ (_22532_, _22531_, _22528_);
  and _74049_ (_22533_, _22532_, _07339_);
  or _74050_ (_22535_, _22482_, _08308_);
  and _74051_ (_22536_, _22519_, _06507_);
  and _74052_ (_22537_, _22536_, _22535_);
  or _74053_ (_22538_, _22537_, _22533_);
  and _74054_ (_22539_, _22538_, _07331_);
  and _74055_ (_22540_, _22487_, _06610_);
  and _74056_ (_22541_, _22540_, _22535_);
  or _74057_ (_22542_, _22541_, _06509_);
  or _74058_ (_22543_, _22542_, _22539_);
  and _74059_ (_22544_, _15663_, _07991_);
  or _74060_ (_22546_, _22482_, _09107_);
  or _74061_ (_22547_, _22546_, _22544_);
  and _74062_ (_22548_, _22547_, _09112_);
  and _74063_ (_22549_, _22548_, _22543_);
  nor _74064_ (_22550_, _10570_, _11771_);
  or _74065_ (_22551_, _22550_, _22482_);
  and _74066_ (_22552_, _22551_, _06602_);
  or _74067_ (_22553_, _22552_, _06639_);
  or _74068_ (_22554_, _22553_, _22549_);
  or _74069_ (_22555_, _22484_, _07048_);
  and _74070_ (_22557_, _22555_, _06651_);
  and _74071_ (_22558_, _22557_, _22554_);
  and _74072_ (_22559_, _15721_, _07991_);
  or _74073_ (_22560_, _22559_, _22482_);
  and _74074_ (_22561_, _22560_, _06646_);
  or _74075_ (_22562_, _22561_, _01446_);
  or _74076_ (_22563_, _22562_, _22558_);
  or _74077_ (_22564_, _01442_, \oc8051_golden_model_1.TL1 [5]);
  and _74078_ (_22565_, _22564_, _43634_);
  and _74079_ (_44170_, _22565_, _22563_);
  and _74080_ (_22566_, _11771_, \oc8051_golden_model_1.TL1 [6]);
  and _74081_ (_22567_, _15759_, _07991_);
  or _74082_ (_22568_, _22567_, _22566_);
  or _74083_ (_22569_, _22568_, _07275_);
  and _74084_ (_22570_, _07991_, \oc8051_golden_model_1.ACC [6]);
  or _74085_ (_22571_, _22570_, _22566_);
  and _74086_ (_22572_, _22571_, _07259_);
  and _74087_ (_22573_, _07260_, \oc8051_golden_model_1.TL1 [6]);
  or _74088_ (_22574_, _22573_, _06474_);
  or _74089_ (_22575_, _22574_, _22572_);
  and _74090_ (_22578_, _22575_, _06772_);
  and _74091_ (_22579_, _22578_, _22569_);
  nor _74092_ (_22580_, _08209_, _11771_);
  or _74093_ (_22581_, _22580_, _22566_);
  and _74094_ (_22582_, _22581_, _06410_);
  or _74095_ (_22583_, _22582_, _22579_);
  and _74096_ (_22584_, _22583_, _06426_);
  and _74097_ (_22585_, _22571_, _06417_);
  or _74098_ (_22586_, _22585_, _10153_);
  or _74099_ (_22587_, _22586_, _22584_);
  or _74100_ (_22589_, _22581_, _06327_);
  and _74101_ (_22590_, _22589_, _22587_);
  or _74102_ (_22591_, _22590_, _09572_);
  and _74103_ (_22592_, _09172_, _07991_);
  or _74104_ (_22593_, _22566_, _06333_);
  or _74105_ (_22594_, _22593_, _22592_);
  and _74106_ (_22595_, _22594_, _06313_);
  and _74107_ (_22596_, _22595_, _22591_);
  and _74108_ (_22597_, _15846_, _07991_);
  or _74109_ (_22598_, _22597_, _22566_);
  and _74110_ (_22600_, _22598_, _06037_);
  or _74111_ (_22601_, _22600_, _06277_);
  or _74112_ (_22602_, _22601_, _22596_);
  and _74113_ (_22603_, _15853_, _07991_);
  or _74114_ (_22604_, _22603_, _22566_);
  or _74115_ (_22605_, _22604_, _06278_);
  and _74116_ (_22606_, _22605_, _22602_);
  or _74117_ (_22607_, _22606_, _06502_);
  and _74118_ (_22608_, _15862_, _07991_);
  or _74119_ (_22609_, _22566_, _07334_);
  or _74120_ (_22611_, _22609_, _22608_);
  and _74121_ (_22612_, _22611_, _07337_);
  and _74122_ (_22613_, _22612_, _22607_);
  and _74123_ (_22614_, _10596_, _07991_);
  or _74124_ (_22615_, _22614_, _22566_);
  and _74125_ (_22616_, _22615_, _06615_);
  or _74126_ (_22617_, _22616_, _22613_);
  and _74127_ (_22618_, _22617_, _07339_);
  or _74128_ (_22619_, _22566_, _08212_);
  and _74129_ (_22620_, _22604_, _06507_);
  and _74130_ (_22622_, _22620_, _22619_);
  or _74131_ (_22623_, _22622_, _22618_);
  and _74132_ (_22624_, _22623_, _07331_);
  and _74133_ (_22625_, _22571_, _06610_);
  and _74134_ (_22626_, _22625_, _22619_);
  or _74135_ (_22627_, _22626_, _06509_);
  or _74136_ (_22628_, _22627_, _22624_);
  and _74137_ (_22629_, _15859_, _07991_);
  or _74138_ (_22630_, _22566_, _09107_);
  or _74139_ (_22631_, _22630_, _22629_);
  and _74140_ (_22633_, _22631_, _09112_);
  and _74141_ (_22634_, _22633_, _22628_);
  nor _74142_ (_22635_, _10595_, _11771_);
  or _74143_ (_22636_, _22635_, _22566_);
  and _74144_ (_22637_, _22636_, _06602_);
  or _74145_ (_22638_, _22637_, _06639_);
  or _74146_ (_22639_, _22638_, _22634_);
  or _74147_ (_22640_, _22568_, _07048_);
  and _74148_ (_22641_, _22640_, _06651_);
  and _74149_ (_22642_, _22641_, _22639_);
  and _74150_ (_22644_, _15921_, _07991_);
  or _74151_ (_22645_, _22644_, _22566_);
  and _74152_ (_22646_, _22645_, _06646_);
  or _74153_ (_22647_, _22646_, _01446_);
  or _74154_ (_22648_, _22647_, _22642_);
  or _74155_ (_22649_, _01442_, \oc8051_golden_model_1.TL1 [6]);
  and _74156_ (_22650_, _22649_, _43634_);
  and _74157_ (_44171_, _22650_, _22648_);
  and _74158_ (_22651_, _01446_, \oc8051_golden_model_1.TL0 [0]);
  and _74159_ (_22652_, _11849_, \oc8051_golden_model_1.TL0 [0]);
  nor _74160_ (_22654_, _12622_, _11854_);
  or _74161_ (_22655_, _22654_, _22652_);
  and _74162_ (_22656_, _08133_, \oc8051_golden_model_1.ACC [0]);
  and _74163_ (_22657_, _22656_, _08453_);
  nor _74164_ (_22658_, _22657_, _07337_);
  and _74165_ (_22659_, _22658_, _22655_);
  or _74166_ (_22660_, _22656_, _22652_);
  and _74167_ (_22661_, _22660_, _06417_);
  or _74168_ (_22662_, _22661_, _10153_);
  nor _74169_ (_22663_, _08453_, _11854_);
  or _74170_ (_22665_, _22663_, _22652_);
  and _74171_ (_22666_, _22665_, _06474_);
  and _74172_ (_22667_, _07260_, \oc8051_golden_model_1.TL0 [0]);
  and _74173_ (_22668_, _22660_, _07259_);
  or _74174_ (_22669_, _22668_, _22667_);
  and _74175_ (_22670_, _22669_, _07275_);
  or _74176_ (_22671_, _22670_, _06410_);
  or _74177_ (_22672_, _22671_, _22666_);
  and _74178_ (_22673_, _22672_, _06426_);
  or _74179_ (_22674_, _22673_, _22662_);
  and _74180_ (_22676_, _07976_, _07250_);
  or _74181_ (_22677_, _22652_, _19597_);
  or _74182_ (_22678_, _22677_, _22676_);
  and _74183_ (_22679_, _22678_, _22674_);
  or _74184_ (_22680_, _22679_, _09572_);
  and _74185_ (_22681_, _09447_, _08133_);
  or _74186_ (_22682_, _22652_, _06333_);
  or _74187_ (_22683_, _22682_, _22681_);
  and _74188_ (_22684_, _22683_, _22680_);
  or _74189_ (_22685_, _22684_, _06037_);
  and _74190_ (_22687_, _14666_, _07976_);
  or _74191_ (_22688_, _22652_, _06313_);
  or _74192_ (_22689_, _22688_, _22687_);
  and _74193_ (_22690_, _22689_, _06278_);
  and _74194_ (_22691_, _22690_, _22685_);
  and _74195_ (_22692_, _08133_, _09008_);
  or _74196_ (_22693_, _22692_, _22652_);
  and _74197_ (_22694_, _22693_, _06277_);
  or _74198_ (_22695_, _22694_, _06502_);
  or _74199_ (_22696_, _22695_, _22691_);
  and _74200_ (_22698_, _14566_, _07976_);
  or _74201_ (_22699_, _22652_, _07334_);
  or _74202_ (_22700_, _22699_, _22698_);
  and _74203_ (_22701_, _22700_, _07337_);
  and _74204_ (_22702_, _22701_, _22696_);
  or _74205_ (_22703_, _22702_, _22659_);
  and _74206_ (_22704_, _22703_, _07339_);
  nand _74207_ (_22705_, _22693_, _06507_);
  nor _74208_ (_22706_, _22705_, _22663_);
  or _74209_ (_22707_, _22706_, _06610_);
  or _74210_ (_22709_, _22707_, _22704_);
  or _74211_ (_22710_, _22657_, _22652_);
  or _74212_ (_22711_, _22710_, _07331_);
  and _74213_ (_22712_, _22711_, _22709_);
  or _74214_ (_22713_, _22712_, _06509_);
  and _74215_ (_22714_, _14563_, _07976_);
  or _74216_ (_22715_, _22652_, _09107_);
  or _74217_ (_22716_, _22715_, _22714_);
  and _74218_ (_22717_, _22716_, _09112_);
  and _74219_ (_22718_, _22717_, _22713_);
  and _74220_ (_22720_, _22655_, _06602_);
  or _74221_ (_22721_, _22720_, _19642_);
  or _74222_ (_22722_, _22721_, _22718_);
  or _74223_ (_22723_, _22665_, _19641_);
  and _74224_ (_22724_, _22723_, _01442_);
  and _74225_ (_22725_, _22724_, _22722_);
  or _74226_ (_22726_, _22725_, _22651_);
  and _74227_ (_44172_, _22726_, _43634_);
  and _74228_ (_22727_, _01446_, \oc8051_golden_model_1.TL0 [1]);
  or _74229_ (_22728_, _08133_, \oc8051_golden_model_1.TL0 [1]);
  nand _74230_ (_22730_, _14744_, _07976_);
  and _74231_ (_22731_, _22730_, _22728_);
  or _74232_ (_22732_, _22731_, _07275_);
  and _74233_ (_22733_, _11849_, \oc8051_golden_model_1.TL0 [1]);
  and _74234_ (_22734_, _08133_, \oc8051_golden_model_1.ACC [1]);
  or _74235_ (_22735_, _22734_, _22733_);
  and _74236_ (_22736_, _22735_, _07259_);
  and _74237_ (_22737_, _07260_, \oc8051_golden_model_1.TL0 [1]);
  or _74238_ (_22738_, _22737_, _06474_);
  or _74239_ (_22739_, _22738_, _22736_);
  and _74240_ (_22741_, _22739_, _06772_);
  and _74241_ (_22742_, _22741_, _22732_);
  nor _74242_ (_22743_, _11854_, _07448_);
  or _74243_ (_22744_, _22743_, _22733_);
  and _74244_ (_22745_, _22744_, _06410_);
  or _74245_ (_22746_, _22745_, _22742_);
  and _74246_ (_22747_, _22746_, _06426_);
  and _74247_ (_22748_, _22735_, _06417_);
  or _74248_ (_22749_, _22748_, _10153_);
  or _74249_ (_22750_, _22749_, _22747_);
  or _74250_ (_22752_, _22744_, _06327_);
  and _74251_ (_22753_, _22752_, _22750_);
  or _74252_ (_22754_, _22753_, _09572_);
  and _74253_ (_22755_, _22754_, _06313_);
  and _74254_ (_22756_, _09402_, _08133_);
  or _74255_ (_22757_, _22733_, _06333_);
  or _74256_ (_22758_, _22757_, _22756_);
  and _74257_ (_22759_, _22758_, _22755_);
  and _74258_ (_22760_, _14851_, _08133_);
  or _74259_ (_22761_, _22760_, _22733_);
  and _74260_ (_22763_, _22761_, _06037_);
  or _74261_ (_22764_, _22763_, _22759_);
  and _74262_ (_22765_, _22764_, _06278_);
  and _74263_ (_22766_, _22728_, _06277_);
  nand _74264_ (_22767_, _07976_, _07160_);
  and _74265_ (_22768_, _22767_, _22766_);
  or _74266_ (_22769_, _22768_, _22765_);
  and _74267_ (_22770_, _22769_, _07334_);
  or _74268_ (_22771_, _14749_, _11854_);
  and _74269_ (_22772_, _22728_, _06502_);
  and _74270_ (_22774_, _22772_, _22771_);
  or _74271_ (_22775_, _22774_, _06615_);
  or _74272_ (_22776_, _22775_, _22770_);
  nor _74273_ (_22777_, _10578_, _11854_);
  or _74274_ (_22778_, _22777_, _22733_);
  nand _74275_ (_22779_, _10576_, _07976_);
  and _74276_ (_22780_, _22779_, _22778_);
  or _74277_ (_22781_, _22780_, _07337_);
  and _74278_ (_22782_, _22781_, _07339_);
  and _74279_ (_22783_, _22782_, _22776_);
  or _74280_ (_22784_, _14747_, _11854_);
  and _74281_ (_22785_, _22728_, _06507_);
  and _74282_ (_22786_, _22785_, _22784_);
  or _74283_ (_22787_, _22786_, _06610_);
  or _74284_ (_22788_, _22787_, _22783_);
  nor _74285_ (_22789_, _22733_, _07331_);
  nand _74286_ (_22790_, _22789_, _22779_);
  and _74287_ (_22791_, _22790_, _09107_);
  and _74288_ (_22792_, _22791_, _22788_);
  or _74289_ (_22793_, _22767_, _08404_);
  and _74290_ (_22796_, _22728_, _06509_);
  and _74291_ (_22797_, _22796_, _22793_);
  or _74292_ (_22798_, _22797_, _06602_);
  or _74293_ (_22799_, _22798_, _22792_);
  or _74294_ (_22800_, _22778_, _09112_);
  and _74295_ (_22801_, _22800_, _07048_);
  and _74296_ (_22802_, _22801_, _22799_);
  and _74297_ (_22803_, _22731_, _06639_);
  or _74298_ (_22804_, _22803_, _06646_);
  or _74299_ (_22805_, _22804_, _22802_);
  nor _74300_ (_22807_, _22733_, _06651_);
  nand _74301_ (_22808_, _22807_, _22730_);
  and _74302_ (_22809_, _22808_, _01442_);
  and _74303_ (_22810_, _22809_, _22805_);
  or _74304_ (_22811_, _22810_, _22727_);
  and _74305_ (_44173_, _22811_, _43634_);
  and _74306_ (_22812_, _01446_, \oc8051_golden_model_1.TL0 [2]);
  and _74307_ (_22813_, _11849_, \oc8051_golden_model_1.TL0 [2]);
  or _74308_ (_22814_, _22813_, _08503_);
  and _74309_ (_22815_, _08133_, _09057_);
  or _74310_ (_22817_, _22815_, _22813_);
  and _74311_ (_22818_, _22817_, _06507_);
  and _74312_ (_22819_, _22818_, _22814_);
  and _74313_ (_22820_, _09356_, _08133_);
  or _74314_ (_22821_, _22820_, _22813_);
  and _74315_ (_22822_, _22821_, _14025_);
  and _74316_ (_22823_, _14959_, _07976_);
  or _74317_ (_22824_, _22823_, _22813_);
  or _74318_ (_22825_, _22824_, _07275_);
  and _74319_ (_22826_, _08133_, \oc8051_golden_model_1.ACC [2]);
  or _74320_ (_22828_, _22826_, _22813_);
  and _74321_ (_22829_, _22828_, _07259_);
  and _74322_ (_22830_, _07260_, \oc8051_golden_model_1.TL0 [2]);
  or _74323_ (_22831_, _22830_, _06474_);
  or _74324_ (_22832_, _22831_, _22829_);
  and _74325_ (_22833_, _22832_, _06772_);
  and _74326_ (_22834_, _22833_, _22825_);
  nor _74327_ (_22835_, _11854_, _07854_);
  or _74328_ (_22836_, _22835_, _22813_);
  and _74329_ (_22837_, _22836_, _06410_);
  or _74330_ (_22839_, _22837_, _22834_);
  and _74331_ (_22840_, _22839_, _06426_);
  and _74332_ (_22841_, _22828_, _06417_);
  or _74333_ (_22842_, _22841_, _10153_);
  or _74334_ (_22843_, _22842_, _22840_);
  or _74335_ (_22844_, _22836_, _06327_);
  and _74336_ (_22845_, _22844_, _16672_);
  and _74337_ (_22846_, _22845_, _22843_);
  or _74338_ (_22847_, _22846_, _06037_);
  or _74339_ (_22848_, _22847_, _22822_);
  and _74340_ (_22850_, _15056_, _07976_);
  or _74341_ (_22851_, _22813_, _06313_);
  or _74342_ (_22852_, _22851_, _22850_);
  and _74343_ (_22853_, _22852_, _06278_);
  and _74344_ (_22854_, _22853_, _22848_);
  and _74345_ (_22855_, _22817_, _06277_);
  or _74346_ (_22856_, _22855_, _06502_);
  or _74347_ (_22857_, _22856_, _22854_);
  and _74348_ (_22858_, _14948_, _07976_);
  or _74349_ (_22859_, _22813_, _07334_);
  or _74350_ (_22861_, _22859_, _22858_);
  and _74351_ (_22862_, _22861_, _07337_);
  and _74352_ (_22863_, _22862_, _22857_);
  and _74353_ (_22864_, _10583_, _08133_);
  or _74354_ (_22865_, _22864_, _22813_);
  and _74355_ (_22866_, _22865_, _06615_);
  or _74356_ (_22867_, _22866_, _22863_);
  and _74357_ (_22868_, _22867_, _07339_);
  or _74358_ (_22869_, _22868_, _22819_);
  and _74359_ (_22870_, _22869_, _07331_);
  and _74360_ (_22872_, _22828_, _06610_);
  and _74361_ (_22873_, _22872_, _22814_);
  or _74362_ (_22874_, _22873_, _06509_);
  or _74363_ (_22875_, _22874_, _22870_);
  and _74364_ (_22876_, _14945_, _07976_);
  or _74365_ (_22877_, _22813_, _09107_);
  or _74366_ (_22878_, _22877_, _22876_);
  and _74367_ (_22879_, _22878_, _09112_);
  and _74368_ (_22880_, _22879_, _22875_);
  nor _74369_ (_22881_, _10582_, _11854_);
  or _74370_ (_22883_, _22881_, _22813_);
  and _74371_ (_22884_, _22883_, _06602_);
  or _74372_ (_22885_, _22884_, _22880_);
  and _74373_ (_22886_, _22885_, _07048_);
  and _74374_ (_22887_, _22824_, _06639_);
  or _74375_ (_22888_, _22887_, _06646_);
  or _74376_ (_22889_, _22888_, _22886_);
  and _74377_ (_22890_, _15129_, _07976_);
  or _74378_ (_22891_, _22813_, _06651_);
  or _74379_ (_22892_, _22891_, _22890_);
  and _74380_ (_22894_, _22892_, _01442_);
  and _74381_ (_22895_, _22894_, _22889_);
  or _74382_ (_22896_, _22895_, _22812_);
  and _74383_ (_44174_, _22896_, _43634_);
  and _74384_ (_22897_, _11849_, \oc8051_golden_model_1.TL0 [3]);
  or _74385_ (_22898_, _22897_, _08359_);
  and _74386_ (_22899_, _08133_, _09014_);
  or _74387_ (_22900_, _22899_, _22897_);
  and _74388_ (_22901_, _22900_, _06507_);
  and _74389_ (_22902_, _22901_, _22898_);
  nor _74390_ (_22904_, _10574_, _11854_);
  or _74391_ (_22905_, _22904_, _22897_);
  and _74392_ (_22906_, _08133_, \oc8051_golden_model_1.ACC [3]);
  nand _74393_ (_22907_, _22906_, _08359_);
  and _74394_ (_22908_, _22907_, _06615_);
  and _74395_ (_22909_, _22908_, _22905_);
  and _74396_ (_22910_, _15153_, _07976_);
  or _74397_ (_22911_, _22910_, _22897_);
  or _74398_ (_22912_, _22911_, _07275_);
  or _74399_ (_22913_, _22906_, _22897_);
  and _74400_ (_22915_, _22913_, _07259_);
  and _74401_ (_22916_, _07260_, \oc8051_golden_model_1.TL0 [3]);
  or _74402_ (_22917_, _22916_, _06474_);
  or _74403_ (_22918_, _22917_, _22915_);
  and _74404_ (_22919_, _22918_, _06772_);
  and _74405_ (_22920_, _22919_, _22912_);
  nor _74406_ (_22921_, _11854_, _07680_);
  or _74407_ (_22922_, _22921_, _22897_);
  and _74408_ (_22923_, _22922_, _06410_);
  or _74409_ (_22924_, _22923_, _22920_);
  and _74410_ (_22926_, _22924_, _06426_);
  and _74411_ (_22927_, _22913_, _06417_);
  or _74412_ (_22928_, _22927_, _10153_);
  or _74413_ (_22929_, _22928_, _22926_);
  or _74414_ (_22930_, _22922_, _06327_);
  and _74415_ (_22931_, _22930_, _22929_);
  or _74416_ (_22932_, _22931_, _09572_);
  and _74417_ (_22933_, _09310_, _08133_);
  or _74418_ (_22934_, _22897_, _06333_);
  or _74419_ (_22935_, _22934_, _22933_);
  and _74420_ (_22937_, _22935_, _06313_);
  and _74421_ (_22938_, _22937_, _22932_);
  and _74422_ (_22939_, _15251_, _08133_);
  or _74423_ (_22940_, _22939_, _22897_);
  and _74424_ (_22941_, _22940_, _06037_);
  or _74425_ (_22942_, _22941_, _06277_);
  or _74426_ (_22943_, _22942_, _22938_);
  or _74427_ (_22944_, _22900_, _06278_);
  and _74428_ (_22945_, _22944_, _22943_);
  or _74429_ (_22946_, _22945_, _06502_);
  and _74430_ (_22948_, _15266_, _07976_);
  or _74431_ (_22949_, _22897_, _07334_);
  or _74432_ (_22950_, _22949_, _22948_);
  and _74433_ (_22951_, _22950_, _07337_);
  and _74434_ (_22952_, _22951_, _22946_);
  or _74435_ (_22953_, _22952_, _22909_);
  and _74436_ (_22954_, _22953_, _07339_);
  or _74437_ (_22955_, _22954_, _22902_);
  and _74438_ (_22956_, _22955_, _07331_);
  and _74439_ (_22957_, _22913_, _06610_);
  and _74440_ (_22959_, _22957_, _22898_);
  or _74441_ (_22960_, _22959_, _06509_);
  or _74442_ (_22961_, _22960_, _22956_);
  and _74443_ (_22962_, _15263_, _07976_);
  or _74444_ (_22963_, _22897_, _09107_);
  or _74445_ (_22964_, _22963_, _22962_);
  and _74446_ (_22965_, _22964_, _09112_);
  and _74447_ (_22966_, _22965_, _22961_);
  and _74448_ (_22967_, _22905_, _06602_);
  or _74449_ (_22968_, _22967_, _06639_);
  or _74450_ (_22970_, _22968_, _22966_);
  or _74451_ (_22971_, _22911_, _07048_);
  and _74452_ (_22972_, _22971_, _06651_);
  and _74453_ (_22973_, _22972_, _22970_);
  and _74454_ (_22974_, _15321_, _07976_);
  or _74455_ (_22975_, _22974_, _22897_);
  and _74456_ (_22976_, _22975_, _06646_);
  or _74457_ (_22977_, _22976_, _01446_);
  or _74458_ (_22978_, _22977_, _22973_);
  or _74459_ (_22979_, _01442_, \oc8051_golden_model_1.TL0 [3]);
  and _74460_ (_22981_, _22979_, _43634_);
  and _74461_ (_44175_, _22981_, _22978_);
  and _74462_ (_22982_, _11849_, \oc8051_golden_model_1.TL0 [4]);
  or _74463_ (_22983_, _22982_, _08599_);
  and _74464_ (_22984_, _08995_, _08133_);
  or _74465_ (_22985_, _22984_, _22982_);
  and _74466_ (_22986_, _22985_, _06507_);
  and _74467_ (_22987_, _22986_, _22983_);
  nor _74468_ (_22988_, _10589_, _11854_);
  or _74469_ (_22989_, _22988_, _22982_);
  and _74470_ (_22991_, _08133_, \oc8051_golden_model_1.ACC [4]);
  nand _74471_ (_22992_, _22991_, _08599_);
  and _74472_ (_22993_, _22992_, _06615_);
  and _74473_ (_22994_, _22993_, _22989_);
  nor _74474_ (_22995_, _08596_, _11854_);
  or _74475_ (_22996_, _22995_, _22982_);
  or _74476_ (_22997_, _22996_, _06327_);
  and _74477_ (_22998_, _15367_, _07976_);
  or _74478_ (_22999_, _22998_, _22982_);
  or _74479_ (_23000_, _22999_, _07275_);
  or _74480_ (_23002_, _22991_, _22982_);
  and _74481_ (_23003_, _23002_, _07259_);
  and _74482_ (_23004_, _07260_, \oc8051_golden_model_1.TL0 [4]);
  or _74483_ (_23005_, _23004_, _06474_);
  or _74484_ (_23006_, _23005_, _23003_);
  and _74485_ (_23007_, _23006_, _06772_);
  and _74486_ (_23008_, _23007_, _23000_);
  and _74487_ (_23009_, _22996_, _06410_);
  or _74488_ (_23010_, _23009_, _23008_);
  and _74489_ (_23011_, _23010_, _06426_);
  and _74490_ (_23013_, _23002_, _06417_);
  or _74491_ (_23014_, _23013_, _10153_);
  or _74492_ (_23015_, _23014_, _23011_);
  and _74493_ (_23016_, _23015_, _22997_);
  or _74494_ (_23017_, _23016_, _09572_);
  and _74495_ (_23018_, _09264_, _07976_);
  or _74496_ (_23019_, _22982_, _16672_);
  or _74497_ (_23020_, _23019_, _23018_);
  and _74498_ (_23021_, _23020_, _23017_);
  or _74499_ (_23022_, _23021_, _06037_);
  and _74500_ (_23024_, _15452_, _07976_);
  or _74501_ (_23025_, _22982_, _06313_);
  or _74502_ (_23026_, _23025_, _23024_);
  and _74503_ (_23027_, _23026_, _06278_);
  and _74504_ (_23028_, _23027_, _23022_);
  and _74505_ (_23029_, _22985_, _06277_);
  or _74506_ (_23030_, _23029_, _06502_);
  or _74507_ (_23031_, _23030_, _23028_);
  and _74508_ (_23032_, _15345_, _07976_);
  or _74509_ (_23033_, _22982_, _07334_);
  or _74510_ (_23035_, _23033_, _23032_);
  and _74511_ (_23036_, _23035_, _07337_);
  and _74512_ (_23037_, _23036_, _23031_);
  or _74513_ (_23038_, _23037_, _22994_);
  and _74514_ (_23039_, _23038_, _07339_);
  or _74515_ (_23040_, _23039_, _22987_);
  and _74516_ (_23041_, _23040_, _07331_);
  and _74517_ (_23042_, _23002_, _06610_);
  and _74518_ (_23043_, _23042_, _22983_);
  or _74519_ (_23044_, _23043_, _06509_);
  or _74520_ (_23045_, _23044_, _23041_);
  and _74521_ (_23046_, _15342_, _07976_);
  or _74522_ (_23047_, _22982_, _09107_);
  or _74523_ (_23048_, _23047_, _23046_);
  and _74524_ (_23049_, _23048_, _09112_);
  and _74525_ (_23050_, _23049_, _23045_);
  and _74526_ (_23051_, _22989_, _06602_);
  or _74527_ (_23052_, _23051_, _06639_);
  or _74528_ (_23053_, _23052_, _23050_);
  or _74529_ (_23054_, _22999_, _07048_);
  and _74530_ (_23057_, _23054_, _06651_);
  and _74531_ (_23058_, _23057_, _23053_);
  and _74532_ (_23059_, _15524_, _07976_);
  or _74533_ (_23060_, _23059_, _22982_);
  and _74534_ (_23061_, _23060_, _06646_);
  or _74535_ (_23062_, _23061_, _01446_);
  or _74536_ (_23063_, _23062_, _23058_);
  or _74537_ (_23064_, _01442_, \oc8051_golden_model_1.TL0 [4]);
  and _74538_ (_23065_, _23064_, _43634_);
  and _74539_ (_44176_, _23065_, _23063_);
  and _74540_ (_23067_, _11849_, \oc8051_golden_model_1.TL0 [5]);
  nor _74541_ (_23068_, _10570_, _11854_);
  or _74542_ (_23069_, _23068_, _23067_);
  and _74543_ (_23070_, _08133_, \oc8051_golden_model_1.ACC [5]);
  nand _74544_ (_23071_, _23070_, _08308_);
  and _74545_ (_23072_, _23071_, _06615_);
  and _74546_ (_23073_, _23072_, _23069_);
  and _74547_ (_23074_, _15550_, _07976_);
  or _74548_ (_23075_, _23074_, _23067_);
  or _74549_ (_23076_, _23075_, _07275_);
  or _74550_ (_23078_, _23070_, _23067_);
  and _74551_ (_23079_, _23078_, _07259_);
  and _74552_ (_23080_, _07260_, \oc8051_golden_model_1.TL0 [5]);
  or _74553_ (_23081_, _23080_, _06474_);
  or _74554_ (_23082_, _23081_, _23079_);
  and _74555_ (_23083_, _23082_, _06772_);
  and _74556_ (_23084_, _23083_, _23076_);
  nor _74557_ (_23085_, _08305_, _11854_);
  or _74558_ (_23086_, _23085_, _23067_);
  and _74559_ (_23087_, _23086_, _06410_);
  or _74560_ (_23089_, _23087_, _23084_);
  and _74561_ (_23090_, _23089_, _06426_);
  and _74562_ (_23091_, _23078_, _06417_);
  or _74563_ (_23092_, _23091_, _10153_);
  or _74564_ (_23093_, _23092_, _23090_);
  or _74565_ (_23094_, _23086_, _06327_);
  and _74566_ (_23095_, _23094_, _23093_);
  or _74567_ (_23096_, _23095_, _09572_);
  and _74568_ (_23097_, _09218_, _08133_);
  or _74569_ (_23098_, _23067_, _06333_);
  or _74570_ (_23100_, _23098_, _23097_);
  and _74571_ (_23101_, _23100_, _06313_);
  and _74572_ (_23102_, _23101_, _23096_);
  and _74573_ (_23103_, _15649_, _08133_);
  or _74574_ (_23104_, _23103_, _23067_);
  and _74575_ (_23105_, _23104_, _06037_);
  or _74576_ (_23106_, _23105_, _06277_);
  or _74577_ (_23107_, _23106_, _23102_);
  and _74578_ (_23108_, _08954_, _08133_);
  or _74579_ (_23109_, _23108_, _23067_);
  or _74580_ (_23111_, _23109_, _06278_);
  and _74581_ (_23112_, _23111_, _23107_);
  or _74582_ (_23113_, _23112_, _06502_);
  and _74583_ (_23114_, _15664_, _07976_);
  or _74584_ (_23115_, _23067_, _07334_);
  or _74585_ (_23116_, _23115_, _23114_);
  and _74586_ (_23117_, _23116_, _07337_);
  and _74587_ (_23118_, _23117_, _23113_);
  or _74588_ (_23119_, _23118_, _23073_);
  and _74589_ (_23120_, _23119_, _07339_);
  or _74590_ (_23122_, _23067_, _08308_);
  and _74591_ (_23123_, _23109_, _06507_);
  and _74592_ (_23124_, _23123_, _23122_);
  or _74593_ (_23125_, _23124_, _23120_);
  and _74594_ (_23126_, _23125_, _07331_);
  and _74595_ (_23127_, _23078_, _06610_);
  and _74596_ (_23128_, _23127_, _23122_);
  or _74597_ (_23129_, _23128_, _06509_);
  or _74598_ (_23130_, _23129_, _23126_);
  and _74599_ (_23131_, _15663_, _07976_);
  or _74600_ (_23133_, _23067_, _09107_);
  or _74601_ (_23134_, _23133_, _23131_);
  and _74602_ (_23135_, _23134_, _09112_);
  and _74603_ (_23136_, _23135_, _23130_);
  and _74604_ (_23137_, _23069_, _06602_);
  or _74605_ (_23138_, _23137_, _06639_);
  or _74606_ (_23139_, _23138_, _23136_);
  or _74607_ (_23140_, _23075_, _07048_);
  and _74608_ (_23141_, _23140_, _06651_);
  and _74609_ (_23142_, _23141_, _23139_);
  and _74610_ (_23144_, _15721_, _07976_);
  or _74611_ (_23145_, _23144_, _23067_);
  and _74612_ (_23146_, _23145_, _06646_);
  or _74613_ (_23147_, _23146_, _01446_);
  or _74614_ (_23148_, _23147_, _23142_);
  or _74615_ (_23149_, _01442_, \oc8051_golden_model_1.TL0 [5]);
  and _74616_ (_23150_, _23149_, _43634_);
  and _74617_ (_44177_, _23150_, _23148_);
  and _74618_ (_23151_, _11849_, \oc8051_golden_model_1.TL0 [6]);
  nor _74619_ (_23152_, _08209_, _11854_);
  or _74620_ (_23154_, _23152_, _23151_);
  or _74621_ (_23155_, _23154_, _06327_);
  and _74622_ (_23156_, _15759_, _07976_);
  or _74623_ (_23157_, _23156_, _23151_);
  or _74624_ (_23158_, _23157_, _07275_);
  and _74625_ (_23159_, _08133_, \oc8051_golden_model_1.ACC [6]);
  or _74626_ (_23160_, _23159_, _23151_);
  and _74627_ (_23161_, _23160_, _07259_);
  and _74628_ (_23162_, _07260_, \oc8051_golden_model_1.TL0 [6]);
  or _74629_ (_23163_, _23162_, _06474_);
  or _74630_ (_23165_, _23163_, _23161_);
  and _74631_ (_23166_, _23165_, _06772_);
  and _74632_ (_23167_, _23166_, _23158_);
  and _74633_ (_23168_, _23154_, _06410_);
  or _74634_ (_23169_, _23168_, _23167_);
  and _74635_ (_23170_, _23169_, _06426_);
  and _74636_ (_23171_, _23160_, _06417_);
  or _74637_ (_23172_, _23171_, _10153_);
  or _74638_ (_23173_, _23172_, _23170_);
  and _74639_ (_23174_, _23173_, _23155_);
  or _74640_ (_23176_, _23174_, _09572_);
  and _74641_ (_23177_, _09172_, _08133_);
  or _74642_ (_23178_, _23151_, _06333_);
  or _74643_ (_23179_, _23178_, _23177_);
  and _74644_ (_23180_, _23179_, _06313_);
  and _74645_ (_23181_, _23180_, _23176_);
  and _74646_ (_23182_, _15846_, _08133_);
  or _74647_ (_23183_, _23182_, _23151_);
  and _74648_ (_23184_, _23183_, _06037_);
  or _74649_ (_23185_, _23184_, _06277_);
  or _74650_ (_23187_, _23185_, _23181_);
  and _74651_ (_23188_, _15853_, _08133_);
  or _74652_ (_23189_, _23188_, _23151_);
  or _74653_ (_23190_, _23189_, _06278_);
  and _74654_ (_23191_, _23190_, _23187_);
  or _74655_ (_23192_, _23191_, _06502_);
  and _74656_ (_23193_, _15862_, _07976_);
  or _74657_ (_23194_, _23151_, _07334_);
  or _74658_ (_23195_, _23194_, _23193_);
  and _74659_ (_23196_, _23195_, _07337_);
  and _74660_ (_23198_, _23196_, _23192_);
  and _74661_ (_23199_, _10596_, _08133_);
  or _74662_ (_23200_, _23199_, _23151_);
  and _74663_ (_23201_, _23200_, _06615_);
  or _74664_ (_23202_, _23201_, _23198_);
  and _74665_ (_23203_, _23202_, _07339_);
  or _74666_ (_23204_, _23151_, _08212_);
  and _74667_ (_23205_, _23189_, _06507_);
  and _74668_ (_23206_, _23205_, _23204_);
  or _74669_ (_23207_, _23206_, _23203_);
  and _74670_ (_23209_, _23207_, _07331_);
  and _74671_ (_23210_, _23160_, _06610_);
  and _74672_ (_23211_, _23210_, _23204_);
  or _74673_ (_23212_, _23211_, _06509_);
  or _74674_ (_23213_, _23212_, _23209_);
  and _74675_ (_23214_, _15859_, _07976_);
  or _74676_ (_23215_, _23151_, _09107_);
  or _74677_ (_23216_, _23215_, _23214_);
  and _74678_ (_23217_, _23216_, _09112_);
  and _74679_ (_23218_, _23217_, _23213_);
  nor _74680_ (_23220_, _10595_, _11854_);
  or _74681_ (_23221_, _23220_, _23151_);
  and _74682_ (_23222_, _23221_, _06602_);
  or _74683_ (_23223_, _23222_, _06639_);
  or _74684_ (_23224_, _23223_, _23218_);
  or _74685_ (_23225_, _23157_, _07048_);
  and _74686_ (_23226_, _23225_, _06651_);
  and _74687_ (_23227_, _23226_, _23224_);
  and _74688_ (_23228_, _15921_, _07976_);
  or _74689_ (_23229_, _23228_, _23151_);
  and _74690_ (_23231_, _23229_, _06646_);
  or _74691_ (_23232_, _23231_, _01446_);
  or _74692_ (_23233_, _23232_, _23227_);
  or _74693_ (_23234_, _01442_, \oc8051_golden_model_1.TL0 [6]);
  and _74694_ (_23235_, _23234_, _43634_);
  and _74695_ (_44178_, _23235_, _23233_);
  and _74696_ (_23236_, _01446_, \oc8051_golden_model_1.TCON [0]);
  and _74697_ (_23237_, _11929_, \oc8051_golden_model_1.TCON [0]);
  nor _74698_ (_23238_, _12622_, _11929_);
  or _74699_ (_23239_, _23238_, _23237_);
  and _74700_ (_23241_, _10577_, _08006_);
  nor _74701_ (_23242_, _23241_, _07337_);
  and _74702_ (_23243_, _23242_, _23239_);
  nor _74703_ (_23244_, _08453_, _11929_);
  or _74704_ (_23245_, _23244_, _23237_);
  or _74705_ (_23246_, _23245_, _07275_);
  and _74706_ (_23247_, _08006_, \oc8051_golden_model_1.ACC [0]);
  or _74707_ (_23248_, _23247_, _23237_);
  and _74708_ (_23249_, _23248_, _07259_);
  and _74709_ (_23250_, _07260_, \oc8051_golden_model_1.TCON [0]);
  or _74710_ (_23252_, _23250_, _06474_);
  or _74711_ (_23253_, _23252_, _23249_);
  and _74712_ (_23254_, _23253_, _06357_);
  and _74713_ (_23255_, _23254_, _23246_);
  and _74714_ (_23256_, _11937_, \oc8051_golden_model_1.TCON [0]);
  and _74715_ (_23257_, _14581_, _08633_);
  or _74716_ (_23258_, _23257_, _23256_);
  and _74717_ (_23259_, _23258_, _06356_);
  or _74718_ (_23260_, _23259_, _23255_);
  and _74719_ (_23261_, _23260_, _06772_);
  and _74720_ (_23263_, _08006_, _07250_);
  or _74721_ (_23264_, _23263_, _23237_);
  and _74722_ (_23265_, _23264_, _06410_);
  or _74723_ (_23266_, _23265_, _06417_);
  or _74724_ (_23267_, _23266_, _23261_);
  or _74725_ (_23268_, _23248_, _06426_);
  and _74726_ (_23269_, _23268_, _06353_);
  and _74727_ (_23270_, _23269_, _23267_);
  and _74728_ (_23271_, _23237_, _06352_);
  or _74729_ (_23272_, _23271_, _06345_);
  or _74730_ (_23274_, _23272_, _23270_);
  or _74731_ (_23275_, _23245_, _06346_);
  and _74732_ (_23276_, _23275_, _06340_);
  and _74733_ (_23277_, _23276_, _23274_);
  or _74734_ (_23278_, _23256_, _16663_);
  and _74735_ (_23279_, _23278_, _06339_);
  and _74736_ (_23280_, _23279_, _23258_);
  or _74737_ (_23281_, _23280_, _10153_);
  or _74738_ (_23282_, _23281_, _23277_);
  or _74739_ (_23283_, _23264_, _06327_);
  and _74740_ (_23285_, _23283_, _23282_);
  or _74741_ (_23286_, _23285_, _09572_);
  and _74742_ (_23287_, _09447_, _08006_);
  or _74743_ (_23288_, _23237_, _06333_);
  or _74744_ (_23289_, _23288_, _23287_);
  and _74745_ (_23290_, _23289_, _06313_);
  and _74746_ (_23291_, _23290_, _23286_);
  and _74747_ (_23292_, _14666_, _08006_);
  or _74748_ (_23293_, _23292_, _23237_);
  and _74749_ (_23294_, _23293_, _06037_);
  or _74750_ (_23296_, _23294_, _06277_);
  or _74751_ (_23297_, _23296_, _23291_);
  and _74752_ (_23298_, _08006_, _09008_);
  or _74753_ (_23299_, _23298_, _23237_);
  or _74754_ (_23300_, _23299_, _06278_);
  and _74755_ (_23301_, _23300_, _23297_);
  or _74756_ (_23302_, _23301_, _06502_);
  and _74757_ (_23303_, _14566_, _08006_);
  or _74758_ (_23304_, _23237_, _07334_);
  or _74759_ (_23305_, _23304_, _23303_);
  and _74760_ (_23307_, _23305_, _07337_);
  and _74761_ (_23308_, _23307_, _23302_);
  or _74762_ (_23309_, _23308_, _23243_);
  and _74763_ (_23310_, _23309_, _07339_);
  nand _74764_ (_23311_, _23299_, _06507_);
  nor _74765_ (_23312_, _23311_, _23244_);
  or _74766_ (_23313_, _23312_, _06610_);
  or _74767_ (_23314_, _23313_, _23310_);
  or _74768_ (_23315_, _23241_, _23237_);
  or _74769_ (_23316_, _23315_, _07331_);
  and _74770_ (_23318_, _23316_, _23314_);
  or _74771_ (_23319_, _23318_, _06509_);
  and _74772_ (_23320_, _14563_, _08006_);
  or _74773_ (_23321_, _23237_, _09107_);
  or _74774_ (_23322_, _23321_, _23320_);
  and _74775_ (_23323_, _23322_, _09112_);
  and _74776_ (_23324_, _23323_, _23319_);
  and _74777_ (_23325_, _23239_, _06602_);
  or _74778_ (_23326_, _23325_, _06639_);
  or _74779_ (_23327_, _23326_, _23324_);
  or _74780_ (_23328_, _23245_, _07048_);
  and _74781_ (_23329_, _23328_, _23327_);
  or _74782_ (_23330_, _23329_, _05989_);
  or _74783_ (_23331_, _23237_, _05990_);
  and _74784_ (_23332_, _23331_, _23330_);
  or _74785_ (_23333_, _23332_, _06646_);
  or _74786_ (_23334_, _23245_, _06651_);
  and _74787_ (_23335_, _23334_, _01442_);
  and _74788_ (_23336_, _23335_, _23333_);
  or _74789_ (_23337_, _23336_, _23236_);
  and _74790_ (_44180_, _23337_, _43634_);
  and _74791_ (_23340_, _01446_, \oc8051_golden_model_1.TCON [1]);
  and _74792_ (_23341_, _11929_, \oc8051_golden_model_1.TCON [1]);
  nor _74793_ (_23342_, _10578_, _11929_);
  or _74794_ (_23343_, _23342_, _23341_);
  or _74795_ (_23344_, _23343_, _09112_);
  nand _74796_ (_23345_, _08006_, _07160_);
  or _74797_ (_23346_, _08006_, \oc8051_golden_model_1.TCON [1]);
  and _74798_ (_23347_, _23346_, _06277_);
  and _74799_ (_23348_, _23347_, _23345_);
  or _74800_ (_23350_, _14851_, _11929_);
  and _74801_ (_23351_, _23346_, _06037_);
  and _74802_ (_23352_, _23351_, _23350_);
  nor _74803_ (_23353_, _11929_, _07448_);
  or _74804_ (_23354_, _23353_, _23341_);
  or _74805_ (_23355_, _23354_, _06772_);
  and _74806_ (_23356_, _14744_, _08006_);
  not _74807_ (_23357_, _23356_);
  and _74808_ (_23358_, _23357_, _23346_);
  or _74809_ (_23359_, _23358_, _07275_);
  and _74810_ (_23361_, _08006_, \oc8051_golden_model_1.ACC [1]);
  or _74811_ (_23362_, _23361_, _23341_);
  and _74812_ (_23363_, _23362_, _07259_);
  and _74813_ (_23364_, _07260_, \oc8051_golden_model_1.TCON [1]);
  or _74814_ (_23365_, _23364_, _06474_);
  or _74815_ (_23366_, _23365_, _23363_);
  and _74816_ (_23367_, _23366_, _06357_);
  and _74817_ (_23368_, _23367_, _23359_);
  and _74818_ (_23369_, _11937_, \oc8051_golden_model_1.TCON [1]);
  and _74819_ (_23370_, _14767_, _08633_);
  or _74820_ (_23372_, _23370_, _23369_);
  and _74821_ (_23373_, _23372_, _06356_);
  or _74822_ (_23374_, _23373_, _06410_);
  or _74823_ (_23375_, _23374_, _23368_);
  and _74824_ (_23376_, _23375_, _23355_);
  or _74825_ (_23377_, _23376_, _06417_);
  or _74826_ (_23378_, _23362_, _06426_);
  and _74827_ (_23379_, _23378_, _06353_);
  and _74828_ (_23380_, _23379_, _23377_);
  and _74829_ (_23381_, _14754_, _08633_);
  or _74830_ (_23383_, _23381_, _23369_);
  and _74831_ (_23384_, _23383_, _06352_);
  or _74832_ (_23385_, _23384_, _06345_);
  or _74833_ (_23386_, _23385_, _23380_);
  and _74834_ (_23387_, _23370_, _14782_);
  or _74835_ (_23388_, _23369_, _06346_);
  or _74836_ (_23389_, _23388_, _23387_);
  and _74837_ (_23390_, _23389_, _23386_);
  and _74838_ (_23391_, _23390_, _06340_);
  and _74839_ (_23392_, _14796_, _08633_);
  or _74840_ (_23394_, _23369_, _23392_);
  and _74841_ (_23395_, _23394_, _06339_);
  or _74842_ (_23396_, _23395_, _10153_);
  or _74843_ (_23397_, _23396_, _23391_);
  or _74844_ (_23398_, _23354_, _06327_);
  and _74845_ (_23399_, _23398_, _23397_);
  or _74846_ (_23400_, _23399_, _09572_);
  and _74847_ (_23401_, _09402_, _08006_);
  or _74848_ (_23402_, _23341_, _06333_);
  or _74849_ (_23403_, _23402_, _23401_);
  and _74850_ (_23405_, _23403_, _06313_);
  and _74851_ (_23406_, _23405_, _23400_);
  or _74852_ (_23407_, _23406_, _23352_);
  and _74853_ (_23408_, _23407_, _06278_);
  or _74854_ (_23409_, _23408_, _23348_);
  and _74855_ (_23410_, _23409_, _07334_);
  or _74856_ (_23411_, _14749_, _11929_);
  and _74857_ (_23412_, _23346_, _06502_);
  and _74858_ (_23413_, _23412_, _23411_);
  or _74859_ (_23414_, _23413_, _06615_);
  or _74860_ (_23416_, _23414_, _23410_);
  and _74861_ (_23417_, _10579_, _08006_);
  or _74862_ (_23418_, _23417_, _23341_);
  or _74863_ (_23419_, _23418_, _07337_);
  and _74864_ (_23420_, _23419_, _07339_);
  and _74865_ (_23421_, _23420_, _23416_);
  or _74866_ (_23422_, _14747_, _11929_);
  and _74867_ (_23423_, _23346_, _06507_);
  and _74868_ (_23424_, _23423_, _23422_);
  or _74869_ (_23425_, _23424_, _06610_);
  or _74870_ (_23427_, _23425_, _23421_);
  and _74871_ (_23428_, _23361_, _08404_);
  or _74872_ (_23429_, _23341_, _07331_);
  or _74873_ (_23430_, _23429_, _23428_);
  and _74874_ (_23431_, _23430_, _09107_);
  and _74875_ (_23432_, _23431_, _23427_);
  or _74876_ (_23433_, _23345_, _08404_);
  and _74877_ (_23434_, _23346_, _06509_);
  and _74878_ (_23435_, _23434_, _23433_);
  or _74879_ (_23436_, _23435_, _06602_);
  or _74880_ (_23438_, _23436_, _23432_);
  and _74881_ (_23439_, _23438_, _23344_);
  or _74882_ (_23440_, _23439_, _06639_);
  or _74883_ (_23441_, _23358_, _07048_);
  and _74884_ (_23442_, _23441_, _05990_);
  and _74885_ (_23443_, _23442_, _23440_);
  and _74886_ (_23444_, _23383_, _05989_);
  or _74887_ (_23445_, _23444_, _06646_);
  or _74888_ (_23446_, _23445_, _23443_);
  or _74889_ (_23447_, _23341_, _06651_);
  or _74890_ (_23449_, _23447_, _23356_);
  and _74891_ (_23450_, _23449_, _01442_);
  and _74892_ (_23451_, _23450_, _23446_);
  or _74893_ (_23452_, _23451_, _23340_);
  and _74894_ (_44181_, _23452_, _43634_);
  and _74895_ (_23453_, _01446_, \oc8051_golden_model_1.TCON [2]);
  and _74896_ (_23454_, _11929_, \oc8051_golden_model_1.TCON [2]);
  nor _74897_ (_23455_, _11929_, _07854_);
  or _74898_ (_23456_, _23455_, _23454_);
  or _74899_ (_23457_, _23456_, _06327_);
  or _74900_ (_23459_, _23456_, _06772_);
  and _74901_ (_23460_, _14959_, _08006_);
  or _74902_ (_23461_, _23460_, _23454_);
  or _74903_ (_23462_, _23461_, _07275_);
  and _74904_ (_23463_, _08006_, \oc8051_golden_model_1.ACC [2]);
  or _74905_ (_23464_, _23463_, _23454_);
  and _74906_ (_23465_, _23464_, _07259_);
  and _74907_ (_23466_, _07260_, \oc8051_golden_model_1.TCON [2]);
  or _74908_ (_23467_, _23466_, _06474_);
  or _74909_ (_23468_, _23467_, _23465_);
  and _74910_ (_23470_, _23468_, _06357_);
  and _74911_ (_23471_, _23470_, _23462_);
  and _74912_ (_23472_, _11937_, \oc8051_golden_model_1.TCON [2]);
  and _74913_ (_23473_, _14955_, _08633_);
  or _74914_ (_23474_, _23473_, _23472_);
  and _74915_ (_23475_, _23474_, _06356_);
  or _74916_ (_23476_, _23475_, _06410_);
  or _74917_ (_23477_, _23476_, _23471_);
  and _74918_ (_23478_, _23477_, _23459_);
  or _74919_ (_23479_, _23478_, _06417_);
  or _74920_ (_23481_, _23464_, _06426_);
  and _74921_ (_23482_, _23481_, _06353_);
  and _74922_ (_23483_, _23482_, _23479_);
  and _74923_ (_23484_, _14953_, _08633_);
  or _74924_ (_23485_, _23484_, _23472_);
  and _74925_ (_23486_, _23485_, _06352_);
  or _74926_ (_23487_, _23486_, _06345_);
  or _74927_ (_23488_, _23487_, _23483_);
  and _74928_ (_23489_, _23473_, _14986_);
  or _74929_ (_23490_, _23472_, _06346_);
  or _74930_ (_23492_, _23490_, _23489_);
  and _74931_ (_23493_, _23492_, _06340_);
  and _74932_ (_23494_, _23493_, _23488_);
  and _74933_ (_23495_, _15000_, _08633_);
  or _74934_ (_23496_, _23495_, _23472_);
  and _74935_ (_23497_, _23496_, _06339_);
  or _74936_ (_23498_, _23497_, _10153_);
  or _74937_ (_23499_, _23498_, _23494_);
  and _74938_ (_23500_, _23499_, _23457_);
  or _74939_ (_23501_, _23500_, _09572_);
  and _74940_ (_23503_, _09356_, _08006_);
  or _74941_ (_23504_, _23454_, _06333_);
  or _74942_ (_23505_, _23504_, _23503_);
  and _74943_ (_23506_, _23505_, _06313_);
  and _74944_ (_23507_, _23506_, _23501_);
  and _74945_ (_23508_, _15056_, _08006_);
  or _74946_ (_23509_, _23508_, _23454_);
  and _74947_ (_23510_, _23509_, _06037_);
  or _74948_ (_23511_, _23510_, _06277_);
  or _74949_ (_23512_, _23511_, _23507_);
  and _74950_ (_23514_, _08006_, _09057_);
  or _74951_ (_23515_, _23514_, _23454_);
  or _74952_ (_23516_, _23515_, _06278_);
  and _74953_ (_23517_, _23516_, _23512_);
  or _74954_ (_23518_, _23517_, _06502_);
  and _74955_ (_23519_, _14948_, _08006_);
  or _74956_ (_23520_, _23454_, _07334_);
  or _74957_ (_23521_, _23520_, _23519_);
  and _74958_ (_23522_, _23521_, _07337_);
  and _74959_ (_23523_, _23522_, _23518_);
  and _74960_ (_23525_, _10583_, _08006_);
  or _74961_ (_23526_, _23525_, _23454_);
  and _74962_ (_23527_, _23526_, _06615_);
  or _74963_ (_23528_, _23527_, _23523_);
  and _74964_ (_23529_, _23528_, _07339_);
  or _74965_ (_23530_, _23454_, _08503_);
  and _74966_ (_23531_, _23515_, _06507_);
  and _74967_ (_23532_, _23531_, _23530_);
  or _74968_ (_23533_, _23532_, _23529_);
  and _74969_ (_23534_, _23533_, _07331_);
  and _74970_ (_23536_, _23464_, _06610_);
  and _74971_ (_23537_, _23536_, _23530_);
  or _74972_ (_23538_, _23537_, _06509_);
  or _74973_ (_23539_, _23538_, _23534_);
  and _74974_ (_23540_, _14945_, _08006_);
  or _74975_ (_23541_, _23454_, _09107_);
  or _74976_ (_23542_, _23541_, _23540_);
  and _74977_ (_23543_, _23542_, _09112_);
  and _74978_ (_23544_, _23543_, _23539_);
  nor _74979_ (_23545_, _10582_, _11929_);
  or _74980_ (_23547_, _23545_, _23454_);
  and _74981_ (_23548_, _23547_, _06602_);
  or _74982_ (_23549_, _23548_, _06639_);
  or _74983_ (_23550_, _23549_, _23544_);
  or _74984_ (_23551_, _23461_, _07048_);
  and _74985_ (_23552_, _23551_, _05990_);
  and _74986_ (_23553_, _23552_, _23550_);
  and _74987_ (_23554_, _23485_, _05989_);
  or _74988_ (_23555_, _23554_, _06646_);
  or _74989_ (_23556_, _23555_, _23553_);
  and _74990_ (_23558_, _15129_, _08006_);
  or _74991_ (_23559_, _23454_, _06651_);
  or _74992_ (_23560_, _23559_, _23558_);
  and _74993_ (_23561_, _23560_, _01442_);
  and _74994_ (_23562_, _23561_, _23556_);
  or _74995_ (_23563_, _23562_, _23453_);
  and _74996_ (_44182_, _23563_, _43634_);
  and _74997_ (_23564_, _01446_, \oc8051_golden_model_1.TCON [3]);
  and _74998_ (_23565_, _11929_, \oc8051_golden_model_1.TCON [3]);
  nor _74999_ (_23566_, _11929_, _07680_);
  or _75000_ (_23568_, _23566_, _23565_);
  or _75001_ (_23569_, _23568_, _06327_);
  and _75002_ (_23570_, _15153_, _08006_);
  or _75003_ (_23571_, _23570_, _23565_);
  or _75004_ (_23572_, _23571_, _07275_);
  and _75005_ (_23573_, _08006_, \oc8051_golden_model_1.ACC [3]);
  or _75006_ (_23574_, _23573_, _23565_);
  and _75007_ (_23575_, _23574_, _07259_);
  and _75008_ (_23576_, _07260_, \oc8051_golden_model_1.TCON [3]);
  or _75009_ (_23577_, _23576_, _06474_);
  or _75010_ (_23579_, _23577_, _23575_);
  and _75011_ (_23580_, _23579_, _06357_);
  and _75012_ (_23581_, _23580_, _23572_);
  and _75013_ (_23582_, _11937_, \oc8051_golden_model_1.TCON [3]);
  and _75014_ (_23583_, _15150_, _08633_);
  or _75015_ (_23584_, _23583_, _23582_);
  and _75016_ (_23585_, _23584_, _06356_);
  or _75017_ (_23586_, _23585_, _06410_);
  or _75018_ (_23587_, _23586_, _23581_);
  or _75019_ (_23588_, _23568_, _06772_);
  and _75020_ (_23590_, _23588_, _23587_);
  or _75021_ (_23591_, _23590_, _06417_);
  or _75022_ (_23592_, _23574_, _06426_);
  and _75023_ (_23593_, _23592_, _06353_);
  and _75024_ (_23594_, _23593_, _23591_);
  and _75025_ (_23595_, _15148_, _08633_);
  or _75026_ (_23596_, _23595_, _23582_);
  and _75027_ (_23597_, _23596_, _06352_);
  or _75028_ (_23598_, _23597_, _06345_);
  or _75029_ (_23599_, _23598_, _23594_);
  or _75030_ (_23601_, _23582_, _15180_);
  and _75031_ (_23602_, _23601_, _23584_);
  or _75032_ (_23603_, _23602_, _06346_);
  and _75033_ (_23604_, _23603_, _06340_);
  and _75034_ (_23605_, _23604_, _23599_);
  and _75035_ (_23606_, _15197_, _08633_);
  or _75036_ (_23607_, _23606_, _23582_);
  and _75037_ (_23608_, _23607_, _06339_);
  or _75038_ (_23609_, _23608_, _10153_);
  or _75039_ (_23610_, _23609_, _23605_);
  and _75040_ (_23612_, _23610_, _23569_);
  or _75041_ (_23613_, _23612_, _09572_);
  and _75042_ (_23614_, _09310_, _08006_);
  or _75043_ (_23615_, _23565_, _06333_);
  or _75044_ (_23616_, _23615_, _23614_);
  and _75045_ (_23617_, _23616_, _06313_);
  and _75046_ (_23618_, _23617_, _23613_);
  and _75047_ (_23619_, _15251_, _08006_);
  or _75048_ (_23620_, _23619_, _23565_);
  and _75049_ (_23621_, _23620_, _06037_);
  or _75050_ (_23623_, _23621_, _06277_);
  or _75051_ (_23624_, _23623_, _23618_);
  and _75052_ (_23625_, _08006_, _09014_);
  or _75053_ (_23626_, _23625_, _23565_);
  or _75054_ (_23627_, _23626_, _06278_);
  and _75055_ (_23628_, _23627_, _23624_);
  or _75056_ (_23629_, _23628_, _06502_);
  and _75057_ (_23630_, _15266_, _08006_);
  or _75058_ (_23631_, _23565_, _07334_);
  or _75059_ (_23632_, _23631_, _23630_);
  and _75060_ (_23634_, _23632_, _07337_);
  and _75061_ (_23635_, _23634_, _23629_);
  and _75062_ (_23636_, _12619_, _08006_);
  or _75063_ (_23637_, _23636_, _23565_);
  and _75064_ (_23638_, _23637_, _06615_);
  or _75065_ (_23639_, _23638_, _23635_);
  and _75066_ (_23640_, _23639_, _07339_);
  or _75067_ (_23641_, _23565_, _08359_);
  and _75068_ (_23642_, _23626_, _06507_);
  and _75069_ (_23643_, _23642_, _23641_);
  or _75070_ (_23645_, _23643_, _23640_);
  and _75071_ (_23646_, _23645_, _07331_);
  and _75072_ (_23647_, _23574_, _06610_);
  and _75073_ (_23648_, _23647_, _23641_);
  or _75074_ (_23649_, _23648_, _06509_);
  or _75075_ (_23650_, _23649_, _23646_);
  and _75076_ (_23651_, _15263_, _08006_);
  or _75077_ (_23652_, _23565_, _09107_);
  or _75078_ (_23653_, _23652_, _23651_);
  and _75079_ (_23654_, _23653_, _09112_);
  and _75080_ (_23656_, _23654_, _23650_);
  nor _75081_ (_23657_, _10574_, _11929_);
  or _75082_ (_23658_, _23657_, _23565_);
  and _75083_ (_23659_, _23658_, _06602_);
  or _75084_ (_23660_, _23659_, _06639_);
  or _75085_ (_23661_, _23660_, _23656_);
  or _75086_ (_23662_, _23571_, _07048_);
  and _75087_ (_23663_, _23662_, _05990_);
  and _75088_ (_23664_, _23663_, _23661_);
  and _75089_ (_23665_, _23596_, _05989_);
  or _75090_ (_23667_, _23665_, _06646_);
  or _75091_ (_23668_, _23667_, _23664_);
  and _75092_ (_23669_, _15321_, _08006_);
  or _75093_ (_23670_, _23565_, _06651_);
  or _75094_ (_23671_, _23670_, _23669_);
  and _75095_ (_23672_, _23671_, _01442_);
  and _75096_ (_23673_, _23672_, _23668_);
  or _75097_ (_23674_, _23673_, _23564_);
  and _75098_ (_44184_, _23674_, _43634_);
  and _75099_ (_23675_, _01446_, \oc8051_golden_model_1.TCON [4]);
  and _75100_ (_23677_, _11929_, \oc8051_golden_model_1.TCON [4]);
  nor _75101_ (_23678_, _10589_, _11929_);
  or _75102_ (_23679_, _23678_, _23677_);
  and _75103_ (_23680_, _08006_, \oc8051_golden_model_1.ACC [4]);
  nand _75104_ (_23681_, _23680_, _08599_);
  and _75105_ (_23682_, _23681_, _06615_);
  and _75106_ (_23683_, _23682_, _23679_);
  nor _75107_ (_23684_, _08596_, _11929_);
  or _75108_ (_23685_, _23684_, _23677_);
  or _75109_ (_23686_, _23685_, _06327_);
  and _75110_ (_23688_, _11937_, \oc8051_golden_model_1.TCON [4]);
  and _75111_ (_23689_, _15348_, _08633_);
  or _75112_ (_23690_, _23689_, _23688_);
  and _75113_ (_23691_, _23690_, _06352_);
  and _75114_ (_23692_, _15367_, _08006_);
  or _75115_ (_23693_, _23692_, _23677_);
  or _75116_ (_23694_, _23693_, _07275_);
  or _75117_ (_23695_, _23680_, _23677_);
  and _75118_ (_23696_, _23695_, _07259_);
  and _75119_ (_23697_, _07260_, \oc8051_golden_model_1.TCON [4]);
  or _75120_ (_23699_, _23697_, _06474_);
  or _75121_ (_23700_, _23699_, _23696_);
  and _75122_ (_23701_, _23700_, _06357_);
  and _75123_ (_23702_, _23701_, _23694_);
  and _75124_ (_23703_, _15353_, _08633_);
  or _75125_ (_23704_, _23703_, _23688_);
  and _75126_ (_23705_, _23704_, _06356_);
  or _75127_ (_23706_, _23705_, _06410_);
  or _75128_ (_23707_, _23706_, _23702_);
  or _75129_ (_23708_, _23685_, _06772_);
  and _75130_ (_23710_, _23708_, _23707_);
  or _75131_ (_23711_, _23710_, _06417_);
  or _75132_ (_23712_, _23695_, _06426_);
  and _75133_ (_23713_, _23712_, _06353_);
  and _75134_ (_23714_, _23713_, _23711_);
  or _75135_ (_23715_, _23714_, _23691_);
  and _75136_ (_23716_, _23715_, _06346_);
  and _75137_ (_23717_, _15385_, _08633_);
  or _75138_ (_23718_, _23717_, _23688_);
  and _75139_ (_23719_, _23718_, _06345_);
  or _75140_ (_23721_, _23719_, _23716_);
  and _75141_ (_23722_, _23721_, _06340_);
  and _75142_ (_23723_, _15350_, _08633_);
  or _75143_ (_23724_, _23723_, _23688_);
  and _75144_ (_23725_, _23724_, _06339_);
  or _75145_ (_23726_, _23725_, _10153_);
  or _75146_ (_23727_, _23726_, _23722_);
  and _75147_ (_23728_, _23727_, _23686_);
  or _75148_ (_23729_, _23728_, _09572_);
  and _75149_ (_23730_, _09264_, _08006_);
  or _75150_ (_23732_, _23677_, _06333_);
  or _75151_ (_23733_, _23732_, _23730_);
  and _75152_ (_23734_, _23733_, _06313_);
  and _75153_ (_23735_, _23734_, _23729_);
  and _75154_ (_23736_, _15452_, _08006_);
  or _75155_ (_23737_, _23736_, _23677_);
  and _75156_ (_23738_, _23737_, _06037_);
  or _75157_ (_23739_, _23738_, _06277_);
  or _75158_ (_23740_, _23739_, _23735_);
  and _75159_ (_23741_, _08995_, _08006_);
  or _75160_ (_23743_, _23741_, _23677_);
  or _75161_ (_23744_, _23743_, _06278_);
  and _75162_ (_23745_, _23744_, _23740_);
  or _75163_ (_23746_, _23745_, _06502_);
  and _75164_ (_23747_, _15345_, _08006_);
  or _75165_ (_23748_, _23677_, _07334_);
  or _75166_ (_23749_, _23748_, _23747_);
  and _75167_ (_23750_, _23749_, _07337_);
  and _75168_ (_23751_, _23750_, _23746_);
  or _75169_ (_23752_, _23751_, _23683_);
  and _75170_ (_23754_, _23752_, _07339_);
  or _75171_ (_23755_, _23677_, _08599_);
  and _75172_ (_23756_, _23743_, _06507_);
  and _75173_ (_23757_, _23756_, _23755_);
  or _75174_ (_23758_, _23757_, _23754_);
  and _75175_ (_23759_, _23758_, _07331_);
  and _75176_ (_23760_, _23695_, _06610_);
  and _75177_ (_23761_, _23760_, _23755_);
  or _75178_ (_23762_, _23761_, _06509_);
  or _75179_ (_23763_, _23762_, _23759_);
  and _75180_ (_23764_, _15342_, _08006_);
  or _75181_ (_23765_, _23677_, _09107_);
  or _75182_ (_23766_, _23765_, _23764_);
  and _75183_ (_23767_, _23766_, _09112_);
  and _75184_ (_23768_, _23767_, _23763_);
  and _75185_ (_23769_, _23679_, _06602_);
  or _75186_ (_23770_, _23769_, _06639_);
  or _75187_ (_23771_, _23770_, _23768_);
  or _75188_ (_23772_, _23693_, _07048_);
  and _75189_ (_23773_, _23772_, _05990_);
  and _75190_ (_23776_, _23773_, _23771_);
  and _75191_ (_23777_, _23690_, _05989_);
  or _75192_ (_23778_, _23777_, _06646_);
  or _75193_ (_23779_, _23778_, _23776_);
  and _75194_ (_23780_, _15524_, _08006_);
  or _75195_ (_23781_, _23677_, _06651_);
  or _75196_ (_23782_, _23781_, _23780_);
  and _75197_ (_23783_, _23782_, _01442_);
  and _75198_ (_23784_, _23783_, _23779_);
  or _75199_ (_23785_, _23784_, _23675_);
  and _75200_ (_44185_, _23785_, _43634_);
  and _75201_ (_23787_, _01446_, \oc8051_golden_model_1.TCON [5]);
  and _75202_ (_23788_, _11929_, \oc8051_golden_model_1.TCON [5]);
  and _75203_ (_23789_, _15550_, _08006_);
  or _75204_ (_23790_, _23789_, _23788_);
  or _75205_ (_23791_, _23790_, _07275_);
  and _75206_ (_23792_, _08006_, \oc8051_golden_model_1.ACC [5]);
  or _75207_ (_23793_, _23792_, _23788_);
  and _75208_ (_23794_, _23793_, _07259_);
  and _75209_ (_23795_, _07260_, \oc8051_golden_model_1.TCON [5]);
  or _75210_ (_23797_, _23795_, _06474_);
  or _75211_ (_23798_, _23797_, _23794_);
  and _75212_ (_23799_, _23798_, _06357_);
  and _75213_ (_23800_, _23799_, _23791_);
  and _75214_ (_23801_, _11937_, \oc8051_golden_model_1.TCON [5]);
  and _75215_ (_23802_, _15566_, _08633_);
  or _75216_ (_23803_, _23802_, _23801_);
  and _75217_ (_23804_, _23803_, _06356_);
  or _75218_ (_23805_, _23804_, _06410_);
  or _75219_ (_23806_, _23805_, _23800_);
  nor _75220_ (_23808_, _08305_, _11929_);
  or _75221_ (_23809_, _23808_, _23788_);
  or _75222_ (_23810_, _23809_, _06772_);
  and _75223_ (_23811_, _23810_, _23806_);
  or _75224_ (_23812_, _23811_, _06417_);
  or _75225_ (_23813_, _23793_, _06426_);
  and _75226_ (_23814_, _23813_, _06353_);
  and _75227_ (_23815_, _23814_, _23812_);
  and _75228_ (_23816_, _15544_, _08633_);
  or _75229_ (_23817_, _23816_, _23801_);
  and _75230_ (_23819_, _23817_, _06352_);
  or _75231_ (_23820_, _23819_, _06345_);
  or _75232_ (_23821_, _23820_, _23815_);
  or _75233_ (_23822_, _23801_, _15581_);
  and _75234_ (_23823_, _23822_, _23803_);
  or _75235_ (_23824_, _23823_, _06346_);
  and _75236_ (_23825_, _23824_, _06340_);
  and _75237_ (_23826_, _23825_, _23821_);
  and _75238_ (_23827_, _15546_, _08633_);
  or _75239_ (_23828_, _23827_, _23801_);
  and _75240_ (_23830_, _23828_, _06339_);
  or _75241_ (_23831_, _23830_, _10153_);
  or _75242_ (_23832_, _23831_, _23826_);
  or _75243_ (_23833_, _23809_, _06327_);
  and _75244_ (_23834_, _23833_, _23832_);
  or _75245_ (_23835_, _23834_, _09572_);
  and _75246_ (_23836_, _09218_, _08006_);
  or _75247_ (_23837_, _23788_, _06333_);
  or _75248_ (_23838_, _23837_, _23836_);
  and _75249_ (_23839_, _23838_, _06313_);
  and _75250_ (_23841_, _23839_, _23835_);
  and _75251_ (_23842_, _15649_, _08006_);
  or _75252_ (_23843_, _23842_, _23788_);
  and _75253_ (_23844_, _23843_, _06037_);
  or _75254_ (_23845_, _23844_, _06277_);
  or _75255_ (_23846_, _23845_, _23841_);
  and _75256_ (_23847_, _08954_, _08006_);
  or _75257_ (_23848_, _23847_, _23788_);
  or _75258_ (_23849_, _23848_, _06278_);
  and _75259_ (_23850_, _23849_, _23846_);
  or _75260_ (_23852_, _23850_, _06502_);
  and _75261_ (_23853_, _15664_, _08006_);
  or _75262_ (_23854_, _23788_, _07334_);
  or _75263_ (_23855_, _23854_, _23853_);
  and _75264_ (_23856_, _23855_, _07337_);
  and _75265_ (_23857_, _23856_, _23852_);
  and _75266_ (_23858_, _12626_, _08006_);
  or _75267_ (_23859_, _23858_, _23788_);
  and _75268_ (_23860_, _23859_, _06615_);
  or _75269_ (_23861_, _23860_, _23857_);
  and _75270_ (_23863_, _23861_, _07339_);
  or _75271_ (_23864_, _23788_, _08308_);
  and _75272_ (_23865_, _23848_, _06507_);
  and _75273_ (_23866_, _23865_, _23864_);
  or _75274_ (_23867_, _23866_, _23863_);
  and _75275_ (_23868_, _23867_, _07331_);
  and _75276_ (_23869_, _23793_, _06610_);
  and _75277_ (_23870_, _23869_, _23864_);
  or _75278_ (_23871_, _23870_, _06509_);
  or _75279_ (_23872_, _23871_, _23868_);
  and _75280_ (_23874_, _15663_, _08006_);
  or _75281_ (_23875_, _23788_, _09107_);
  or _75282_ (_23876_, _23875_, _23874_);
  and _75283_ (_23877_, _23876_, _09112_);
  and _75284_ (_23878_, _23877_, _23872_);
  nor _75285_ (_23879_, _10570_, _11929_);
  or _75286_ (_23880_, _23879_, _23788_);
  and _75287_ (_23881_, _23880_, _06602_);
  or _75288_ (_23882_, _23881_, _06639_);
  or _75289_ (_23883_, _23882_, _23878_);
  or _75290_ (_23885_, _23790_, _07048_);
  and _75291_ (_23886_, _23885_, _05990_);
  and _75292_ (_23887_, _23886_, _23883_);
  and _75293_ (_23888_, _23817_, _05989_);
  or _75294_ (_23889_, _23888_, _06646_);
  or _75295_ (_23890_, _23889_, _23887_);
  and _75296_ (_23891_, _15721_, _08006_);
  or _75297_ (_23892_, _23788_, _06651_);
  or _75298_ (_23893_, _23892_, _23891_);
  and _75299_ (_23894_, _23893_, _01442_);
  and _75300_ (_23896_, _23894_, _23890_);
  or _75301_ (_23897_, _23896_, _23787_);
  and _75302_ (_44186_, _23897_, _43634_);
  and _75303_ (_23898_, _01446_, \oc8051_golden_model_1.TCON [6]);
  and _75304_ (_23899_, _11929_, \oc8051_golden_model_1.TCON [6]);
  nor _75305_ (_23900_, _10595_, _11929_);
  or _75306_ (_23901_, _23900_, _23899_);
  and _75307_ (_23902_, _08006_, \oc8051_golden_model_1.ACC [6]);
  nand _75308_ (_23903_, _23902_, _08212_);
  and _75309_ (_23904_, _23903_, _06615_);
  and _75310_ (_23906_, _23904_, _23901_);
  and _75311_ (_23907_, _15759_, _08006_);
  or _75312_ (_23908_, _23907_, _23899_);
  or _75313_ (_23909_, _23908_, _07275_);
  or _75314_ (_23910_, _23902_, _23899_);
  and _75315_ (_23911_, _23910_, _07259_);
  and _75316_ (_23912_, _07260_, \oc8051_golden_model_1.TCON [6]);
  or _75317_ (_23913_, _23912_, _06474_);
  or _75318_ (_23914_, _23913_, _23911_);
  and _75319_ (_23915_, _23914_, _06357_);
  and _75320_ (_23917_, _23915_, _23909_);
  and _75321_ (_23918_, _11937_, \oc8051_golden_model_1.TCON [6]);
  and _75322_ (_23919_, _15763_, _08633_);
  or _75323_ (_23920_, _23919_, _23918_);
  and _75324_ (_23921_, _23920_, _06356_);
  or _75325_ (_23922_, _23921_, _06410_);
  or _75326_ (_23923_, _23922_, _23917_);
  nor _75327_ (_23924_, _08209_, _11929_);
  or _75328_ (_23925_, _23924_, _23899_);
  or _75329_ (_23926_, _23925_, _06772_);
  and _75330_ (_23928_, _23926_, _23923_);
  or _75331_ (_23929_, _23928_, _06417_);
  or _75332_ (_23930_, _23910_, _06426_);
  and _75333_ (_23931_, _23930_, _06353_);
  and _75334_ (_23932_, _23931_, _23929_);
  and _75335_ (_23933_, _15743_, _08633_);
  or _75336_ (_23934_, _23933_, _23918_);
  and _75337_ (_23935_, _23934_, _06352_);
  or _75338_ (_23936_, _23935_, _06345_);
  or _75339_ (_23937_, _23936_, _23932_);
  or _75340_ (_23939_, _23918_, _15778_);
  and _75341_ (_23940_, _23939_, _23920_);
  or _75342_ (_23941_, _23940_, _06346_);
  and _75343_ (_23942_, _23941_, _06340_);
  and _75344_ (_23943_, _23942_, _23937_);
  and _75345_ (_23944_, _15745_, _08633_);
  or _75346_ (_23945_, _23944_, _23918_);
  and _75347_ (_23946_, _23945_, _06339_);
  or _75348_ (_23947_, _23946_, _10153_);
  or _75349_ (_23948_, _23947_, _23943_);
  or _75350_ (_23949_, _23925_, _06327_);
  and _75351_ (_23950_, _23949_, _23948_);
  or _75352_ (_23951_, _23950_, _09572_);
  and _75353_ (_23952_, _09172_, _08006_);
  or _75354_ (_23953_, _23899_, _06333_);
  or _75355_ (_23954_, _23953_, _23952_);
  and _75356_ (_23955_, _23954_, _06313_);
  and _75357_ (_23956_, _23955_, _23951_);
  and _75358_ (_23957_, _15846_, _08006_);
  or _75359_ (_23958_, _23957_, _23899_);
  and _75360_ (_23961_, _23958_, _06037_);
  or _75361_ (_23962_, _23961_, _06277_);
  or _75362_ (_23963_, _23962_, _23956_);
  and _75363_ (_23964_, _15853_, _08006_);
  or _75364_ (_23965_, _23964_, _23899_);
  or _75365_ (_23966_, _23965_, _06278_);
  and _75366_ (_23967_, _23966_, _23963_);
  or _75367_ (_23968_, _23967_, _06502_);
  and _75368_ (_23969_, _15862_, _08006_);
  or _75369_ (_23970_, _23899_, _07334_);
  or _75370_ (_23972_, _23970_, _23969_);
  and _75371_ (_23973_, _23972_, _07337_);
  and _75372_ (_23974_, _23973_, _23968_);
  or _75373_ (_23975_, _23974_, _23906_);
  and _75374_ (_23976_, _23975_, _07339_);
  or _75375_ (_23977_, _23899_, _08212_);
  and _75376_ (_23978_, _23965_, _06507_);
  and _75377_ (_23979_, _23978_, _23977_);
  or _75378_ (_23980_, _23979_, _23976_);
  and _75379_ (_23981_, _23980_, _07331_);
  and _75380_ (_23983_, _23910_, _06610_);
  and _75381_ (_23984_, _23983_, _23977_);
  or _75382_ (_23985_, _23984_, _06509_);
  or _75383_ (_23986_, _23985_, _23981_);
  and _75384_ (_23987_, _15859_, _08006_);
  or _75385_ (_23988_, _23899_, _09107_);
  or _75386_ (_23989_, _23988_, _23987_);
  and _75387_ (_23990_, _23989_, _09112_);
  and _75388_ (_23991_, _23990_, _23986_);
  and _75389_ (_23992_, _23901_, _06602_);
  or _75390_ (_23994_, _23992_, _06639_);
  or _75391_ (_23995_, _23994_, _23991_);
  or _75392_ (_23996_, _23908_, _07048_);
  and _75393_ (_23997_, _23996_, _05990_);
  and _75394_ (_23998_, _23997_, _23995_);
  and _75395_ (_23999_, _23934_, _05989_);
  or _75396_ (_24000_, _23999_, _06646_);
  or _75397_ (_24001_, _24000_, _23998_);
  and _75398_ (_24002_, _15921_, _08006_);
  or _75399_ (_24003_, _23899_, _06651_);
  or _75400_ (_24005_, _24003_, _24002_);
  and _75401_ (_24006_, _24005_, _01442_);
  and _75402_ (_24007_, _24006_, _24001_);
  or _75403_ (_24008_, _24007_, _23898_);
  and _75404_ (_44187_, _24008_, _43634_);
  and _75405_ (_24009_, _01446_, \oc8051_golden_model_1.TH1 [0]);
  and _75406_ (_24010_, _12031_, \oc8051_golden_model_1.TH1 [0]);
  nor _75407_ (_24011_, _12622_, _12031_);
  or _75408_ (_24012_, _24011_, _24010_);
  and _75409_ (_24013_, _10577_, _07981_);
  nor _75410_ (_24015_, _24013_, _07337_);
  and _75411_ (_24016_, _24015_, _24012_);
  and _75412_ (_24017_, _07981_, _07250_);
  or _75413_ (_24018_, _24017_, _24010_);
  or _75414_ (_24019_, _24018_, _06327_);
  nor _75415_ (_24020_, _08453_, _12031_);
  or _75416_ (_24021_, _24020_, _24010_);
  or _75417_ (_24022_, _24021_, _07275_);
  and _75418_ (_24023_, _07981_, \oc8051_golden_model_1.ACC [0]);
  or _75419_ (_24024_, _24023_, _24010_);
  and _75420_ (_24026_, _24024_, _07259_);
  and _75421_ (_24027_, _07260_, \oc8051_golden_model_1.TH1 [0]);
  or _75422_ (_24028_, _24027_, _06474_);
  or _75423_ (_24029_, _24028_, _24026_);
  and _75424_ (_24030_, _24029_, _06772_);
  and _75425_ (_24031_, _24030_, _24022_);
  and _75426_ (_24032_, _24018_, _06410_);
  or _75427_ (_24033_, _24032_, _24031_);
  and _75428_ (_24034_, _24033_, _06426_);
  and _75429_ (_24035_, _24024_, _06417_);
  or _75430_ (_24037_, _24035_, _10153_);
  or _75431_ (_24038_, _24037_, _24034_);
  and _75432_ (_24039_, _24038_, _24019_);
  or _75433_ (_24040_, _24039_, _09572_);
  and _75434_ (_24041_, _09447_, _07981_);
  or _75435_ (_24042_, _24010_, _06333_);
  or _75436_ (_24043_, _24042_, _24041_);
  and _75437_ (_24044_, _24043_, _24040_);
  or _75438_ (_24045_, _24044_, _06037_);
  and _75439_ (_24046_, _14666_, _07981_);
  or _75440_ (_24048_, _24010_, _06313_);
  or _75441_ (_24049_, _24048_, _24046_);
  and _75442_ (_24050_, _24049_, _06278_);
  and _75443_ (_24051_, _24050_, _24045_);
  and _75444_ (_24052_, _07981_, _09008_);
  or _75445_ (_24053_, _24052_, _24010_);
  and _75446_ (_24054_, _24053_, _06277_);
  or _75447_ (_24055_, _24054_, _06502_);
  or _75448_ (_24056_, _24055_, _24051_);
  and _75449_ (_24057_, _14566_, _07981_);
  or _75450_ (_24059_, _24010_, _07334_);
  or _75451_ (_24060_, _24059_, _24057_);
  and _75452_ (_24061_, _24060_, _07337_);
  and _75453_ (_24062_, _24061_, _24056_);
  or _75454_ (_24063_, _24062_, _24016_);
  and _75455_ (_24064_, _24063_, _07339_);
  nand _75456_ (_24065_, _24053_, _06507_);
  nor _75457_ (_24066_, _24065_, _24020_);
  or _75458_ (_24067_, _24066_, _06610_);
  or _75459_ (_24068_, _24067_, _24064_);
  or _75460_ (_24070_, _24013_, _24010_);
  or _75461_ (_24071_, _24070_, _07331_);
  and _75462_ (_24072_, _24071_, _24068_);
  or _75463_ (_24073_, _24072_, _06509_);
  and _75464_ (_24074_, _14563_, _07981_);
  or _75465_ (_24075_, _24010_, _09107_);
  or _75466_ (_24076_, _24075_, _24074_);
  and _75467_ (_24077_, _24076_, _09112_);
  and _75468_ (_24078_, _24077_, _24073_);
  and _75469_ (_24079_, _24012_, _06602_);
  or _75470_ (_24081_, _24079_, _19642_);
  or _75471_ (_24082_, _24081_, _24078_);
  or _75472_ (_24083_, _24021_, _19641_);
  and _75473_ (_24084_, _24083_, _01442_);
  and _75474_ (_24085_, _24084_, _24082_);
  or _75475_ (_24086_, _24085_, _24009_);
  and _75476_ (_44189_, _24086_, _43634_);
  not _75477_ (_24087_, \oc8051_golden_model_1.TH1 [1]);
  nor _75478_ (_24088_, _01442_, _24087_);
  nand _75479_ (_24089_, _07981_, _07160_);
  or _75480_ (_24091_, _07981_, \oc8051_golden_model_1.TH1 [1]);
  and _75481_ (_24092_, _24091_, _06277_);
  and _75482_ (_24093_, _24092_, _24089_);
  nor _75483_ (_24094_, _12031_, _07448_);
  nor _75484_ (_24095_, _07981_, _24087_);
  or _75485_ (_24096_, _24095_, _19597_);
  or _75486_ (_24097_, _24096_, _24094_);
  and _75487_ (_24098_, _07981_, \oc8051_golden_model_1.ACC [1]);
  or _75488_ (_24099_, _24098_, _24095_);
  and _75489_ (_24100_, _24099_, _06417_);
  or _75490_ (_24102_, _24100_, _10153_);
  and _75491_ (_24103_, _14744_, _07981_);
  not _75492_ (_24104_, _24103_);
  and _75493_ (_24105_, _24104_, _24091_);
  and _75494_ (_24106_, _24105_, _06474_);
  nor _75495_ (_24107_, _07259_, _24087_);
  and _75496_ (_24108_, _24099_, _07259_);
  or _75497_ (_24109_, _24108_, _24107_);
  and _75498_ (_24110_, _24109_, _07275_);
  or _75499_ (_24111_, _24110_, _06410_);
  or _75500_ (_24113_, _24111_, _24106_);
  and _75501_ (_24114_, _24113_, _06426_);
  or _75502_ (_24115_, _24114_, _24102_);
  and _75503_ (_24116_, _24115_, _24097_);
  or _75504_ (_24117_, _24116_, _09572_);
  and _75505_ (_24118_, _24117_, _06313_);
  and _75506_ (_24119_, _09402_, _07981_);
  or _75507_ (_24120_, _24095_, _06333_);
  or _75508_ (_24121_, _24120_, _24119_);
  and _75509_ (_24122_, _24121_, _24118_);
  or _75510_ (_24124_, _14851_, _12031_);
  and _75511_ (_24125_, _24091_, _06037_);
  and _75512_ (_24126_, _24125_, _24124_);
  or _75513_ (_24127_, _24126_, _24122_);
  and _75514_ (_24128_, _24127_, _06278_);
  or _75515_ (_24129_, _24128_, _24093_);
  and _75516_ (_24130_, _24129_, _07334_);
  or _75517_ (_24131_, _14749_, _12031_);
  and _75518_ (_24132_, _24091_, _06502_);
  and _75519_ (_24133_, _24132_, _24131_);
  or _75520_ (_24135_, _24133_, _06615_);
  or _75521_ (_24136_, _24135_, _24130_);
  nor _75522_ (_24137_, _10578_, _12031_);
  or _75523_ (_24138_, _24137_, _24095_);
  nand _75524_ (_24139_, _10576_, _07981_);
  and _75525_ (_24140_, _24139_, _24138_);
  or _75526_ (_24141_, _24140_, _07337_);
  and _75527_ (_24142_, _24141_, _07339_);
  and _75528_ (_24143_, _24142_, _24136_);
  or _75529_ (_24144_, _14747_, _12031_);
  and _75530_ (_24146_, _24091_, _06507_);
  and _75531_ (_24147_, _24146_, _24144_);
  or _75532_ (_24148_, _24147_, _06610_);
  or _75533_ (_24149_, _24148_, _24143_);
  nor _75534_ (_24150_, _24095_, _07331_);
  nand _75535_ (_24151_, _24150_, _24139_);
  and _75536_ (_24152_, _24151_, _09107_);
  and _75537_ (_24153_, _24152_, _24149_);
  or _75538_ (_24154_, _24089_, _08404_);
  and _75539_ (_24155_, _24091_, _06509_);
  and _75540_ (_24157_, _24155_, _24154_);
  or _75541_ (_24158_, _24157_, _06602_);
  or _75542_ (_24159_, _24158_, _24153_);
  or _75543_ (_24160_, _24138_, _09112_);
  and _75544_ (_24161_, _24160_, _07048_);
  and _75545_ (_24162_, _24161_, _24159_);
  and _75546_ (_24163_, _24105_, _06639_);
  or _75547_ (_24164_, _24163_, _06646_);
  or _75548_ (_24165_, _24164_, _24162_);
  or _75549_ (_24166_, _24095_, _06651_);
  or _75550_ (_24168_, _24166_, _24103_);
  and _75551_ (_24169_, _24168_, _01442_);
  and _75552_ (_24170_, _24169_, _24165_);
  or _75553_ (_24171_, _24170_, _24088_);
  and _75554_ (_44190_, _24171_, _43634_);
  and _75555_ (_24172_, _01446_, \oc8051_golden_model_1.TH1 [2]);
  and _75556_ (_24173_, _12031_, \oc8051_golden_model_1.TH1 [2]);
  and _75557_ (_24174_, _09356_, _07981_);
  or _75558_ (_24175_, _24174_, _24173_);
  and _75559_ (_24176_, _24175_, _14025_);
  and _75560_ (_24178_, _14959_, _07981_);
  or _75561_ (_24179_, _24178_, _24173_);
  or _75562_ (_24180_, _24179_, _07275_);
  and _75563_ (_24181_, _07981_, \oc8051_golden_model_1.ACC [2]);
  or _75564_ (_24182_, _24181_, _24173_);
  and _75565_ (_24183_, _24182_, _07259_);
  and _75566_ (_24184_, _07260_, \oc8051_golden_model_1.TH1 [2]);
  or _75567_ (_24185_, _24184_, _06474_);
  or _75568_ (_24186_, _24185_, _24183_);
  and _75569_ (_24187_, _24186_, _06772_);
  and _75570_ (_24189_, _24187_, _24180_);
  nor _75571_ (_24190_, _12031_, _07854_);
  or _75572_ (_24191_, _24190_, _24173_);
  and _75573_ (_24192_, _24191_, _06410_);
  or _75574_ (_24193_, _24192_, _24189_);
  and _75575_ (_24194_, _24193_, _06426_);
  and _75576_ (_24195_, _24182_, _06417_);
  or _75577_ (_24196_, _24195_, _10153_);
  or _75578_ (_24197_, _24196_, _24194_);
  or _75579_ (_24198_, _24191_, _06327_);
  and _75580_ (_24200_, _24198_, _16672_);
  and _75581_ (_24201_, _24200_, _24197_);
  or _75582_ (_24202_, _24201_, _06037_);
  or _75583_ (_24203_, _24202_, _24176_);
  and _75584_ (_24204_, _15056_, _07981_);
  or _75585_ (_24205_, _24173_, _06313_);
  or _75586_ (_24206_, _24205_, _24204_);
  and _75587_ (_24207_, _24206_, _06278_);
  and _75588_ (_24208_, _24207_, _24203_);
  and _75589_ (_24209_, _07981_, _09057_);
  or _75590_ (_24211_, _24209_, _24173_);
  and _75591_ (_24212_, _24211_, _06277_);
  or _75592_ (_24213_, _24212_, _06502_);
  or _75593_ (_24214_, _24213_, _24208_);
  and _75594_ (_24215_, _14948_, _07981_);
  or _75595_ (_24216_, _24173_, _07334_);
  or _75596_ (_24217_, _24216_, _24215_);
  and _75597_ (_24218_, _24217_, _07337_);
  and _75598_ (_24219_, _24218_, _24214_);
  and _75599_ (_24220_, _10583_, _07981_);
  or _75600_ (_24222_, _24220_, _24173_);
  and _75601_ (_24223_, _24222_, _06615_);
  or _75602_ (_24224_, _24223_, _24219_);
  and _75603_ (_24225_, _24224_, _07339_);
  or _75604_ (_24226_, _24173_, _08503_);
  and _75605_ (_24227_, _24211_, _06507_);
  and _75606_ (_24228_, _24227_, _24226_);
  or _75607_ (_24229_, _24228_, _24225_);
  and _75608_ (_24230_, _24229_, _07331_);
  and _75609_ (_24231_, _24182_, _06610_);
  and _75610_ (_24233_, _24231_, _24226_);
  or _75611_ (_24234_, _24233_, _06509_);
  or _75612_ (_24235_, _24234_, _24230_);
  and _75613_ (_24236_, _14945_, _07981_);
  or _75614_ (_24237_, _24173_, _09107_);
  or _75615_ (_24238_, _24237_, _24236_);
  and _75616_ (_24239_, _24238_, _09112_);
  and _75617_ (_24240_, _24239_, _24235_);
  nor _75618_ (_24241_, _10582_, _12031_);
  or _75619_ (_24242_, _24241_, _24173_);
  and _75620_ (_24244_, _24242_, _06602_);
  or _75621_ (_24245_, _24244_, _24240_);
  and _75622_ (_24246_, _24245_, _07048_);
  and _75623_ (_24247_, _24179_, _06639_);
  or _75624_ (_24248_, _24247_, _06646_);
  or _75625_ (_24249_, _24248_, _24246_);
  and _75626_ (_24250_, _15129_, _07981_);
  or _75627_ (_24251_, _24173_, _06651_);
  or _75628_ (_24252_, _24251_, _24250_);
  and _75629_ (_24253_, _24252_, _01442_);
  and _75630_ (_24256_, _24253_, _24249_);
  or _75631_ (_24257_, _24256_, _24172_);
  and _75632_ (_44191_, _24257_, _43634_);
  and _75633_ (_24258_, _12031_, \oc8051_golden_model_1.TH1 [3]);
  or _75634_ (_24259_, _24258_, _08359_);
  and _75635_ (_24260_, _07981_, _09014_);
  or _75636_ (_24261_, _24260_, _24258_);
  and _75637_ (_24262_, _24261_, _06507_);
  and _75638_ (_24263_, _24262_, _24259_);
  and _75639_ (_24264_, _15153_, _07981_);
  or _75640_ (_24266_, _24264_, _24258_);
  or _75641_ (_24267_, _24266_, _07275_);
  and _75642_ (_24268_, _07981_, \oc8051_golden_model_1.ACC [3]);
  or _75643_ (_24269_, _24268_, _24258_);
  and _75644_ (_24270_, _24269_, _07259_);
  and _75645_ (_24271_, _07260_, \oc8051_golden_model_1.TH1 [3]);
  or _75646_ (_24272_, _24271_, _06474_);
  or _75647_ (_24273_, _24272_, _24270_);
  and _75648_ (_24274_, _24273_, _06772_);
  and _75649_ (_24275_, _24274_, _24267_);
  nor _75650_ (_24277_, _12031_, _07680_);
  or _75651_ (_24278_, _24277_, _24258_);
  and _75652_ (_24279_, _24278_, _06410_);
  or _75653_ (_24280_, _24279_, _24275_);
  and _75654_ (_24281_, _24280_, _06426_);
  and _75655_ (_24282_, _24269_, _06417_);
  or _75656_ (_24283_, _24282_, _10153_);
  or _75657_ (_24284_, _24283_, _24281_);
  or _75658_ (_24285_, _24278_, _06327_);
  and _75659_ (_24286_, _24285_, _24284_);
  or _75660_ (_24287_, _24286_, _09572_);
  and _75661_ (_24288_, _09310_, _07981_);
  or _75662_ (_24289_, _24258_, _06333_);
  or _75663_ (_24290_, _24289_, _24288_);
  and _75664_ (_24291_, _24290_, _06313_);
  and _75665_ (_24292_, _24291_, _24287_);
  and _75666_ (_24293_, _15251_, _07981_);
  or _75667_ (_24294_, _24293_, _24258_);
  and _75668_ (_24295_, _24294_, _06037_);
  or _75669_ (_24296_, _24295_, _06277_);
  or _75670_ (_24298_, _24296_, _24292_);
  or _75671_ (_24299_, _24261_, _06278_);
  and _75672_ (_24300_, _24299_, _24298_);
  or _75673_ (_24301_, _24300_, _06502_);
  and _75674_ (_24302_, _15266_, _07981_);
  or _75675_ (_24303_, _24258_, _07334_);
  or _75676_ (_24304_, _24303_, _24302_);
  and _75677_ (_24305_, _24304_, _07337_);
  and _75678_ (_24306_, _24305_, _24301_);
  and _75679_ (_24307_, _12619_, _07981_);
  or _75680_ (_24309_, _24307_, _24258_);
  and _75681_ (_24310_, _24309_, _06615_);
  or _75682_ (_24311_, _24310_, _24306_);
  and _75683_ (_24312_, _24311_, _07339_);
  or _75684_ (_24313_, _24312_, _24263_);
  and _75685_ (_24314_, _24313_, _07331_);
  and _75686_ (_24315_, _24269_, _06610_);
  and _75687_ (_24316_, _24315_, _24259_);
  or _75688_ (_24317_, _24316_, _06509_);
  or _75689_ (_24318_, _24317_, _24314_);
  and _75690_ (_24320_, _15263_, _07981_);
  or _75691_ (_24321_, _24258_, _09107_);
  or _75692_ (_24322_, _24321_, _24320_);
  and _75693_ (_24323_, _24322_, _09112_);
  and _75694_ (_24324_, _24323_, _24318_);
  nor _75695_ (_24325_, _10574_, _12031_);
  or _75696_ (_24326_, _24325_, _24258_);
  and _75697_ (_24327_, _24326_, _06602_);
  or _75698_ (_24328_, _24327_, _06639_);
  or _75699_ (_24329_, _24328_, _24324_);
  or _75700_ (_24330_, _24266_, _07048_);
  and _75701_ (_24331_, _24330_, _06651_);
  and _75702_ (_24332_, _24331_, _24329_);
  and _75703_ (_24333_, _15321_, _07981_);
  or _75704_ (_24334_, _24333_, _24258_);
  and _75705_ (_24335_, _24334_, _06646_);
  or _75706_ (_24336_, _24335_, _01446_);
  or _75707_ (_24337_, _24336_, _24332_);
  or _75708_ (_24338_, _01442_, \oc8051_golden_model_1.TH1 [3]);
  and _75709_ (_24339_, _24338_, _43634_);
  and _75710_ (_44192_, _24339_, _24337_);
  and _75711_ (_24341_, _12031_, \oc8051_golden_model_1.TH1 [4]);
  or _75712_ (_24342_, _24341_, _08599_);
  and _75713_ (_24343_, _08995_, _07981_);
  or _75714_ (_24344_, _24343_, _24341_);
  and _75715_ (_24345_, _24344_, _06507_);
  and _75716_ (_24346_, _24345_, _24342_);
  and _75717_ (_24347_, _15367_, _07981_);
  or _75718_ (_24348_, _24347_, _24341_);
  or _75719_ (_24349_, _24348_, _07275_);
  and _75720_ (_24350_, _07981_, \oc8051_golden_model_1.ACC [4]);
  or _75721_ (_24351_, _24350_, _24341_);
  and _75722_ (_24352_, _24351_, _07259_);
  and _75723_ (_24353_, _07260_, \oc8051_golden_model_1.TH1 [4]);
  or _75724_ (_24354_, _24353_, _06474_);
  or _75725_ (_24355_, _24354_, _24352_);
  and _75726_ (_24356_, _24355_, _06772_);
  and _75727_ (_24357_, _24356_, _24349_);
  nor _75728_ (_24358_, _08596_, _12031_);
  or _75729_ (_24359_, _24358_, _24341_);
  and _75730_ (_24361_, _24359_, _06410_);
  or _75731_ (_24362_, _24361_, _24357_);
  and _75732_ (_24363_, _24362_, _06426_);
  and _75733_ (_24364_, _24351_, _06417_);
  or _75734_ (_24365_, _24364_, _10153_);
  or _75735_ (_24366_, _24365_, _24363_);
  or _75736_ (_24367_, _24359_, _06327_);
  and _75737_ (_24368_, _24367_, _24366_);
  or _75738_ (_24369_, _24368_, _09572_);
  and _75739_ (_24370_, _09264_, _07981_);
  or _75740_ (_24372_, _24341_, _16672_);
  or _75741_ (_24373_, _24372_, _24370_);
  and _75742_ (_24374_, _24373_, _24369_);
  or _75743_ (_24375_, _24374_, _06037_);
  and _75744_ (_24376_, _15452_, _07981_);
  or _75745_ (_24377_, _24341_, _06313_);
  or _75746_ (_24378_, _24377_, _24376_);
  and _75747_ (_24379_, _24378_, _06278_);
  and _75748_ (_24380_, _24379_, _24375_);
  and _75749_ (_24381_, _24344_, _06277_);
  or _75750_ (_24382_, _24381_, _06502_);
  or _75751_ (_24383_, _24382_, _24380_);
  and _75752_ (_24384_, _15345_, _07981_);
  or _75753_ (_24385_, _24341_, _07334_);
  or _75754_ (_24386_, _24385_, _24384_);
  and _75755_ (_24387_, _24386_, _07337_);
  and _75756_ (_24388_, _24387_, _24383_);
  and _75757_ (_24389_, _10590_, _07981_);
  or _75758_ (_24390_, _24389_, _24341_);
  and _75759_ (_24391_, _24390_, _06615_);
  or _75760_ (_24393_, _24391_, _24388_);
  and _75761_ (_24394_, _24393_, _07339_);
  or _75762_ (_24395_, _24394_, _24346_);
  and _75763_ (_24396_, _24395_, _07331_);
  and _75764_ (_24397_, _24351_, _06610_);
  and _75765_ (_24398_, _24397_, _24342_);
  or _75766_ (_24399_, _24398_, _06509_);
  or _75767_ (_24400_, _24399_, _24396_);
  and _75768_ (_24401_, _15342_, _07981_);
  or _75769_ (_24402_, _24341_, _09107_);
  or _75770_ (_24404_, _24402_, _24401_);
  and _75771_ (_24405_, _24404_, _09112_);
  and _75772_ (_24406_, _24405_, _24400_);
  nor _75773_ (_24407_, _10589_, _12031_);
  or _75774_ (_24408_, _24407_, _24341_);
  and _75775_ (_24409_, _24408_, _06602_);
  or _75776_ (_24410_, _24409_, _06639_);
  or _75777_ (_24411_, _24410_, _24406_);
  or _75778_ (_24412_, _24348_, _07048_);
  and _75779_ (_24413_, _24412_, _06651_);
  and _75780_ (_24414_, _24413_, _24411_);
  and _75781_ (_24415_, _15524_, _07981_);
  or _75782_ (_24416_, _24415_, _24341_);
  and _75783_ (_24417_, _24416_, _06646_);
  or _75784_ (_24418_, _24417_, _01446_);
  or _75785_ (_24419_, _24418_, _24414_);
  or _75786_ (_24420_, _01442_, \oc8051_golden_model_1.TH1 [4]);
  and _75787_ (_24421_, _24420_, _43634_);
  and _75788_ (_44193_, _24421_, _24419_);
  and _75789_ (_24422_, _12031_, \oc8051_golden_model_1.TH1 [5]);
  nor _75790_ (_24424_, _10570_, _12031_);
  or _75791_ (_24425_, _24424_, _24422_);
  and _75792_ (_24426_, _07981_, \oc8051_golden_model_1.ACC [5]);
  nand _75793_ (_24427_, _24426_, _08308_);
  and _75794_ (_24428_, _24427_, _06615_);
  and _75795_ (_24429_, _24428_, _24425_);
  nor _75796_ (_24430_, _08305_, _12031_);
  or _75797_ (_24431_, _24430_, _24422_);
  or _75798_ (_24432_, _24431_, _06327_);
  and _75799_ (_24433_, _15550_, _07981_);
  or _75800_ (_24435_, _24433_, _24422_);
  or _75801_ (_24436_, _24435_, _07275_);
  or _75802_ (_24437_, _24426_, _24422_);
  and _75803_ (_24438_, _24437_, _07259_);
  and _75804_ (_24439_, _07260_, \oc8051_golden_model_1.TH1 [5]);
  or _75805_ (_24440_, _24439_, _06474_);
  or _75806_ (_24441_, _24440_, _24438_);
  and _75807_ (_24442_, _24441_, _06772_);
  and _75808_ (_24443_, _24442_, _24436_);
  and _75809_ (_24444_, _24431_, _06410_);
  or _75810_ (_24445_, _24444_, _24443_);
  and _75811_ (_24446_, _24445_, _06426_);
  and _75812_ (_24447_, _24437_, _06417_);
  or _75813_ (_24448_, _24447_, _10153_);
  or _75814_ (_24449_, _24448_, _24446_);
  and _75815_ (_24450_, _24449_, _24432_);
  or _75816_ (_24451_, _24450_, _09572_);
  and _75817_ (_24452_, _09218_, _07981_);
  or _75818_ (_24453_, _24422_, _06333_);
  or _75819_ (_24454_, _24453_, _24452_);
  and _75820_ (_24456_, _24454_, _06313_);
  and _75821_ (_24457_, _24456_, _24451_);
  and _75822_ (_24458_, _15649_, _07981_);
  or _75823_ (_24459_, _24458_, _24422_);
  and _75824_ (_24460_, _24459_, _06037_);
  or _75825_ (_24461_, _24460_, _06277_);
  or _75826_ (_24462_, _24461_, _24457_);
  and _75827_ (_24463_, _08954_, _07981_);
  or _75828_ (_24464_, _24463_, _24422_);
  or _75829_ (_24465_, _24464_, _06278_);
  and _75830_ (_24467_, _24465_, _24462_);
  or _75831_ (_24468_, _24467_, _06502_);
  and _75832_ (_24469_, _15664_, _07981_);
  or _75833_ (_24470_, _24422_, _07334_);
  or _75834_ (_24471_, _24470_, _24469_);
  and _75835_ (_24472_, _24471_, _07337_);
  and _75836_ (_24473_, _24472_, _24468_);
  or _75837_ (_24474_, _24473_, _24429_);
  and _75838_ (_24475_, _24474_, _07339_);
  or _75839_ (_24476_, _24422_, _08308_);
  and _75840_ (_24477_, _24464_, _06507_);
  and _75841_ (_24478_, _24477_, _24476_);
  or _75842_ (_24479_, _24478_, _24475_);
  and _75843_ (_24480_, _24479_, _07331_);
  and _75844_ (_24481_, _24437_, _06610_);
  and _75845_ (_24482_, _24481_, _24476_);
  or _75846_ (_24483_, _24482_, _06509_);
  or _75847_ (_24484_, _24483_, _24480_);
  and _75848_ (_24485_, _15663_, _07981_);
  or _75849_ (_24486_, _24422_, _09107_);
  or _75850_ (_24488_, _24486_, _24485_);
  and _75851_ (_24489_, _24488_, _09112_);
  and _75852_ (_24490_, _24489_, _24484_);
  and _75853_ (_24491_, _24425_, _06602_);
  or _75854_ (_24492_, _24491_, _06639_);
  or _75855_ (_24493_, _24492_, _24490_);
  or _75856_ (_24494_, _24435_, _07048_);
  and _75857_ (_24495_, _24494_, _06651_);
  and _75858_ (_24496_, _24495_, _24493_);
  and _75859_ (_24497_, _15721_, _07981_);
  or _75860_ (_24499_, _24497_, _24422_);
  and _75861_ (_24500_, _24499_, _06646_);
  or _75862_ (_24501_, _24500_, _01446_);
  or _75863_ (_24502_, _24501_, _24496_);
  or _75864_ (_24503_, _01442_, \oc8051_golden_model_1.TH1 [5]);
  and _75865_ (_24504_, _24503_, _43634_);
  and _75866_ (_44194_, _24504_, _24502_);
  and _75867_ (_24505_, _12031_, \oc8051_golden_model_1.TH1 [6]);
  and _75868_ (_24506_, _15759_, _07981_);
  or _75869_ (_24507_, _24506_, _24505_);
  or _75870_ (_24508_, _24507_, _07275_);
  and _75871_ (_24509_, _07981_, \oc8051_golden_model_1.ACC [6]);
  or _75872_ (_24510_, _24509_, _24505_);
  and _75873_ (_24511_, _24510_, _07259_);
  and _75874_ (_24512_, _07260_, \oc8051_golden_model_1.TH1 [6]);
  or _75875_ (_24513_, _24512_, _06474_);
  or _75876_ (_24514_, _24513_, _24511_);
  and _75877_ (_24515_, _24514_, _06772_);
  and _75878_ (_24516_, _24515_, _24508_);
  nor _75879_ (_24517_, _08209_, _12031_);
  or _75880_ (_24519_, _24517_, _24505_);
  and _75881_ (_24520_, _24519_, _06410_);
  or _75882_ (_24521_, _24520_, _24516_);
  and _75883_ (_24522_, _24521_, _06426_);
  and _75884_ (_24523_, _24510_, _06417_);
  or _75885_ (_24524_, _24523_, _10153_);
  or _75886_ (_24525_, _24524_, _24522_);
  or _75887_ (_24526_, _24519_, _06327_);
  and _75888_ (_24527_, _24526_, _24525_);
  or _75889_ (_24528_, _24527_, _09572_);
  and _75890_ (_24530_, _09172_, _07981_);
  or _75891_ (_24531_, _24505_, _06333_);
  or _75892_ (_24532_, _24531_, _24530_);
  and _75893_ (_24533_, _24532_, _06313_);
  and _75894_ (_24534_, _24533_, _24528_);
  and _75895_ (_24535_, _15846_, _07981_);
  or _75896_ (_24536_, _24535_, _24505_);
  and _75897_ (_24537_, _24536_, _06037_);
  or _75898_ (_24538_, _24537_, _06277_);
  or _75899_ (_24539_, _24538_, _24534_);
  and _75900_ (_24540_, _15853_, _07981_);
  or _75901_ (_24541_, _24540_, _24505_);
  or _75902_ (_24542_, _24541_, _06278_);
  and _75903_ (_24543_, _24542_, _24539_);
  or _75904_ (_24544_, _24543_, _06502_);
  and _75905_ (_24545_, _15862_, _07981_);
  or _75906_ (_24546_, _24505_, _07334_);
  or _75907_ (_24547_, _24546_, _24545_);
  and _75908_ (_24548_, _24547_, _07337_);
  and _75909_ (_24549_, _24548_, _24544_);
  and _75910_ (_24551_, _10596_, _07981_);
  or _75911_ (_24552_, _24551_, _24505_);
  and _75912_ (_24553_, _24552_, _06615_);
  or _75913_ (_24554_, _24553_, _24549_);
  and _75914_ (_24555_, _24554_, _07339_);
  or _75915_ (_24556_, _24505_, _08212_);
  and _75916_ (_24557_, _24541_, _06507_);
  and _75917_ (_24558_, _24557_, _24556_);
  or _75918_ (_24559_, _24558_, _24555_);
  and _75919_ (_24560_, _24559_, _07331_);
  and _75920_ (_24562_, _24510_, _06610_);
  and _75921_ (_24563_, _24562_, _24556_);
  or _75922_ (_24564_, _24563_, _06509_);
  or _75923_ (_24565_, _24564_, _24560_);
  and _75924_ (_24566_, _15859_, _07981_);
  or _75925_ (_24567_, _24505_, _09107_);
  or _75926_ (_24568_, _24567_, _24566_);
  and _75927_ (_24569_, _24568_, _09112_);
  and _75928_ (_24570_, _24569_, _24565_);
  nor _75929_ (_24571_, _10595_, _12031_);
  or _75930_ (_24572_, _24571_, _24505_);
  and _75931_ (_24573_, _24572_, _06602_);
  or _75932_ (_24574_, _24573_, _06639_);
  or _75933_ (_24575_, _24574_, _24570_);
  or _75934_ (_24576_, _24507_, _07048_);
  and _75935_ (_24577_, _24576_, _06651_);
  and _75936_ (_24578_, _24577_, _24575_);
  and _75937_ (_24579_, _15921_, _07981_);
  or _75938_ (_24580_, _24579_, _24505_);
  and _75939_ (_24581_, _24580_, _06646_);
  or _75940_ (_24583_, _24581_, _01446_);
  or _75941_ (_24584_, _24583_, _24578_);
  or _75942_ (_24585_, _01442_, \oc8051_golden_model_1.TH1 [6]);
  and _75943_ (_24586_, _24585_, _43634_);
  and _75944_ (_44195_, _24586_, _24584_);
  and _75945_ (_24587_, _01446_, \oc8051_golden_model_1.TH0 [0]);
  and _75946_ (_24588_, _12109_, \oc8051_golden_model_1.TH0 [0]);
  and _75947_ (_24589_, _07954_, _07250_);
  or _75948_ (_24590_, _24589_, _24588_);
  or _75949_ (_24591_, _24590_, _06327_);
  nor _75950_ (_24593_, _08453_, _12109_);
  or _75951_ (_24594_, _24593_, _24588_);
  or _75952_ (_24595_, _24594_, _07275_);
  and _75953_ (_24596_, _07954_, \oc8051_golden_model_1.ACC [0]);
  or _75954_ (_24597_, _24596_, _24588_);
  and _75955_ (_24598_, _24597_, _07259_);
  and _75956_ (_24599_, _07260_, \oc8051_golden_model_1.TH0 [0]);
  or _75957_ (_24600_, _24599_, _06474_);
  or _75958_ (_24601_, _24600_, _24598_);
  and _75959_ (_24602_, _24601_, _06772_);
  and _75960_ (_24603_, _24602_, _24595_);
  and _75961_ (_24604_, _24590_, _06410_);
  or _75962_ (_24605_, _24604_, _24603_);
  and _75963_ (_24606_, _24605_, _06426_);
  and _75964_ (_24607_, _24597_, _06417_);
  or _75965_ (_24608_, _24607_, _10153_);
  or _75966_ (_24609_, _24608_, _24606_);
  and _75967_ (_24610_, _24609_, _24591_);
  or _75968_ (_24611_, _24610_, _09572_);
  and _75969_ (_24612_, _09447_, _07954_);
  or _75970_ (_24614_, _24588_, _06333_);
  or _75971_ (_24615_, _24614_, _24612_);
  and _75972_ (_24616_, _24615_, _24611_);
  or _75973_ (_24617_, _24616_, _06037_);
  and _75974_ (_24618_, _14666_, _07954_);
  or _75975_ (_24619_, _24588_, _06313_);
  or _75976_ (_24620_, _24619_, _24618_);
  and _75977_ (_24621_, _24620_, _06278_);
  and _75978_ (_24622_, _24621_, _24617_);
  and _75979_ (_24623_, _07954_, _09008_);
  or _75980_ (_24625_, _24623_, _24588_);
  and _75981_ (_24626_, _24625_, _06277_);
  or _75982_ (_24627_, _24626_, _06502_);
  or _75983_ (_24628_, _24627_, _24622_);
  and _75984_ (_24629_, _14566_, _07954_);
  or _75985_ (_24630_, _24588_, _07334_);
  or _75986_ (_24631_, _24630_, _24629_);
  and _75987_ (_24632_, _24631_, _07337_);
  and _75988_ (_24633_, _24632_, _24628_);
  nor _75989_ (_24634_, _12622_, _12109_);
  or _75990_ (_24635_, _24634_, _24588_);
  and _75991_ (_24636_, _10577_, _07954_);
  nor _75992_ (_24637_, _24636_, _07337_);
  and _75993_ (_24638_, _24637_, _24635_);
  or _75994_ (_24639_, _24638_, _24633_);
  and _75995_ (_24640_, _24639_, _07339_);
  nand _75996_ (_24641_, _24625_, _06507_);
  nor _75997_ (_24642_, _24641_, _24593_);
  or _75998_ (_24643_, _24642_, _06610_);
  or _75999_ (_24644_, _24643_, _24640_);
  or _76000_ (_24646_, _24636_, _24588_);
  or _76001_ (_24647_, _24646_, _07331_);
  and _76002_ (_24648_, _24647_, _24644_);
  or _76003_ (_24649_, _24648_, _06509_);
  and _76004_ (_24650_, _14563_, _07954_);
  or _76005_ (_24651_, _24588_, _09107_);
  or _76006_ (_24652_, _24651_, _24650_);
  and _76007_ (_24653_, _24652_, _09112_);
  and _76008_ (_24654_, _24653_, _24649_);
  and _76009_ (_24655_, _24635_, _06602_);
  or _76010_ (_24657_, _24655_, _19642_);
  or _76011_ (_24658_, _24657_, _24654_);
  or _76012_ (_24659_, _24594_, _19641_);
  and _76013_ (_24660_, _24659_, _01442_);
  and _76014_ (_24661_, _24660_, _24658_);
  or _76015_ (_24662_, _24661_, _24587_);
  and _76016_ (_44197_, _24662_, _43634_);
  and _76017_ (_24663_, _12109_, \oc8051_golden_model_1.TH0 [1]);
  nor _76018_ (_24664_, _10578_, _12109_);
  or _76019_ (_24665_, _24664_, _24663_);
  or _76020_ (_24666_, _24665_, _09112_);
  or _76021_ (_24667_, _07954_, \oc8051_golden_model_1.TH0 [1]);
  and _76022_ (_24668_, _14744_, _07954_);
  not _76023_ (_24669_, _24668_);
  and _76024_ (_24670_, _24669_, _24667_);
  or _76025_ (_24671_, _24670_, _07275_);
  and _76026_ (_24672_, _07954_, \oc8051_golden_model_1.ACC [1]);
  or _76027_ (_24673_, _24672_, _24663_);
  and _76028_ (_24674_, _24673_, _07259_);
  and _76029_ (_24675_, _07260_, \oc8051_golden_model_1.TH0 [1]);
  or _76030_ (_24677_, _24675_, _06474_);
  or _76031_ (_24678_, _24677_, _24674_);
  and _76032_ (_24679_, _24678_, _06772_);
  and _76033_ (_24680_, _24679_, _24671_);
  nor _76034_ (_24681_, _12109_, _07448_);
  or _76035_ (_24682_, _24681_, _24663_);
  and _76036_ (_24683_, _24682_, _06410_);
  or _76037_ (_24684_, _24683_, _24680_);
  and _76038_ (_24685_, _24684_, _06426_);
  and _76039_ (_24686_, _24673_, _06417_);
  or _76040_ (_24688_, _24686_, _10153_);
  or _76041_ (_24689_, _24688_, _24685_);
  or _76042_ (_24690_, _24682_, _06327_);
  and _76043_ (_24691_, _24690_, _16672_);
  and _76044_ (_24692_, _24691_, _24689_);
  or _76045_ (_24693_, _09402_, _12109_);
  and _76046_ (_24694_, _24667_, _14025_);
  and _76047_ (_24695_, _24694_, _24693_);
  or _76048_ (_24696_, _24695_, _24692_);
  and _76049_ (_24697_, _24696_, _06313_);
  or _76050_ (_24699_, _14851_, _12109_);
  and _76051_ (_24700_, _24667_, _06037_);
  and _76052_ (_24701_, _24700_, _24699_);
  or _76053_ (_24702_, _24701_, _24697_);
  and _76054_ (_24703_, _24702_, _06278_);
  nand _76055_ (_24704_, _07954_, _07160_);
  and _76056_ (_24705_, _24667_, _06277_);
  and _76057_ (_24706_, _24705_, _24704_);
  or _76058_ (_24707_, _24706_, _24703_);
  and _76059_ (_24708_, _24707_, _07334_);
  or _76060_ (_24709_, _14749_, _12109_);
  and _76061_ (_24710_, _24667_, _06502_);
  and _76062_ (_24711_, _24710_, _24709_);
  or _76063_ (_24712_, _24711_, _06615_);
  or _76064_ (_24713_, _24712_, _24708_);
  nand _76065_ (_24714_, _10576_, _07954_);
  and _76066_ (_24715_, _24714_, _24665_);
  or _76067_ (_24716_, _24715_, _07337_);
  and _76068_ (_24717_, _24716_, _07339_);
  and _76069_ (_24718_, _24717_, _24713_);
  or _76070_ (_24720_, _14747_, _12109_);
  and _76071_ (_24721_, _24667_, _06507_);
  and _76072_ (_24722_, _24721_, _24720_);
  or _76073_ (_24723_, _24722_, _06610_);
  or _76074_ (_24724_, _24723_, _24718_);
  nor _76075_ (_24725_, _24663_, _07331_);
  nand _76076_ (_24726_, _24725_, _24714_);
  and _76077_ (_24727_, _24726_, _09107_);
  and _76078_ (_24728_, _24727_, _24724_);
  or _76079_ (_24729_, _24704_, _08404_);
  and _76080_ (_24731_, _24667_, _06509_);
  and _76081_ (_24732_, _24731_, _24729_);
  or _76082_ (_24733_, _24732_, _06602_);
  or _76083_ (_24734_, _24733_, _24728_);
  and _76084_ (_24735_, _24734_, _24666_);
  or _76085_ (_24736_, _24735_, _06639_);
  or _76086_ (_24737_, _24670_, _07048_);
  and _76087_ (_24738_, _24737_, _06651_);
  and _76088_ (_24739_, _24738_, _24736_);
  or _76089_ (_24740_, _24668_, _24663_);
  and _76090_ (_24741_, _24740_, _06646_);
  or _76091_ (_24742_, _24741_, _01446_);
  or _76092_ (_24743_, _24742_, _24739_);
  or _76093_ (_24744_, _01442_, \oc8051_golden_model_1.TH0 [1]);
  and _76094_ (_24745_, _24744_, _43634_);
  and _76095_ (_44198_, _24745_, _24743_);
  and _76096_ (_24746_, _01446_, \oc8051_golden_model_1.TH0 [2]);
  and _76097_ (_24747_, _12109_, \oc8051_golden_model_1.TH0 [2]);
  nor _76098_ (_24748_, _10582_, _12109_);
  or _76099_ (_24749_, _24748_, _24747_);
  and _76100_ (_24751_, _07954_, \oc8051_golden_model_1.ACC [2]);
  nand _76101_ (_24752_, _24751_, _08503_);
  and _76102_ (_24753_, _24752_, _06615_);
  and _76103_ (_24754_, _24753_, _24749_);
  and _76104_ (_24755_, _09356_, _07954_);
  or _76105_ (_24756_, _24755_, _24747_);
  and _76106_ (_24757_, _24756_, _14025_);
  and _76107_ (_24758_, _14959_, _07954_);
  or _76108_ (_24759_, _24758_, _24747_);
  or _76109_ (_24760_, _24759_, _07275_);
  or _76110_ (_24762_, _24751_, _24747_);
  and _76111_ (_24763_, _24762_, _07259_);
  and _76112_ (_24764_, _07260_, \oc8051_golden_model_1.TH0 [2]);
  or _76113_ (_24765_, _24764_, _06474_);
  or _76114_ (_24766_, _24765_, _24763_);
  and _76115_ (_24767_, _24766_, _06772_);
  and _76116_ (_24768_, _24767_, _24760_);
  nor _76117_ (_24769_, _12109_, _07854_);
  or _76118_ (_24770_, _24769_, _24747_);
  and _76119_ (_24771_, _24770_, _06410_);
  or _76120_ (_24773_, _24771_, _24768_);
  and _76121_ (_24774_, _24773_, _06426_);
  and _76122_ (_24775_, _24762_, _06417_);
  or _76123_ (_24776_, _24775_, _10153_);
  or _76124_ (_24777_, _24776_, _24774_);
  or _76125_ (_24778_, _24770_, _06327_);
  and _76126_ (_24779_, _24778_, _16672_);
  and _76127_ (_24780_, _24779_, _24777_);
  or _76128_ (_24781_, _24780_, _06037_);
  or _76129_ (_24782_, _24781_, _24757_);
  and _76130_ (_24783_, _15056_, _07954_);
  or _76131_ (_24784_, _24747_, _06313_);
  or _76132_ (_24785_, _24784_, _24783_);
  and _76133_ (_24786_, _24785_, _06278_);
  and _76134_ (_24787_, _24786_, _24782_);
  and _76135_ (_24788_, _07954_, _09057_);
  or _76136_ (_24789_, _24788_, _24747_);
  and _76137_ (_24790_, _24789_, _06277_);
  or _76138_ (_24791_, _24790_, _06502_);
  or _76139_ (_24792_, _24791_, _24787_);
  and _76140_ (_24794_, _14948_, _07954_);
  or _76141_ (_24795_, _24747_, _07334_);
  or _76142_ (_24796_, _24795_, _24794_);
  and _76143_ (_24797_, _24796_, _07337_);
  and _76144_ (_24798_, _24797_, _24792_);
  or _76145_ (_24799_, _24798_, _24754_);
  and _76146_ (_24800_, _24799_, _07339_);
  or _76147_ (_24801_, _24747_, _08503_);
  and _76148_ (_24802_, _24789_, _06507_);
  and _76149_ (_24803_, _24802_, _24801_);
  or _76150_ (_24805_, _24803_, _24800_);
  and _76151_ (_24806_, _24805_, _07331_);
  and _76152_ (_24807_, _24762_, _06610_);
  and _76153_ (_24808_, _24807_, _24801_);
  or _76154_ (_24809_, _24808_, _06509_);
  or _76155_ (_24810_, _24809_, _24806_);
  and _76156_ (_24811_, _14945_, _07954_);
  or _76157_ (_24812_, _24747_, _09107_);
  or _76158_ (_24813_, _24812_, _24811_);
  and _76159_ (_24814_, _24813_, _09112_);
  and _76160_ (_24815_, _24814_, _24810_);
  and _76161_ (_24816_, _24749_, _06602_);
  or _76162_ (_24817_, _24816_, _24815_);
  and _76163_ (_24818_, _24817_, _07048_);
  and _76164_ (_24819_, _24759_, _06639_);
  or _76165_ (_24820_, _24819_, _06646_);
  or _76166_ (_24821_, _24820_, _24818_);
  and _76167_ (_24822_, _15129_, _07954_);
  or _76168_ (_24823_, _24747_, _06651_);
  or _76169_ (_24824_, _24823_, _24822_);
  and _76170_ (_24826_, _24824_, _01442_);
  and _76171_ (_24827_, _24826_, _24821_);
  or _76172_ (_24828_, _24827_, _24746_);
  and _76173_ (_44199_, _24828_, _43634_);
  and _76174_ (_24829_, _12109_, \oc8051_golden_model_1.TH0 [3]);
  or _76175_ (_24830_, _24829_, _08359_);
  and _76176_ (_24831_, _07954_, _09014_);
  or _76177_ (_24832_, _24831_, _24829_);
  and _76178_ (_24833_, _24832_, _06507_);
  and _76179_ (_24834_, _24833_, _24830_);
  nor _76180_ (_24836_, _10574_, _12109_);
  or _76181_ (_24837_, _24836_, _24829_);
  and _76182_ (_24838_, _07954_, \oc8051_golden_model_1.ACC [3]);
  nand _76183_ (_24839_, _24838_, _08359_);
  and _76184_ (_24840_, _24839_, _06615_);
  and _76185_ (_24841_, _24840_, _24837_);
  and _76186_ (_24842_, _15153_, _07954_);
  or _76187_ (_24843_, _24842_, _24829_);
  or _76188_ (_24844_, _24843_, _07275_);
  or _76189_ (_24845_, _24838_, _24829_);
  and _76190_ (_24847_, _24845_, _07259_);
  and _76191_ (_24848_, _07260_, \oc8051_golden_model_1.TH0 [3]);
  or _76192_ (_24849_, _24848_, _06474_);
  or _76193_ (_24850_, _24849_, _24847_);
  and _76194_ (_24851_, _24850_, _06772_);
  and _76195_ (_24852_, _24851_, _24844_);
  nor _76196_ (_24853_, _12109_, _07680_);
  or _76197_ (_24854_, _24853_, _24829_);
  and _76198_ (_24855_, _24854_, _06410_);
  or _76199_ (_24856_, _24855_, _24852_);
  and _76200_ (_24858_, _24856_, _06426_);
  and _76201_ (_24859_, _24845_, _06417_);
  or _76202_ (_24860_, _24859_, _10153_);
  or _76203_ (_24861_, _24860_, _24858_);
  or _76204_ (_24862_, _24854_, _06327_);
  and _76205_ (_24863_, _24862_, _24861_);
  or _76206_ (_24864_, _24863_, _09572_);
  and _76207_ (_24865_, _09310_, _07954_);
  or _76208_ (_24866_, _24829_, _06333_);
  or _76209_ (_24867_, _24866_, _24865_);
  and _76210_ (_24869_, _24867_, _06313_);
  and _76211_ (_24870_, _24869_, _24864_);
  and _76212_ (_24871_, _15251_, _07954_);
  or _76213_ (_24872_, _24871_, _24829_);
  and _76214_ (_24873_, _24872_, _06037_);
  or _76215_ (_24874_, _24873_, _06277_);
  or _76216_ (_24875_, _24874_, _24870_);
  or _76217_ (_24876_, _24832_, _06278_);
  and _76218_ (_24877_, _24876_, _24875_);
  or _76219_ (_24878_, _24877_, _06502_);
  and _76220_ (_24880_, _15266_, _07954_);
  or _76221_ (_24881_, _24829_, _07334_);
  or _76222_ (_24882_, _24881_, _24880_);
  and _76223_ (_24883_, _24882_, _07337_);
  and _76224_ (_24884_, _24883_, _24878_);
  or _76225_ (_24885_, _24884_, _24841_);
  and _76226_ (_24886_, _24885_, _07339_);
  or _76227_ (_24887_, _24886_, _24834_);
  and _76228_ (_24888_, _24887_, _07331_);
  and _76229_ (_24889_, _24845_, _06610_);
  and _76230_ (_24891_, _24889_, _24830_);
  or _76231_ (_24892_, _24891_, _06509_);
  or _76232_ (_24893_, _24892_, _24888_);
  and _76233_ (_24894_, _15263_, _07954_);
  or _76234_ (_24895_, _24829_, _09107_);
  or _76235_ (_24896_, _24895_, _24894_);
  and _76236_ (_24897_, _24896_, _09112_);
  and _76237_ (_24898_, _24897_, _24893_);
  and _76238_ (_24899_, _24837_, _06602_);
  or _76239_ (_24900_, _24899_, _06639_);
  or _76240_ (_24902_, _24900_, _24898_);
  or _76241_ (_24903_, _24843_, _07048_);
  and _76242_ (_24904_, _24903_, _06651_);
  and _76243_ (_24905_, _24904_, _24902_);
  and _76244_ (_24906_, _15321_, _07954_);
  or _76245_ (_24907_, _24906_, _24829_);
  and _76246_ (_24908_, _24907_, _06646_);
  or _76247_ (_24909_, _24908_, _01446_);
  or _76248_ (_24910_, _24909_, _24905_);
  or _76249_ (_24911_, _01442_, \oc8051_golden_model_1.TH0 [3]);
  and _76250_ (_24913_, _24911_, _43634_);
  and _76251_ (_44200_, _24913_, _24910_);
  and _76252_ (_24914_, _12109_, \oc8051_golden_model_1.TH0 [4]);
  nor _76253_ (_24915_, _10589_, _12109_);
  or _76254_ (_24916_, _24915_, _24914_);
  and _76255_ (_24917_, _07954_, \oc8051_golden_model_1.ACC [4]);
  nand _76256_ (_24918_, _24917_, _08599_);
  and _76257_ (_24919_, _24918_, _06615_);
  and _76258_ (_24920_, _24919_, _24916_);
  and _76259_ (_24921_, _15367_, _07954_);
  or _76260_ (_24922_, _24921_, _24914_);
  or _76261_ (_24923_, _24922_, _07275_);
  or _76262_ (_24924_, _24917_, _24914_);
  and _76263_ (_24925_, _24924_, _07259_);
  and _76264_ (_24926_, _07260_, \oc8051_golden_model_1.TH0 [4]);
  or _76265_ (_24927_, _24926_, _06474_);
  or _76266_ (_24928_, _24927_, _24925_);
  and _76267_ (_24929_, _24928_, _06772_);
  and _76268_ (_24930_, _24929_, _24923_);
  nor _76269_ (_24931_, _08596_, _12109_);
  or _76270_ (_24932_, _24931_, _24914_);
  and _76271_ (_24933_, _24932_, _06410_);
  or _76272_ (_24934_, _24933_, _24930_);
  and _76273_ (_24935_, _24934_, _06426_);
  and _76274_ (_24936_, _24924_, _06417_);
  or _76275_ (_24937_, _24936_, _10153_);
  or _76276_ (_24938_, _24937_, _24935_);
  or _76277_ (_24939_, _24932_, _06327_);
  and _76278_ (_24940_, _24939_, _24938_);
  or _76279_ (_24941_, _24940_, _09572_);
  and _76280_ (_24943_, _09264_, _07954_);
  or _76281_ (_24944_, _24914_, _16672_);
  or _76282_ (_24945_, _24944_, _24943_);
  and _76283_ (_24946_, _24945_, _24941_);
  or _76284_ (_24947_, _24946_, _06037_);
  and _76285_ (_24948_, _15452_, _07954_);
  or _76286_ (_24949_, _24914_, _06313_);
  or _76287_ (_24950_, _24949_, _24948_);
  and _76288_ (_24951_, _24950_, _06278_);
  and _76289_ (_24952_, _24951_, _24947_);
  and _76290_ (_24954_, _08995_, _07954_);
  or _76291_ (_24955_, _24954_, _24914_);
  and _76292_ (_24956_, _24955_, _06277_);
  or _76293_ (_24957_, _24956_, _06502_);
  or _76294_ (_24958_, _24957_, _24952_);
  and _76295_ (_24959_, _15345_, _07954_);
  or _76296_ (_24960_, _24914_, _07334_);
  or _76297_ (_24961_, _24960_, _24959_);
  and _76298_ (_24962_, _24961_, _07337_);
  and _76299_ (_24963_, _24962_, _24958_);
  or _76300_ (_24965_, _24963_, _24920_);
  and _76301_ (_24966_, _24965_, _07339_);
  or _76302_ (_24967_, _24914_, _08599_);
  and _76303_ (_24968_, _24955_, _06507_);
  and _76304_ (_24969_, _24968_, _24967_);
  or _76305_ (_24970_, _24969_, _24966_);
  and _76306_ (_24971_, _24970_, _07331_);
  and _76307_ (_24972_, _24924_, _06610_);
  and _76308_ (_24973_, _24972_, _24967_);
  or _76309_ (_24974_, _24973_, _06509_);
  or _76310_ (_24976_, _24974_, _24971_);
  and _76311_ (_24977_, _15342_, _07954_);
  or _76312_ (_24978_, _24914_, _09107_);
  or _76313_ (_24979_, _24978_, _24977_);
  and _76314_ (_24980_, _24979_, _09112_);
  and _76315_ (_24981_, _24980_, _24976_);
  and _76316_ (_24982_, _24916_, _06602_);
  or _76317_ (_24983_, _24982_, _06639_);
  or _76318_ (_24984_, _24983_, _24981_);
  or _76319_ (_24985_, _24922_, _07048_);
  and _76320_ (_24987_, _24985_, _06651_);
  and _76321_ (_24988_, _24987_, _24984_);
  and _76322_ (_24989_, _15524_, _07954_);
  or _76323_ (_24990_, _24989_, _24914_);
  and _76324_ (_24991_, _24990_, _06646_);
  or _76325_ (_24992_, _24991_, _01446_);
  or _76326_ (_24993_, _24992_, _24988_);
  or _76327_ (_24994_, _01442_, \oc8051_golden_model_1.TH0 [4]);
  and _76328_ (_24995_, _24994_, _43634_);
  and _76329_ (_44201_, _24995_, _24993_);
  and _76330_ (_24997_, _12109_, \oc8051_golden_model_1.TH0 [5]);
  nor _76331_ (_24998_, _10570_, _12109_);
  or _76332_ (_24999_, _24998_, _24997_);
  and _76333_ (_25000_, _07954_, \oc8051_golden_model_1.ACC [5]);
  nand _76334_ (_25001_, _25000_, _08308_);
  and _76335_ (_25002_, _25001_, _06615_);
  and _76336_ (_25003_, _25002_, _24999_);
  and _76337_ (_25004_, _15550_, _07954_);
  or _76338_ (_25005_, _25004_, _24997_);
  or _76339_ (_25006_, _25005_, _07275_);
  or _76340_ (_25007_, _25000_, _24997_);
  and _76341_ (_25008_, _25007_, _07259_);
  and _76342_ (_25009_, _07260_, \oc8051_golden_model_1.TH0 [5]);
  or _76343_ (_25010_, _25009_, _06474_);
  or _76344_ (_25011_, _25010_, _25008_);
  and _76345_ (_25012_, _25011_, _06772_);
  and _76346_ (_25013_, _25012_, _25006_);
  nor _76347_ (_25014_, _08305_, _12109_);
  or _76348_ (_25015_, _25014_, _24997_);
  and _76349_ (_25016_, _25015_, _06410_);
  or _76350_ (_25019_, _25016_, _25013_);
  and _76351_ (_25020_, _25019_, _06426_);
  and _76352_ (_25021_, _25007_, _06417_);
  or _76353_ (_25022_, _25021_, _10153_);
  or _76354_ (_25023_, _25022_, _25020_);
  or _76355_ (_25024_, _25015_, _06327_);
  and _76356_ (_25025_, _25024_, _25023_);
  or _76357_ (_25026_, _25025_, _09572_);
  and _76358_ (_25027_, _09218_, _07954_);
  or _76359_ (_25028_, _24997_, _06333_);
  or _76360_ (_25030_, _25028_, _25027_);
  and _76361_ (_25031_, _25030_, _06313_);
  and _76362_ (_25032_, _25031_, _25026_);
  and _76363_ (_25033_, _15649_, _07954_);
  or _76364_ (_25034_, _25033_, _24997_);
  and _76365_ (_25035_, _25034_, _06037_);
  or _76366_ (_25036_, _25035_, _06277_);
  or _76367_ (_25037_, _25036_, _25032_);
  and _76368_ (_25038_, _08954_, _07954_);
  or _76369_ (_25039_, _25038_, _24997_);
  or _76370_ (_25041_, _25039_, _06278_);
  and _76371_ (_25042_, _25041_, _25037_);
  or _76372_ (_25043_, _25042_, _06502_);
  and _76373_ (_25044_, _15664_, _07954_);
  or _76374_ (_25045_, _24997_, _07334_);
  or _76375_ (_25046_, _25045_, _25044_);
  and _76376_ (_25047_, _25046_, _07337_);
  and _76377_ (_25048_, _25047_, _25043_);
  or _76378_ (_25049_, _25048_, _25003_);
  and _76379_ (_25050_, _25049_, _07339_);
  or _76380_ (_25052_, _24997_, _08308_);
  and _76381_ (_25053_, _25039_, _06507_);
  and _76382_ (_25054_, _25053_, _25052_);
  or _76383_ (_25055_, _25054_, _25050_);
  and _76384_ (_25056_, _25055_, _07331_);
  and _76385_ (_25057_, _25007_, _06610_);
  and _76386_ (_25058_, _25057_, _25052_);
  or _76387_ (_25059_, _25058_, _06509_);
  or _76388_ (_25060_, _25059_, _25056_);
  and _76389_ (_25061_, _15663_, _07954_);
  or _76390_ (_25063_, _24997_, _09107_);
  or _76391_ (_25064_, _25063_, _25061_);
  and _76392_ (_25065_, _25064_, _09112_);
  and _76393_ (_25066_, _25065_, _25060_);
  and _76394_ (_25067_, _24999_, _06602_);
  or _76395_ (_25068_, _25067_, _06639_);
  or _76396_ (_25069_, _25068_, _25066_);
  or _76397_ (_25070_, _25005_, _07048_);
  and _76398_ (_25071_, _25070_, _06651_);
  and _76399_ (_25072_, _25071_, _25069_);
  and _76400_ (_25074_, _15721_, _07954_);
  or _76401_ (_25075_, _25074_, _24997_);
  and _76402_ (_25076_, _25075_, _06646_);
  or _76403_ (_25077_, _25076_, _01446_);
  or _76404_ (_25078_, _25077_, _25072_);
  or _76405_ (_25079_, _01442_, \oc8051_golden_model_1.TH0 [5]);
  and _76406_ (_25080_, _25079_, _43634_);
  and _76407_ (_44203_, _25080_, _25078_);
  and _76408_ (_25081_, _12109_, \oc8051_golden_model_1.TH0 [6]);
  and _76409_ (_25082_, _15759_, _07954_);
  or _76410_ (_25084_, _25082_, _25081_);
  or _76411_ (_25085_, _25084_, _07275_);
  and _76412_ (_25086_, _07954_, \oc8051_golden_model_1.ACC [6]);
  or _76413_ (_25087_, _25086_, _25081_);
  and _76414_ (_25088_, _25087_, _07259_);
  and _76415_ (_25089_, _07260_, \oc8051_golden_model_1.TH0 [6]);
  or _76416_ (_25090_, _25089_, _06474_);
  or _76417_ (_25091_, _25090_, _25088_);
  and _76418_ (_25092_, _25091_, _06772_);
  and _76419_ (_25093_, _25092_, _25085_);
  nor _76420_ (_25095_, _08209_, _12109_);
  or _76421_ (_25096_, _25095_, _25081_);
  and _76422_ (_25097_, _25096_, _06410_);
  or _76423_ (_25098_, _25097_, _25093_);
  and _76424_ (_25099_, _25098_, _06426_);
  and _76425_ (_25100_, _25087_, _06417_);
  or _76426_ (_25101_, _25100_, _10153_);
  or _76427_ (_25102_, _25101_, _25099_);
  or _76428_ (_25103_, _25096_, _06327_);
  and _76429_ (_25104_, _25103_, _25102_);
  or _76430_ (_25106_, _25104_, _09572_);
  and _76431_ (_25107_, _09172_, _07954_);
  or _76432_ (_25108_, _25081_, _06333_);
  or _76433_ (_25109_, _25108_, _25107_);
  and _76434_ (_25110_, _25109_, _06313_);
  and _76435_ (_25111_, _25110_, _25106_);
  and _76436_ (_25112_, _15846_, _07954_);
  or _76437_ (_25113_, _25112_, _25081_);
  and _76438_ (_25114_, _25113_, _06037_);
  or _76439_ (_25115_, _25114_, _06277_);
  or _76440_ (_25117_, _25115_, _25111_);
  and _76441_ (_25118_, _15853_, _07954_);
  or _76442_ (_25119_, _25118_, _25081_);
  or _76443_ (_25120_, _25119_, _06278_);
  and _76444_ (_25121_, _25120_, _25117_);
  or _76445_ (_25122_, _25121_, _06502_);
  and _76446_ (_25123_, _15862_, _07954_);
  or _76447_ (_25124_, _25081_, _07334_);
  or _76448_ (_25125_, _25124_, _25123_);
  and _76449_ (_25126_, _25125_, _07337_);
  and _76450_ (_25128_, _25126_, _25122_);
  and _76451_ (_25129_, _10596_, _07954_);
  or _76452_ (_25130_, _25129_, _25081_);
  and _76453_ (_25131_, _25130_, _06615_);
  or _76454_ (_25132_, _25131_, _25128_);
  and _76455_ (_25133_, _25132_, _07339_);
  or _76456_ (_25134_, _25081_, _08212_);
  and _76457_ (_25135_, _25119_, _06507_);
  and _76458_ (_25136_, _25135_, _25134_);
  or _76459_ (_25137_, _25136_, _25133_);
  and _76460_ (_25139_, _25137_, _07331_);
  and _76461_ (_25140_, _25087_, _06610_);
  and _76462_ (_25141_, _25140_, _25134_);
  or _76463_ (_25142_, _25141_, _06509_);
  or _76464_ (_25143_, _25142_, _25139_);
  and _76465_ (_25144_, _15859_, _07954_);
  or _76466_ (_25145_, _25081_, _09107_);
  or _76467_ (_25146_, _25145_, _25144_);
  and _76468_ (_25147_, _25146_, _09112_);
  and _76469_ (_25148_, _25147_, _25143_);
  nor _76470_ (_25150_, _10595_, _12109_);
  or _76471_ (_25151_, _25150_, _25081_);
  and _76472_ (_25152_, _25151_, _06602_);
  or _76473_ (_25153_, _25152_, _06639_);
  or _76474_ (_25154_, _25153_, _25148_);
  or _76475_ (_25155_, _25084_, _07048_);
  and _76476_ (_25156_, _25155_, _06651_);
  and _76477_ (_25157_, _25156_, _25154_);
  and _76478_ (_25158_, _15921_, _07954_);
  or _76479_ (_25159_, _25158_, _25081_);
  and _76480_ (_25161_, _25159_, _06646_);
  or _76481_ (_25162_, _25161_, _01446_);
  or _76482_ (_25163_, _25162_, _25157_);
  or _76483_ (_25164_, _01442_, \oc8051_golden_model_1.TH0 [6]);
  and _76484_ (_25165_, _25164_, _43634_);
  and _76485_ (_44204_, _25165_, _25163_);
  and _76486_ (_25166_, _13105_, _05701_);
  and _76487_ (_25167_, _13037_, \oc8051_golden_model_1.PC [0]);
  and _76488_ (_25168_, _06950_, \oc8051_golden_model_1.PC [0]);
  nor _76489_ (_25169_, _25168_, _12446_);
  nor _76490_ (_25171_, _25169_, _13037_);
  nor _76491_ (_25172_, _25171_, _25167_);
  and _76492_ (_25173_, _25172_, _05989_);
  and _76493_ (_25174_, _13072_, _09123_);
  nor _76494_ (_25175_, _25174_, _05701_);
  and _76495_ (_25176_, _12201_, _13049_);
  nor _76496_ (_25177_, _25176_, _05701_);
  nor _76497_ (_25178_, _10968_, _05701_);
  and _76498_ (_25179_, _10968_, _05701_);
  nor _76499_ (_25180_, _25179_, _25178_);
  nor _76500_ (_25182_, _25180_, _12832_);
  nor _76501_ (_25183_, _06950_, _06023_);
  and _76502_ (_25184_, _12320_, _09107_);
  nor _76503_ (_25185_, _25184_, _05701_);
  nor _76504_ (_25186_, _10975_, _05701_);
  and _76505_ (_25187_, _10975_, _05701_);
  nor _76506_ (_25188_, _25187_, _25186_);
  nor _76507_ (_25189_, _25188_, _12810_);
  and _76508_ (_25190_, _12328_, _07339_);
  nor _76509_ (_25191_, _25190_, _05701_);
  and _76510_ (_25193_, _12333_, _07334_);
  nor _76511_ (_25194_, _25193_, _05701_);
  and _76512_ (_25195_, _06277_, _05701_);
  nor _76513_ (_25196_, _06950_, _06055_);
  nor _76514_ (_25197_, _12379_, \oc8051_golden_model_1.PC [0]);
  and _76515_ (_25198_, _25169_, _12379_);
  or _76516_ (_25199_, _25198_, _06473_);
  nor _76517_ (_25200_, _25199_, _25197_);
  nor _76518_ (_25201_, _06950_, _06057_);
  and _76519_ (_25202_, _12519_, _05701_);
  nor _76520_ (_25204_, _12519_, _05701_);
  nor _76521_ (_25205_, _25204_, _25202_);
  and _76522_ (_25206_, _25205_, _07564_);
  not _76523_ (_25207_, _12516_);
  nor _76524_ (_25208_, _06950_, _07564_);
  or _76525_ (_25209_, _25208_, _25207_);
  nor _76526_ (_25210_, _25209_, _25206_);
  nor _76527_ (_25211_, _12516_, _05701_);
  nor _76528_ (_25212_, _25211_, _25210_);
  nor _76529_ (_25213_, _25212_, _08687_);
  and _76530_ (_25215_, _12539_, \oc8051_golden_model_1.PC [0]);
  and _76531_ (_25216_, _06310_, _05701_);
  nor _76532_ (_25217_, _25216_, _12260_);
  and _76533_ (_25218_, _25217_, _12537_);
  or _76534_ (_25219_, _25218_, _25215_);
  nor _76535_ (_25220_, _25219_, _08685_);
  nor _76536_ (_25221_, _25220_, _25213_);
  nor _76537_ (_25222_, _25221_, _07269_);
  and _76538_ (_25223_, _07269_, \oc8051_golden_model_1.PC [0]);
  nor _76539_ (_25224_, _25223_, _25222_);
  and _76540_ (_25226_, _25224_, _07275_);
  not _76541_ (_25227_, _25226_);
  not _76542_ (_25228_, _12502_);
  and _76543_ (_25229_, _12512_, _05701_);
  and _76544_ (_25230_, _25169_, _12510_);
  or _76545_ (_25231_, _25230_, _25229_);
  and _76546_ (_25232_, _25231_, _06474_);
  nor _76547_ (_25233_, _25232_, _25228_);
  and _76548_ (_25234_, _25233_, _25227_);
  nor _76549_ (_25235_, _12502_, _05701_);
  nor _76550_ (_25237_, _25235_, _07692_);
  not _76551_ (_25238_, _25237_);
  nor _76552_ (_25239_, _25238_, _25234_);
  nor _76553_ (_25240_, _06950_, _06052_);
  and _76554_ (_25241_, _12561_, _12551_);
  not _76555_ (_25242_, _25241_);
  nor _76556_ (_25243_, _25242_, _25240_);
  not _76557_ (_25244_, _25243_);
  nor _76558_ (_25245_, _25244_, _25239_);
  nor _76559_ (_25246_, _25241_, _05701_);
  nor _76560_ (_25248_, _25246_, _12565_);
  not _76561_ (_25249_, _25248_);
  nor _76562_ (_25250_, _25249_, _25245_);
  nor _76563_ (_25251_, _25250_, _25201_);
  or _76564_ (_25252_, _25251_, _12611_);
  and _76565_ (_25253_, _12609_, \oc8051_golden_model_1.PC [0]);
  nor _76566_ (_25254_, _25169_, _12609_);
  or _76567_ (_25255_, _25254_, _12574_);
  or _76568_ (_25256_, _25255_, _25253_);
  and _76569_ (_25257_, _25256_, _06473_);
  and _76570_ (_25259_, _25257_, _25252_);
  nor _76571_ (_25260_, _25259_, _06431_);
  not _76572_ (_25261_, _25260_);
  nor _76573_ (_25262_, _25261_, _25200_);
  and _76574_ (_25263_, _12630_, _05701_);
  not _76575_ (_25264_, _25169_);
  nor _76576_ (_25265_, _25264_, _12630_);
  nor _76577_ (_25266_, _25265_, _25263_);
  nor _76578_ (_25267_, _25266_, _06500_);
  nor _76579_ (_25268_, _25267_, _25262_);
  nor _76580_ (_25269_, _25268_, _06490_);
  and _76581_ (_25270_, _12648_, _05701_);
  nor _76582_ (_25271_, _25264_, _12648_);
  nor _76583_ (_25272_, _25271_, _25270_);
  nor _76584_ (_25273_, _25272_, _12349_);
  or _76585_ (_25274_, _25273_, _25269_);
  and _76586_ (_25275_, _25274_, _12348_);
  and _76587_ (_25276_, _12347_, _05701_);
  or _76588_ (_25277_, _25276_, _25275_);
  and _76589_ (_25278_, _25277_, _06049_);
  nor _76590_ (_25281_, _06950_, _06049_);
  nor _76591_ (_25282_, _25281_, _12345_);
  not _76592_ (_25283_, _25282_);
  nor _76593_ (_25284_, _25283_, _25278_);
  not _76594_ (_25285_, _06055_);
  nor _76595_ (_25286_, _12344_, _05701_);
  nor _76596_ (_25287_, _25286_, _25285_);
  not _76597_ (_25288_, _25287_);
  nor _76598_ (_25289_, _25288_, _25284_);
  and _76599_ (_25290_, _12339_, _06043_);
  not _76600_ (_25292_, _25290_);
  or _76601_ (_25293_, _25292_, _25289_);
  nor _76602_ (_25294_, _25293_, _25196_);
  nor _76603_ (_25295_, _25290_, _05701_);
  nor _76604_ (_25296_, _25295_, _06039_);
  not _76605_ (_25297_, _25296_);
  nor _76606_ (_25298_, _25297_, _25294_);
  nor _76607_ (_25299_, _06950_, _07745_);
  nor _76608_ (_25300_, _06486_, _06037_);
  and _76609_ (_25301_, _25300_, _12694_);
  not _76610_ (_25303_, _25301_);
  nor _76611_ (_25304_, _25303_, _25299_);
  not _76612_ (_25305_, _25304_);
  nor _76613_ (_25306_, _25305_, _25298_);
  nor _76614_ (_25307_, _25301_, _05701_);
  nor _76615_ (_25308_, _25307_, _12696_);
  not _76616_ (_25309_, _25308_);
  nor _76617_ (_25310_, _25309_, _25306_);
  nor _76618_ (_25311_, _06950_, _06004_);
  or _76619_ (_25312_, _25311_, _12704_);
  nor _76620_ (_25314_, _25312_, _25310_);
  nor _76621_ (_25315_, _25217_, _12705_);
  nor _76622_ (_25316_, _25315_, _25314_);
  and _76623_ (_25317_, _25316_, _06278_);
  or _76624_ (_25318_, _25317_, _25195_);
  and _76625_ (_25319_, _25318_, _12719_);
  and _76626_ (_25320_, _12718_, _06046_);
  or _76627_ (_25321_, _25320_, _25319_);
  and _76628_ (_25322_, _25321_, _06009_);
  nor _76629_ (_25323_, _06950_, _06009_);
  or _76630_ (_25325_, _25323_, _25322_);
  and _76631_ (_25326_, _25325_, _12764_);
  not _76632_ (_25327_, _25193_);
  nor _76633_ (_25328_, _25217_, _11389_);
  and _76634_ (_25329_, _11389_, _05701_);
  nor _76635_ (_25330_, _25329_, _12764_);
  not _76636_ (_25331_, _25330_);
  nor _76637_ (_25332_, _25331_, _25328_);
  nor _76638_ (_25333_, _25332_, _25327_);
  not _76639_ (_25334_, _25333_);
  nor _76640_ (_25336_, _25334_, _25326_);
  nor _76641_ (_25337_, _25336_, _25194_);
  and _76642_ (_25338_, _25337_, _06012_);
  nor _76643_ (_25339_, _06950_, _06012_);
  or _76644_ (_25340_, _25339_, _25338_);
  and _76645_ (_25341_, _25340_, _12788_);
  not _76646_ (_25342_, _25190_);
  nor _76647_ (_25343_, _11389_, _05701_);
  and _76648_ (_25344_, _25217_, _11389_);
  or _76649_ (_25345_, _25344_, _25343_);
  and _76650_ (_25347_, _25345_, _12787_);
  nor _76651_ (_25348_, _25347_, _25342_);
  not _76652_ (_25349_, _25348_);
  nor _76653_ (_25350_, _25349_, _25341_);
  nor _76654_ (_25351_, _25350_, _25191_);
  and _76655_ (_25352_, _25351_, _06018_);
  nor _76656_ (_25353_, _06950_, _06018_);
  or _76657_ (_25354_, _25353_, _25352_);
  and _76658_ (_25355_, _25354_, _12810_);
  not _76659_ (_25356_, _25184_);
  or _76660_ (_25358_, _25356_, _25355_);
  nor _76661_ (_25359_, _25358_, _25189_);
  or _76662_ (_25360_, _25359_, _12827_);
  nor _76663_ (_25361_, _25360_, _25185_);
  nor _76664_ (_25362_, _25361_, _25183_);
  nor _76665_ (_25363_, _25362_, _12310_);
  and _76666_ (_25364_, _12837_, _11217_);
  not _76667_ (_25365_, _25364_);
  or _76668_ (_25366_, _25365_, _25363_);
  nor _76669_ (_25367_, _25366_, _25182_);
  nor _76670_ (_25369_, _25364_, _05701_);
  nor _76671_ (_25370_, _25369_, _06621_);
  not _76672_ (_25371_, _25370_);
  nor _76673_ (_25372_, _25371_, _25367_);
  and _76674_ (_25373_, _09447_, _06621_);
  or _76675_ (_25374_, _25373_, _25372_);
  and _76676_ (_25375_, _25374_, _06016_);
  nor _76677_ (_25376_, _06950_, _06016_);
  or _76678_ (_25377_, _25376_, _25375_);
  and _76679_ (_25378_, _25377_, _06629_);
  and _76680_ (_25380_, _25264_, _13037_);
  nor _76681_ (_25381_, _13037_, _05701_);
  or _76682_ (_25382_, _25381_, _06629_);
  or _76683_ (_25383_, _25382_, _25380_);
  and _76684_ (_25384_, _25383_, _25176_);
  not _76685_ (_25385_, _25384_);
  nor _76686_ (_25386_, _25385_, _25378_);
  nor _76687_ (_25387_, _25386_, _25177_);
  and _76688_ (_25388_, _25387_, _06362_);
  and _76689_ (_25389_, _09447_, _06361_);
  or _76690_ (_25391_, _25389_, _25388_);
  and _76691_ (_25392_, _25391_, _06021_);
  nor _76692_ (_25393_, _06950_, _06021_);
  nor _76693_ (_25394_, _25393_, _25392_);
  nor _76694_ (_25395_, _25394_, _06496_);
  not _76695_ (_25396_, _25174_);
  and _76696_ (_25397_, _25172_, _06496_);
  nor _76697_ (_25398_, _25397_, _25396_);
  not _76698_ (_25399_, _25398_);
  nor _76699_ (_25400_, _25399_, _25395_);
  nor _76700_ (_25402_, _25400_, _25175_);
  nor _76701_ (_25403_, _25402_, _07783_);
  and _76702_ (_25404_, _07783_, _06950_);
  nor _76703_ (_25405_, _25404_, _05989_);
  not _76704_ (_25406_, _25405_);
  nor _76705_ (_25407_, _25406_, _25403_);
  nor _76706_ (_25408_, _25407_, _25173_);
  and _76707_ (_25409_, _13095_, _13087_);
  not _76708_ (_25410_, _25409_);
  nor _76709_ (_25411_, _25410_, _25408_);
  nor _76710_ (_25413_, _06488_, _05997_);
  not _76711_ (_25414_, _25413_);
  nor _76712_ (_25415_, _25409_, \oc8051_golden_model_1.PC [0]);
  nor _76713_ (_25416_, _25415_, _25414_);
  not _76714_ (_25417_, _25416_);
  nor _76715_ (_25418_, _25417_, _25411_);
  and _76716_ (_25419_, _25414_, _06950_);
  nor _76717_ (_25420_, _25419_, _13105_);
  not _76718_ (_25421_, _25420_);
  nor _76719_ (_25422_, _25421_, _25418_);
  nor _76720_ (_25424_, _25422_, _25166_);
  nand _76721_ (_25425_, _25424_, _01442_);
  or _76722_ (_25426_, _01442_, \oc8051_golden_model_1.PC [0]);
  and _76723_ (_25427_, _25426_, _43634_);
  and _76724_ (_44206_, _25427_, _25425_);
  and _76725_ (_25428_, _13105_, _12444_);
  and _76726_ (_25429_, _06646_, _05667_);
  and _76727_ (_25430_, _13037_, _12444_);
  nor _76728_ (_25431_, _12448_, _12446_);
  nor _76729_ (_25432_, _25431_, _12449_);
  nor _76730_ (_25434_, _25432_, _13037_);
  nor _76731_ (_25435_, _25434_, _25430_);
  and _76732_ (_25436_, _25435_, _05989_);
  and _76733_ (_25437_, _06639_, _05667_);
  nor _76734_ (_25438_, _12201_, _12444_);
  nor _76735_ (_25439_, _12837_, _12444_);
  and _76736_ (_25440_, _12318_, _06089_);
  and _76737_ (_25441_, _12326_, _06089_);
  nor _76738_ (_25442_, _17563_, _12444_);
  or _76739_ (_25443_, _12339_, _12444_);
  nand _76740_ (_25445_, _12347_, _06089_);
  and _76741_ (_25446_, _07269_, _12444_);
  nor _76742_ (_25447_, _07160_, _07564_);
  nor _76743_ (_25448_, _12518_, _05701_);
  nor _76744_ (_25449_, _25448_, _07259_);
  nor _76745_ (_25450_, _25449_, \oc8051_golden_model_1.PC [1]);
  and _76746_ (_25451_, _25449_, \oc8051_golden_model_1.PC [1]);
  or _76747_ (_25452_, _25451_, _25450_);
  or _76748_ (_25453_, _25452_, _06855_);
  nand _76749_ (_25454_, _06855_, _06089_);
  and _76750_ (_25456_, _25454_, _07564_);
  and _76751_ (_25457_, _25456_, _25453_);
  or _76752_ (_25458_, _25457_, _25207_);
  or _76753_ (_25459_, _25458_, _25447_);
  or _76754_ (_25460_, _12516_, _12444_);
  and _76755_ (_25461_, _25460_, _08685_);
  and _76756_ (_25462_, _25461_, _25459_);
  or _76757_ (_25463_, _12537_, _05667_);
  nor _76758_ (_25464_, _12262_, _12260_);
  nor _76759_ (_25465_, _25464_, _12263_);
  or _76760_ (_25467_, _25465_, _12539_);
  and _76761_ (_25468_, _25467_, _08687_);
  and _76762_ (_25469_, _25468_, _25463_);
  or _76763_ (_25470_, _25469_, _25462_);
  and _76764_ (_25471_, _25470_, _07270_);
  or _76765_ (_25472_, _25471_, _25446_);
  and _76766_ (_25473_, _25472_, _07275_);
  and _76767_ (_25474_, _25432_, _12510_);
  and _76768_ (_25475_, _12512_, _06089_);
  or _76769_ (_25476_, _25475_, _25474_);
  and _76770_ (_25478_, _25476_, _06474_);
  or _76771_ (_25479_, _25478_, _25228_);
  or _76772_ (_25480_, _25479_, _25473_);
  or _76773_ (_25481_, _12502_, _12444_);
  and _76774_ (_25482_, _25481_, _06357_);
  and _76775_ (_25483_, _25482_, _25480_);
  and _76776_ (_25484_, _06356_, _05667_);
  or _76777_ (_25485_, _25484_, _07692_);
  or _76778_ (_25486_, _25485_, _25483_);
  nand _76779_ (_25487_, _07160_, _07692_);
  and _76780_ (_25489_, _25487_, _06772_);
  and _76781_ (_25490_, _25489_, _25486_);
  nand _76782_ (_25491_, _06410_, _05667_);
  nand _76783_ (_25492_, _25491_, _12551_);
  or _76784_ (_25493_, _25492_, _25490_);
  or _76785_ (_25494_, _12551_, _12444_);
  and _76786_ (_25495_, _25494_, _06426_);
  and _76787_ (_25496_, _25495_, _25493_);
  nand _76788_ (_25497_, _06417_, _05667_);
  nand _76789_ (_25498_, _25497_, _12561_);
  or _76790_ (_25500_, _25498_, _25496_);
  or _76791_ (_25501_, _12561_, _12444_);
  and _76792_ (_25502_, _25501_, _06353_);
  and _76793_ (_25503_, _25502_, _25500_);
  and _76794_ (_25504_, _06352_, _05667_);
  or _76795_ (_25505_, _25504_, _12565_);
  or _76796_ (_25506_, _25505_, _25503_);
  nand _76797_ (_25507_, _07160_, _12565_);
  and _76798_ (_25508_, _25507_, _07394_);
  and _76799_ (_25509_, _25508_, _25506_);
  nand _76800_ (_25511_, _06351_, _05667_);
  nand _76801_ (_25512_, _25511_, _12573_);
  or _76802_ (_25513_, _25512_, _25509_);
  or _76803_ (_25514_, _25432_, _12609_);
  nand _76804_ (_25515_, _12609_, _12444_);
  and _76805_ (_25516_, _25515_, _25514_);
  and _76806_ (_25517_, _25516_, _12571_);
  or _76807_ (_25518_, _25517_, _12574_);
  and _76808_ (_25519_, _25518_, _25513_);
  and _76809_ (_25520_, _25516_, _06469_);
  or _76810_ (_25522_, _25520_, _06472_);
  or _76811_ (_25523_, _25522_, _25519_);
  nor _76812_ (_25524_, _12379_, _12444_);
  and _76813_ (_25525_, _25432_, _12379_);
  or _76814_ (_25526_, _25525_, _06473_);
  or _76815_ (_25527_, _25526_, _25524_);
  and _76816_ (_25528_, _25527_, _06500_);
  and _76817_ (_25529_, _25528_, _25523_);
  not _76818_ (_25530_, _25432_);
  nor _76819_ (_25531_, _25530_, _12630_);
  and _76820_ (_25533_, _12630_, _06089_);
  or _76821_ (_25534_, _25533_, _25531_);
  and _76822_ (_25535_, _25534_, _06431_);
  or _76823_ (_25536_, _25535_, _25529_);
  and _76824_ (_25537_, _25536_, _12349_);
  nand _76825_ (_25538_, _12648_, _12444_);
  or _76826_ (_25539_, _25432_, _12648_);
  and _76827_ (_25540_, _25539_, _06490_);
  and _76828_ (_25541_, _25540_, _25538_);
  or _76829_ (_25542_, _25541_, _12347_);
  or _76830_ (_25544_, _25542_, _25537_);
  and _76831_ (_25545_, _25544_, _25445_);
  or _76832_ (_25546_, _25545_, _06345_);
  nand _76833_ (_25547_, _06345_, \oc8051_golden_model_1.PC [1]);
  and _76834_ (_25548_, _25547_, _06049_);
  and _76835_ (_25549_, _25548_, _25546_);
  nor _76836_ (_25550_, _07160_, _06049_);
  and _76837_ (_25551_, _18528_, _07252_);
  nor _76838_ (_25552_, _25551_, _06054_);
  not _76839_ (_25553_, _25552_);
  and _76840_ (_25555_, _25553_, _12659_);
  not _76841_ (_25556_, _25555_);
  or _76842_ (_25557_, _25556_, _25550_);
  or _76843_ (_25558_, _25557_, _25549_);
  or _76844_ (_25559_, _25555_, _05667_);
  and _76845_ (_25560_, _25559_, _12342_);
  and _76846_ (_25561_, _25560_, _25558_);
  nand _76847_ (_25562_, _12341_, _12444_);
  nand _76848_ (_25563_, _25562_, _12343_);
  or _76849_ (_25564_, _25563_, _25561_);
  or _76850_ (_25566_, _12343_, _12444_);
  and _76851_ (_25567_, _25566_, _14252_);
  and _76852_ (_25568_, _25567_, _25564_);
  and _76853_ (_25569_, _06445_, _05667_);
  or _76854_ (_25570_, _25569_, _25285_);
  or _76855_ (_25571_, _25570_, _25568_);
  nand _76856_ (_25572_, _07160_, _25285_);
  and _76857_ (_25573_, _25572_, _14251_);
  and _76858_ (_25574_, _25573_, _25571_);
  nand _76859_ (_25575_, _06444_, _05667_);
  nand _76860_ (_25576_, _25575_, _12339_);
  or _76861_ (_25577_, _25576_, _25574_);
  and _76862_ (_25578_, _25577_, _25443_);
  or _76863_ (_25579_, _25578_, _12337_);
  or _76864_ (_25580_, _12336_, _05667_);
  and _76865_ (_25581_, _25580_, _06043_);
  and _76866_ (_25582_, _25581_, _25579_);
  and _76867_ (_25583_, _12444_, _06042_);
  or _76868_ (_25584_, _25583_, _06339_);
  or _76869_ (_25585_, _25584_, _25582_);
  nand _76870_ (_25588_, _06339_, \oc8051_golden_model_1.PC [1]);
  and _76871_ (_25589_, _25588_, _25585_);
  or _76872_ (_25590_, _25589_, _06039_);
  nand _76873_ (_25591_, _07160_, _06039_);
  and _76874_ (_25592_, _25591_, _06487_);
  and _76875_ (_25593_, _25592_, _25590_);
  nand _76876_ (_25594_, _06486_, _06089_);
  nand _76877_ (_25595_, _25594_, _06334_);
  or _76878_ (_25596_, _25595_, _25593_);
  or _76879_ (_25597_, _06334_, _05667_);
  and _76880_ (_25599_, _25597_, _06313_);
  and _76881_ (_25600_, _25599_, _25596_);
  nand _76882_ (_25601_, _06089_, _06037_);
  nand _76883_ (_25602_, _25601_, _12694_);
  or _76884_ (_25603_, _25602_, _25600_);
  not _76885_ (_25604_, _06401_);
  or _76886_ (_25605_, _12694_, _12444_);
  and _76887_ (_25606_, _25605_, _25604_);
  and _76888_ (_25607_, _25606_, _25603_);
  and _76889_ (_25608_, _06401_, _05667_);
  or _76890_ (_25610_, _25608_, _12696_);
  or _76891_ (_25611_, _25610_, _25607_);
  nand _76892_ (_25612_, _07160_, _12696_);
  and _76893_ (_25613_, _25612_, _12705_);
  and _76894_ (_25614_, _25613_, _25611_);
  and _76895_ (_25615_, _25465_, _12704_);
  or _76896_ (_25616_, _25615_, _08848_);
  or _76897_ (_25617_, _25616_, _25614_);
  nor _76898_ (_25618_, _06277_, \oc8051_golden_model_1.PC [1]);
  or _76899_ (_25619_, _25618_, _08627_);
  and _76900_ (_25621_, _25619_, _25617_);
  and _76901_ (_25622_, _06277_, _06089_);
  or _76902_ (_25623_, _25622_, _11028_);
  or _76903_ (_25624_, _25623_, _25621_);
  nand _76904_ (_25625_, _11028_, \oc8051_golden_model_1.PC [1]);
  nand _76905_ (_25626_, _25625_, _25624_);
  nand _76906_ (_25627_, _25626_, _12719_);
  nor _76907_ (_25628_, _12719_, _06087_);
  nor _76908_ (_25629_, _25628_, _06400_);
  nand _76909_ (_25630_, _25629_, _25627_);
  and _76910_ (_25632_, _06400_, _05667_);
  nor _76911_ (_25633_, _25632_, _06275_);
  nand _76912_ (_25634_, _25633_, _25630_);
  and _76913_ (_25635_, _07160_, _06275_);
  nor _76914_ (_25636_, _25635_, _12763_);
  nand _76915_ (_25637_, _25636_, _25634_);
  nor _76916_ (_25638_, _25465_, _11389_);
  and _76917_ (_25639_, _11389_, \oc8051_golden_model_1.PC [1]);
  nor _76918_ (_25640_, _25639_, _12764_);
  not _76919_ (_25641_, _25640_);
  nor _76920_ (_25643_, _25641_, _25638_);
  nor _76921_ (_25644_, _25643_, _17564_);
  and _76922_ (_25645_, _25644_, _25637_);
  or _76923_ (_25646_, _25645_, _25442_);
  nor _76924_ (_25647_, _17572_, _11042_);
  nand _76925_ (_25648_, _25647_, _25646_);
  nor _76926_ (_25649_, _25647_, _12444_);
  nor _76927_ (_25650_, _25649_, _17457_);
  nand _76928_ (_25651_, _25650_, _25648_);
  and _76929_ (_25652_, _17457_, _12444_);
  nor _76930_ (_25654_, _25652_, _12331_);
  nand _76931_ (_25655_, _25654_, _25651_);
  nor _76932_ (_25656_, _12330_, _05667_);
  nor _76933_ (_25657_, _25656_, _06502_);
  nand _76934_ (_25658_, _25657_, _25655_);
  and _76935_ (_25659_, _06502_, _06089_);
  nor _76936_ (_25660_, _25659_, _06615_);
  and _76937_ (_25661_, _25660_, _25658_);
  and _76938_ (_25662_, _06615_, \oc8051_golden_model_1.PC [1]);
  or _76939_ (_25663_, _25662_, _25661_);
  nand _76940_ (_25665_, _25663_, _06012_);
  and _76941_ (_25666_, _07160_, _12782_);
  nor _76942_ (_25667_, _25666_, _12787_);
  nand _76943_ (_25668_, _25667_, _25665_);
  nor _76944_ (_25669_, _25465_, _12770_);
  nor _76945_ (_25670_, _11389_, _05667_);
  nor _76946_ (_25671_, _25670_, _12788_);
  not _76947_ (_25672_, _25671_);
  nor _76948_ (_25673_, _25672_, _25669_);
  nor _76949_ (_25674_, _25673_, _12326_);
  and _76950_ (_25676_, _25674_, _25668_);
  nor _76951_ (_25677_, _25676_, _25441_);
  and _76952_ (_25678_, _06331_, _06506_);
  or _76953_ (_25679_, _12324_, _25678_);
  or _76954_ (_25680_, _25679_, _25677_);
  and _76955_ (_25681_, _25679_, _06089_);
  nor _76956_ (_25682_, _25681_, _06977_);
  nand _76957_ (_25683_, _25682_, _25680_);
  and _76958_ (_25684_, _06977_, _12444_);
  nor _76959_ (_25685_, _25684_, _12323_);
  nand _76960_ (_25687_, _25685_, _25683_);
  nor _76961_ (_25688_, _12322_, _05667_);
  nor _76962_ (_25689_, _25688_, _06507_);
  nand _76963_ (_25690_, _25689_, _25687_);
  and _76964_ (_25691_, _06507_, _06089_);
  nor _76965_ (_25692_, _25691_, _06610_);
  and _76966_ (_25693_, _25692_, _25690_);
  and _76967_ (_25694_, _06610_, \oc8051_golden_model_1.PC [1]);
  or _76968_ (_25695_, _25694_, _25693_);
  nand _76969_ (_25696_, _25695_, _06018_);
  and _76970_ (_25698_, _07160_, _07330_);
  nor _76971_ (_25699_, _25698_, _12809_);
  nand _76972_ (_25700_, _25699_, _25696_);
  nor _76973_ (_25701_, _25465_, \oc8051_golden_model_1.PSW [7]);
  and _76974_ (_25702_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor _76975_ (_25703_, _25702_, _12810_);
  not _76976_ (_25704_, _25703_);
  nor _76977_ (_25705_, _25704_, _25701_);
  nor _76978_ (_25706_, _25705_, _12318_);
  and _76979_ (_25707_, _25706_, _25700_);
  nor _76980_ (_25709_, _25707_, _25440_);
  and _76981_ (_25710_, _06331_, _06508_);
  or _76982_ (_25711_, _12316_, _25710_);
  or _76983_ (_25712_, _25711_, _25709_);
  and _76984_ (_25713_, _25711_, _06089_);
  nor _76985_ (_25714_, _25713_, _06988_);
  nand _76986_ (_25715_, _25714_, _25712_);
  and _76987_ (_25716_, _06988_, _12444_);
  nor _76988_ (_25717_, _25716_, _12315_);
  nand _76989_ (_25718_, _25717_, _25715_);
  nor _76990_ (_25720_, _12314_, _05667_);
  nor _76991_ (_25721_, _25720_, _06509_);
  nand _76992_ (_25722_, _25721_, _25718_);
  and _76993_ (_25723_, _06509_, _06089_);
  nor _76994_ (_25724_, _25723_, _06602_);
  and _76995_ (_25725_, _25724_, _25722_);
  and _76996_ (_25726_, _06602_, \oc8051_golden_model_1.PC [1]);
  or _76997_ (_25727_, _25726_, _25725_);
  nand _76998_ (_25728_, _25727_, _06023_);
  and _76999_ (_25729_, _07160_, _12827_);
  nor _77000_ (_25731_, _25729_, _12310_);
  nand _77001_ (_25732_, _25731_, _25728_);
  nor _77002_ (_25733_, _25465_, _10967_);
  and _77003_ (_25734_, _10967_, \oc8051_golden_model_1.PC [1]);
  nor _77004_ (_25735_, _25734_, _12832_);
  not _77005_ (_25736_, _25735_);
  nor _77006_ (_25737_, _25736_, _25733_);
  nor _77007_ (_25738_, _25737_, _12839_);
  and _77008_ (_25739_, _25738_, _25732_);
  or _77009_ (_25740_, _25739_, _25439_);
  nand _77010_ (_25742_, _25740_, _11187_);
  nor _77011_ (_25743_, _11187_, _05667_);
  nor _77012_ (_25744_, _25743_, _11216_);
  nand _77013_ (_25745_, _25744_, _25742_);
  and _77014_ (_25746_, _11216_, _12444_);
  nor _77015_ (_25747_, _25746_, _06621_);
  and _77016_ (_25748_, _25747_, _25745_);
  and _77017_ (_25749_, _11310_, _06621_);
  or _77018_ (_25750_, _25749_, _25748_);
  nand _77019_ (_25751_, _25750_, _06016_);
  and _77020_ (_25753_, _07160_, _07350_);
  nor _77021_ (_25754_, _25753_, _06512_);
  nand _77022_ (_25755_, _25754_, _25751_);
  nor _77023_ (_25756_, _13037_, _06089_);
  not _77024_ (_25757_, _25756_);
  and _77025_ (_25758_, _25530_, _13037_);
  nor _77026_ (_25759_, _25758_, _06629_);
  and _77027_ (_25760_, _25759_, _25757_);
  nor _77028_ (_25761_, _25760_, _12854_);
  and _77029_ (_25762_, _25761_, _25755_);
  or _77030_ (_25764_, _25762_, _25438_);
  nand _77031_ (_25765_, _25764_, _13046_);
  nor _77032_ (_25766_, _13046_, _05667_);
  nor _77033_ (_25767_, _25766_, _10564_);
  nand _77034_ (_25768_, _25767_, _25765_);
  and _77035_ (_25769_, _10564_, _12444_);
  nor _77036_ (_25770_, _25769_, _06361_);
  and _77037_ (_25771_, _25770_, _25768_);
  and _77038_ (_25772_, _11310_, _06361_);
  or _77039_ (_25773_, _25772_, _25771_);
  nand _77040_ (_25775_, _25773_, _06021_);
  and _77041_ (_25776_, _07160_, _12187_);
  nor _77042_ (_25777_, _25776_, _06496_);
  nand _77043_ (_25778_, _25777_, _25775_);
  and _77044_ (_25779_, _25435_, _06496_);
  nor _77045_ (_25780_, _25779_, _15091_);
  and _77046_ (_25781_, _25780_, _25778_);
  nor _77047_ (_25782_, _09122_, _12444_);
  or _77048_ (_25783_, _25782_, _25781_);
  nand _77049_ (_25784_, _25783_, _09121_);
  and _77050_ (_25786_, _07561_, _06089_);
  nor _77051_ (_25787_, _25786_, _06639_);
  and _77052_ (_25788_, _25787_, _25784_);
  or _77053_ (_25789_, _25788_, _25437_);
  nand _77054_ (_25790_, _25789_, _13072_);
  nor _77055_ (_25791_, _13072_, _06089_);
  nor _77056_ (_25792_, _25791_, _07783_);
  nand _77057_ (_25793_, _25792_, _25790_);
  and _77058_ (_25794_, _07783_, _07160_);
  nor _77059_ (_25795_, _25794_, _05989_);
  and _77060_ (_25797_, _25795_, _25793_);
  or _77061_ (_25798_, _25797_, _25436_);
  nand _77062_ (_25799_, _25798_, _09473_);
  nor _77063_ (_25800_, _09473_, _06089_);
  nor _77064_ (_25801_, _25800_, _07055_);
  nand _77065_ (_25802_, _25801_, _25799_);
  and _77066_ (_25803_, _07055_, _06089_);
  nor _77067_ (_25804_, _25803_, _06646_);
  and _77068_ (_25805_, _25804_, _25802_);
  or _77069_ (_25806_, _25805_, _25429_);
  nand _77070_ (_25808_, _25806_, _13095_);
  nor _77071_ (_25809_, _13095_, _06089_);
  nor _77072_ (_25810_, _25809_, _25414_);
  nand _77073_ (_25811_, _25810_, _25808_);
  and _77074_ (_25812_, _25414_, _07160_);
  nor _77075_ (_25813_, _25812_, _13105_);
  and _77076_ (_25814_, _25813_, _25811_);
  or _77077_ (_25815_, _25814_, _25428_);
  or _77078_ (_25816_, _25815_, _01446_);
  or _77079_ (_25817_, _01442_, \oc8051_golden_model_1.PC [1]);
  and _77080_ (_25819_, _25817_, _43634_);
  and _77081_ (_44207_, _25819_, _25816_);
  and _77082_ (_25820_, _06646_, _06111_);
  and _77083_ (_25821_, _06639_, _06111_);
  nor _77084_ (_25822_, _12201_, _06127_);
  nor _77085_ (_25823_, _12837_, _06127_);
  nor _77086_ (_25824_, _12320_, _06127_);
  nor _77087_ (_25825_, _12328_, _06127_);
  nor _77088_ (_25826_, _12333_, _06127_);
  nor _77089_ (_25827_, _12694_, _06127_);
  nor _77090_ (_25829_, _06326_, _06111_);
  nor _77091_ (_25830_, _25555_, _06111_);
  and _77092_ (_25831_, _12347_, _06128_);
  and _77093_ (_25832_, _12453_, _12450_);
  nor _77094_ (_25833_, _25832_, _12454_);
  not _77095_ (_25834_, _25833_);
  nand _77096_ (_25835_, _25834_, _12379_);
  or _77097_ (_25836_, _12441_, _12379_);
  nand _77098_ (_25837_, _25836_, _25835_);
  nand _77099_ (_25838_, _25837_, _06472_);
  or _77100_ (_25840_, _25833_, _12512_);
  or _77101_ (_25841_, _12510_, _12441_);
  and _77102_ (_25842_, _25841_, _25840_);
  or _77103_ (_25843_, _25842_, _07275_);
  and _77104_ (_25844_, _12539_, _06111_);
  and _77105_ (_25845_, _12267_, _12264_);
  nor _77106_ (_25846_, _25845_, _12268_);
  and _77107_ (_25847_, _25846_, _12537_);
  nor _77108_ (_25848_, _25847_, _25844_);
  nand _77109_ (_25849_, _25848_, _08687_);
  and _77110_ (_25851_, _12518_, _05673_);
  nor _77111_ (_25852_, _25851_, _07259_);
  and _77112_ (_25853_, _07259_, _06111_);
  nor _77113_ (_25854_, _25853_, _06855_);
  not _77114_ (_25855_, _25854_);
  nor _77115_ (_25856_, _25855_, _25852_);
  not _77116_ (_25857_, _25856_);
  nor _77117_ (_25858_, _12519_, _06127_);
  nor _77118_ (_25859_, _25858_, _06816_);
  and _77119_ (_25860_, _25859_, _25857_);
  nor _77120_ (_25862_, _07564_, _06769_);
  or _77121_ (_25863_, _25862_, _25207_);
  nor _77122_ (_25864_, _25863_, _25860_);
  nor _77123_ (_25865_, _12516_, _06127_);
  nor _77124_ (_25866_, _25865_, _25864_);
  nor _77125_ (_25867_, _25866_, _08687_);
  nor _77126_ (_25868_, _25867_, _07269_);
  and _77127_ (_25869_, _25868_, _25849_);
  and _77128_ (_25870_, _07269_, _06127_);
  or _77129_ (_25871_, _25870_, _06474_);
  or _77130_ (_25873_, _25871_, _25869_);
  nand _77131_ (_25874_, _25873_, _25843_);
  nand _77132_ (_25875_, _25874_, _12502_);
  nor _77133_ (_25876_, _12502_, _06127_);
  nor _77134_ (_25877_, _25876_, _06356_);
  nand _77135_ (_25878_, _25877_, _25875_);
  and _77136_ (_25879_, _06356_, _06111_);
  nor _77137_ (_25880_, _25879_, _07692_);
  nand _77138_ (_25881_, _25880_, _25878_);
  and _77139_ (_25882_, _06769_, _07692_);
  nor _77140_ (_25884_, _25882_, _06410_);
  nand _77141_ (_25885_, _25884_, _25881_);
  and _77142_ (_25886_, _06410_, _06111_);
  nor _77143_ (_25887_, _25886_, _12552_);
  nand _77144_ (_25888_, _25887_, _25885_);
  nor _77145_ (_25889_, _12551_, _06127_);
  nor _77146_ (_25890_, _25889_, _06417_);
  nand _77147_ (_25891_, _25890_, _25888_);
  and _77148_ (_25892_, _06417_, _06111_);
  nor _77149_ (_25893_, _25892_, _12563_);
  nand _77150_ (_25895_, _25893_, _25891_);
  nor _77151_ (_25896_, _12561_, _06127_);
  nor _77152_ (_25897_, _25896_, _06352_);
  nand _77153_ (_25898_, _25897_, _25895_);
  and _77154_ (_25899_, _06352_, _06111_);
  nor _77155_ (_25900_, _25899_, _12565_);
  nand _77156_ (_25901_, _25900_, _25898_);
  and _77157_ (_25902_, _06769_, _12565_);
  nor _77158_ (_25903_, _25902_, _06351_);
  nand _77159_ (_25904_, _25903_, _25901_);
  and _77160_ (_25905_, _06351_, _06111_);
  nor _77161_ (_25906_, _25905_, _12611_);
  and _77162_ (_25907_, _25906_, _25904_);
  nor _77163_ (_25908_, _25834_, _12609_);
  and _77164_ (_25909_, _12609_, _12441_);
  or _77165_ (_25910_, _25909_, _12574_);
  nor _77166_ (_25911_, _25910_, _25908_);
  or _77167_ (_25912_, _25911_, _25907_);
  nand _77168_ (_25913_, _25912_, _06473_);
  and _77169_ (_25914_, _25913_, _25838_);
  or _77170_ (_25917_, _25914_, _06431_);
  and _77171_ (_25918_, _12630_, _12441_);
  nor _77172_ (_25919_, _25834_, _12630_);
  or _77173_ (_25920_, _25919_, _06500_);
  or _77174_ (_25921_, _25920_, _25918_);
  and _77175_ (_25922_, _25921_, _12349_);
  nand _77176_ (_25923_, _25922_, _25917_);
  and _77177_ (_25924_, _12648_, _12442_);
  nor _77178_ (_25925_, _25833_, _12648_);
  or _77179_ (_25926_, _25925_, _12349_);
  nor _77180_ (_25928_, _25926_, _25924_);
  nor _77181_ (_25929_, _25928_, _12347_);
  and _77182_ (_25930_, _25929_, _25923_);
  or _77183_ (_25931_, _25930_, _25831_);
  nand _77184_ (_25932_, _25931_, _06346_);
  and _77185_ (_25933_, _06345_, _06113_);
  nor _77186_ (_25934_, _25933_, _07596_);
  nand _77187_ (_25935_, _25934_, _25932_);
  nor _77188_ (_25936_, _06769_, _06049_);
  nor _77189_ (_25937_, _25936_, _25556_);
  and _77190_ (_25939_, _25937_, _25935_);
  or _77191_ (_25940_, _25939_, _25830_);
  nand _77192_ (_25941_, _25940_, _12344_);
  nor _77193_ (_25942_, _12344_, _06127_);
  nor _77194_ (_25943_, _25942_, _06445_);
  nand _77195_ (_25944_, _25943_, _25941_);
  and _77196_ (_25945_, _06445_, _06111_);
  nor _77197_ (_25946_, _25945_, _25285_);
  nand _77198_ (_25947_, _25946_, _25944_);
  and _77199_ (_25948_, _06769_, _25285_);
  nor _77200_ (_25950_, _25948_, _06444_);
  nand _77201_ (_25951_, _25950_, _25947_);
  and _77202_ (_25952_, _06444_, _06111_);
  nor _77203_ (_25953_, _25952_, _12671_);
  and _77204_ (_25954_, _25953_, _25951_);
  nor _77205_ (_25955_, _12339_, _06127_);
  or _77206_ (_25956_, _25955_, _25954_);
  nand _77207_ (_25957_, _25956_, _12336_);
  nor _77208_ (_25958_, _12336_, _06111_);
  nor _77209_ (_25959_, _25958_, _06042_);
  nand _77210_ (_25961_, _25959_, _25957_);
  and _77211_ (_25962_, _06127_, _06042_);
  nor _77212_ (_25963_, _25962_, _06339_);
  and _77213_ (_25964_, _25963_, _25961_);
  and _77214_ (_25965_, _06339_, _06113_);
  or _77215_ (_25966_, _25965_, _25964_);
  nand _77216_ (_25967_, _25966_, _07745_);
  and _77217_ (_25968_, _06769_, _06039_);
  nor _77218_ (_25969_, _25968_, _06486_);
  nand _77219_ (_25970_, _25969_, _25967_);
  and _77220_ (_25972_, _12441_, _06486_);
  not _77221_ (_25973_, _25972_);
  and _77222_ (_25974_, _25973_, _06326_);
  and _77223_ (_25975_, _25974_, _25970_);
  nor _77224_ (_25976_, _25975_, _25829_);
  nor _77225_ (_25977_, _07252_, _06003_);
  or _77226_ (_25978_, _25977_, _25976_);
  and _77227_ (_25979_, _25977_, _06113_);
  nor _77228_ (_25980_, _25979_, _06037_);
  nand _77229_ (_25981_, _25980_, _25978_);
  and _77230_ (_25983_, _12441_, _06037_);
  nor _77231_ (_25984_, _25983_, _12700_);
  and _77232_ (_25985_, _25984_, _25981_);
  or _77233_ (_25986_, _25985_, _25827_);
  nand _77234_ (_25987_, _25986_, _25604_);
  and _77235_ (_25988_, _06401_, _06113_);
  nor _77236_ (_25989_, _25988_, _12696_);
  nand _77237_ (_25990_, _25989_, _25987_);
  nor _77238_ (_25991_, _06769_, _06004_);
  nor _77239_ (_25992_, _25991_, _12704_);
  and _77240_ (_25994_, _25992_, _25990_);
  nor _77241_ (_25995_, _25846_, _12705_);
  nor _77242_ (_25996_, _25995_, _25994_);
  and _77243_ (_25997_, _06785_, _06276_);
  or _77244_ (_25998_, _25997_, _25996_);
  and _77245_ (_25999_, _06466_, _06276_);
  and _77246_ (_26000_, _25997_, _06113_);
  nor _77247_ (_26001_, _26000_, _25999_);
  nand _77248_ (_26002_, _26001_, _25998_);
  and _77249_ (_26003_, _25999_, _06111_);
  not _77250_ (_26005_, _26003_);
  and _77251_ (_26006_, _26005_, _08625_);
  nand _77252_ (_26007_, _26006_, _26002_);
  nor _77253_ (_26008_, _08625_, _06111_);
  nor _77254_ (_26009_, _26008_, _06277_);
  nand _77255_ (_26010_, _26009_, _26007_);
  and _77256_ (_26011_, _12441_, _06277_);
  nor _77257_ (_26012_, _26011_, _11028_);
  and _77258_ (_26013_, _26012_, _26010_);
  and _77259_ (_26014_, _11028_, _06113_);
  or _77260_ (_26016_, _26014_, _26013_);
  nand _77261_ (_26017_, _26016_, _12719_);
  nor _77262_ (_26018_, _12719_, _06122_);
  nor _77263_ (_26019_, _26018_, _06400_);
  nand _77264_ (_26020_, _26019_, _26017_);
  and _77265_ (_26021_, _06400_, _06111_);
  nor _77266_ (_26022_, _26021_, _06275_);
  nand _77267_ (_26023_, _26022_, _26020_);
  and _77268_ (_26024_, _06769_, _06275_);
  nor _77269_ (_26025_, _26024_, _12763_);
  nand _77270_ (_26027_, _26025_, _26023_);
  nor _77271_ (_26028_, _25846_, _11389_);
  and _77272_ (_26029_, _11389_, _06113_);
  nor _77273_ (_26030_, _26029_, _12764_);
  not _77274_ (_26031_, _26030_);
  nor _77275_ (_26032_, _26031_, _26028_);
  nor _77276_ (_26033_, _26032_, _12768_);
  and _77277_ (_26034_, _26033_, _26027_);
  or _77278_ (_26035_, _26034_, _25826_);
  nand _77279_ (_26036_, _26035_, _12330_);
  nor _77280_ (_26038_, _12330_, _06111_);
  nor _77281_ (_26039_, _26038_, _06502_);
  nand _77282_ (_26040_, _26039_, _26036_);
  and _77283_ (_26041_, _12441_, _06502_);
  nor _77284_ (_26042_, _26041_, _06615_);
  and _77285_ (_26043_, _26042_, _26040_);
  and _77286_ (_26044_, _06615_, _06113_);
  or _77287_ (_26045_, _26044_, _26043_);
  nand _77288_ (_26046_, _26045_, _06012_);
  and _77289_ (_26047_, _06769_, _12782_);
  nor _77290_ (_26049_, _26047_, _12787_);
  nand _77291_ (_26050_, _26049_, _26046_);
  nor _77292_ (_26051_, _11389_, _06113_);
  and _77293_ (_26052_, _25846_, _11389_);
  or _77294_ (_26053_, _26052_, _26051_);
  and _77295_ (_26054_, _26053_, _12787_);
  nor _77296_ (_26055_, _26054_, _12792_);
  and _77297_ (_26056_, _26055_, _26050_);
  or _77298_ (_26057_, _26056_, _25825_);
  nand _77299_ (_26058_, _26057_, _12322_);
  nor _77300_ (_26060_, _12322_, _06111_);
  nor _77301_ (_26061_, _26060_, _06507_);
  nand _77302_ (_26062_, _26061_, _26058_);
  and _77303_ (_26063_, _12441_, _06507_);
  nor _77304_ (_26064_, _26063_, _06610_);
  and _77305_ (_26065_, _26064_, _26062_);
  and _77306_ (_26066_, _06610_, _06113_);
  or _77307_ (_26067_, _26066_, _26065_);
  nand _77308_ (_26068_, _26067_, _06018_);
  and _77309_ (_26069_, _06769_, _07330_);
  nor _77310_ (_26071_, _26069_, _12809_);
  nand _77311_ (_26072_, _26071_, _26068_);
  nor _77312_ (_26073_, _25846_, \oc8051_golden_model_1.PSW [7]);
  nor _77313_ (_26074_, _06111_, _10967_);
  nor _77314_ (_26075_, _26074_, _12810_);
  not _77315_ (_26076_, _26075_);
  nor _77316_ (_26077_, _26076_, _26073_);
  nor _77317_ (_26078_, _26077_, _12814_);
  and _77318_ (_26079_, _26078_, _26072_);
  or _77319_ (_26080_, _26079_, _25824_);
  nand _77320_ (_26082_, _26080_, _12314_);
  nor _77321_ (_26083_, _12314_, _06111_);
  nor _77322_ (_26084_, _26083_, _06509_);
  nand _77323_ (_26085_, _26084_, _26082_);
  and _77324_ (_26086_, _12441_, _06509_);
  nor _77325_ (_26087_, _26086_, _06602_);
  and _77326_ (_26088_, _26087_, _26085_);
  and _77327_ (_26089_, _06602_, _06113_);
  or _77328_ (_26090_, _26089_, _26088_);
  nand _77329_ (_26091_, _26090_, _06023_);
  and _77330_ (_26093_, _06769_, _12827_);
  nor _77331_ (_26094_, _26093_, _12310_);
  nand _77332_ (_26095_, _26094_, _26091_);
  and _77333_ (_26096_, _06111_, _10967_);
  and _77334_ (_26097_, _25846_, \oc8051_golden_model_1.PSW [7]);
  or _77335_ (_26098_, _26097_, _26096_);
  and _77336_ (_26099_, _26098_, _12310_);
  nor _77337_ (_26100_, _26099_, _12839_);
  and _77338_ (_26101_, _26100_, _26095_);
  or _77339_ (_26102_, _26101_, _25823_);
  nand _77340_ (_26104_, _26102_, _11187_);
  nor _77341_ (_26105_, _11187_, _06111_);
  nor _77342_ (_26106_, _26105_, _11216_);
  nand _77343_ (_26107_, _26106_, _26104_);
  and _77344_ (_26108_, _11216_, _06127_);
  nor _77345_ (_26109_, _26108_, _06621_);
  and _77346_ (_26110_, _26109_, _26107_);
  nor _77347_ (_26111_, _09356_, _14116_);
  or _77348_ (_26112_, _26111_, _26110_);
  nand _77349_ (_26113_, _26112_, _06016_);
  and _77350_ (_26115_, _06769_, _07350_);
  nor _77351_ (_26116_, _26115_, _06512_);
  nand _77352_ (_26117_, _26116_, _26113_);
  and _77353_ (_26118_, _25834_, _13037_);
  nor _77354_ (_26119_, _12441_, _13037_);
  or _77355_ (_26120_, _26119_, _06629_);
  or _77356_ (_26121_, _26120_, _26118_);
  and _77357_ (_26122_, _26121_, _12201_);
  and _77358_ (_26123_, _26122_, _26117_);
  or _77359_ (_26124_, _26123_, _25822_);
  nand _77360_ (_26126_, _26124_, _13046_);
  nor _77361_ (_26127_, _13046_, _06111_);
  nor _77362_ (_26128_, _26127_, _10564_);
  nand _77363_ (_26129_, _26128_, _26126_);
  and _77364_ (_26130_, _10564_, _06127_);
  nor _77365_ (_26131_, _26130_, _06361_);
  and _77366_ (_26132_, _26131_, _26129_);
  nor _77367_ (_26133_, _09356_, _06362_);
  or _77368_ (_26134_, _26133_, _26132_);
  nand _77369_ (_26135_, _26134_, _06021_);
  and _77370_ (_26137_, _06769_, _12187_);
  nor _77371_ (_26138_, _26137_, _06496_);
  nand _77372_ (_26139_, _26138_, _26135_);
  nor _77373_ (_26140_, _25833_, _13037_);
  and _77374_ (_26141_, _12442_, _13037_);
  nor _77375_ (_26142_, _26141_, _26140_);
  and _77376_ (_26143_, _26142_, _06496_);
  nor _77377_ (_26144_, _26143_, _13062_);
  nand _77378_ (_26145_, _26144_, _26139_);
  nor _77379_ (_26146_, _09123_, _06127_);
  nor _77380_ (_26148_, _26146_, _06639_);
  and _77381_ (_26149_, _26148_, _26145_);
  or _77382_ (_26150_, _26149_, _25821_);
  nand _77383_ (_26151_, _26150_, _13072_);
  nor _77384_ (_26152_, _13072_, _06128_);
  nor _77385_ (_26153_, _26152_, _07783_);
  nand _77386_ (_26154_, _26153_, _26151_);
  and _77387_ (_26155_, _07783_, _06769_);
  nor _77388_ (_26156_, _26155_, _05989_);
  nand _77389_ (_26157_, _26156_, _26154_);
  and _77390_ (_26159_, _26142_, _05989_);
  nor _77391_ (_26160_, _26159_, _13088_);
  nand _77392_ (_26161_, _26160_, _26157_);
  nor _77393_ (_26162_, _13087_, _06127_);
  nor _77394_ (_26163_, _26162_, _06646_);
  and _77395_ (_26164_, _26163_, _26161_);
  or _77396_ (_26165_, _26164_, _25820_);
  nand _77397_ (_26166_, _26165_, _13095_);
  nor _77398_ (_26167_, _13095_, _06128_);
  nor _77399_ (_26168_, _26167_, _25414_);
  nand _77400_ (_26170_, _26168_, _26166_);
  and _77401_ (_26171_, _25414_, _06769_);
  nor _77402_ (_26172_, _26171_, _13105_);
  and _77403_ (_26173_, _26172_, _26170_);
  and _77404_ (_26174_, _13105_, _06127_);
  or _77405_ (_26175_, _26174_, _26173_);
  or _77406_ (_26176_, _26175_, _01446_);
  or _77407_ (_26177_, _01442_, \oc8051_golden_model_1.PC [2]);
  and _77408_ (_26178_, _26177_, _43634_);
  and _77409_ (_44208_, _26178_, _26176_);
  and _77410_ (_26180_, _06646_, _06150_);
  and _77411_ (_26181_, _06639_, _06150_);
  nor _77412_ (_26182_, _12201_, _06173_);
  nor _77413_ (_26183_, _12837_, _06173_);
  nor _77414_ (_26184_, _12320_, _06173_);
  nor _77415_ (_26185_, _12328_, _06173_);
  nor _77416_ (_26186_, _12333_, _06173_);
  nor _77417_ (_26187_, _25555_, _06150_);
  and _77418_ (_26188_, _12347_, _06155_);
  or _77419_ (_26189_, _12510_, _12436_);
  or _77420_ (_26191_, _12439_, _12438_);
  and _77421_ (_26192_, _26191_, _12455_);
  nor _77422_ (_26193_, _26191_, _12455_);
  nor _77423_ (_26194_, _26193_, _26192_);
  or _77424_ (_26195_, _26194_, _12512_);
  and _77425_ (_26196_, _26195_, _26189_);
  or _77426_ (_26197_, _26196_, _07275_);
  and _77427_ (_26198_, _12539_, _06150_);
  or _77428_ (_26199_, _12257_, _12256_);
  and _77429_ (_26200_, _26199_, _12269_);
  nor _77430_ (_26202_, _26199_, _12269_);
  nor _77431_ (_26203_, _26202_, _26200_);
  and _77432_ (_26204_, _26203_, _12537_);
  nor _77433_ (_26205_, _26204_, _26198_);
  nand _77434_ (_26206_, _26205_, _08687_);
  nor _77435_ (_26207_, _12516_, _06173_);
  and _77436_ (_26208_, _12518_, _05661_);
  nor _77437_ (_26209_, _26208_, _07259_);
  and _77438_ (_26210_, _07259_, _06150_);
  nor _77439_ (_26211_, _26210_, _06855_);
  not _77440_ (_26213_, _26211_);
  nor _77441_ (_26214_, _26213_, _26209_);
  not _77442_ (_26215_, _26214_);
  nor _77443_ (_26216_, _12519_, _06173_);
  nor _77444_ (_26217_, _26216_, _06816_);
  and _77445_ (_26218_, _26217_, _26215_);
  nor _77446_ (_26219_, _07564_, _06595_);
  or _77447_ (_26220_, _26219_, _25207_);
  nor _77448_ (_26221_, _26220_, _26218_);
  nor _77449_ (_26222_, _26221_, _26207_);
  nor _77450_ (_26224_, _26222_, _08687_);
  nor _77451_ (_26225_, _26224_, _07269_);
  and _77452_ (_26226_, _26225_, _26206_);
  and _77453_ (_26227_, _07269_, _06173_);
  or _77454_ (_26228_, _26227_, _06474_);
  or _77455_ (_26229_, _26228_, _26226_);
  nand _77456_ (_26230_, _26229_, _26197_);
  nand _77457_ (_26231_, _26230_, _12502_);
  nor _77458_ (_26232_, _12502_, _06173_);
  nor _77459_ (_26233_, _26232_, _06356_);
  nand _77460_ (_26235_, _26233_, _26231_);
  and _77461_ (_26236_, _06356_, _06150_);
  nor _77462_ (_26237_, _26236_, _07692_);
  nand _77463_ (_26238_, _26237_, _26235_);
  and _77464_ (_26239_, _06595_, _07692_);
  nor _77465_ (_26240_, _26239_, _06410_);
  nand _77466_ (_26241_, _26240_, _26238_);
  and _77467_ (_26242_, _06410_, _06150_);
  nor _77468_ (_26243_, _26242_, _12552_);
  nand _77469_ (_26244_, _26243_, _26241_);
  nor _77470_ (_26246_, _12551_, _06173_);
  nor _77471_ (_26247_, _26246_, _06417_);
  nand _77472_ (_26248_, _26247_, _26244_);
  and _77473_ (_26249_, _06417_, _06150_);
  nor _77474_ (_26250_, _26249_, _12563_);
  nand _77475_ (_26251_, _26250_, _26248_);
  nor _77476_ (_26252_, _12561_, _06173_);
  nor _77477_ (_26253_, _26252_, _06352_);
  nand _77478_ (_26254_, _26253_, _26251_);
  and _77479_ (_26255_, _06352_, _06150_);
  nor _77480_ (_26257_, _26255_, _12565_);
  nand _77481_ (_26258_, _26257_, _26254_);
  and _77482_ (_26259_, _06595_, _12565_);
  nor _77483_ (_26260_, _26259_, _06351_);
  nand _77484_ (_26261_, _26260_, _26258_);
  and _77485_ (_26262_, _06351_, _06150_);
  nor _77486_ (_26263_, _26262_, _12611_);
  and _77487_ (_26264_, _26263_, _26261_);
  and _77488_ (_26265_, _12609_, _12436_);
  not _77489_ (_26266_, _26194_);
  nor _77490_ (_26268_, _26266_, _12609_);
  or _77491_ (_26269_, _26268_, _12574_);
  nor _77492_ (_26270_, _26269_, _26265_);
  or _77493_ (_26271_, _26270_, _26264_);
  nand _77494_ (_26272_, _26271_, _06473_);
  nor _77495_ (_26273_, _12437_, _12379_);
  and _77496_ (_26274_, _26194_, _12379_);
  nor _77497_ (_26275_, _26274_, _26273_);
  nand _77498_ (_26276_, _26275_, _06472_);
  and _77499_ (_26277_, _26276_, _06500_);
  nand _77500_ (_26279_, _26277_, _26272_);
  nor _77501_ (_26280_, _26194_, _12630_);
  and _77502_ (_26281_, _12630_, _12437_);
  or _77503_ (_26282_, _26281_, _06500_);
  or _77504_ (_26283_, _26282_, _26280_);
  nand _77505_ (_26284_, _26283_, _26279_);
  nand _77506_ (_26285_, _26284_, _12349_);
  nor _77507_ (_26286_, _26194_, _12648_);
  and _77508_ (_26287_, _12648_, _12437_);
  or _77509_ (_26288_, _26287_, _12349_);
  nor _77510_ (_26290_, _26288_, _26286_);
  nor _77511_ (_26291_, _26290_, _12347_);
  and _77512_ (_26292_, _26291_, _26285_);
  or _77513_ (_26293_, _26292_, _26188_);
  nand _77514_ (_26294_, _26293_, _06346_);
  and _77515_ (_26295_, _06345_, _06521_);
  nor _77516_ (_26296_, _26295_, _07596_);
  nand _77517_ (_26297_, _26296_, _26294_);
  nor _77518_ (_26298_, _06595_, _06049_);
  nor _77519_ (_26299_, _26298_, _25556_);
  and _77520_ (_26301_, _26299_, _26297_);
  or _77521_ (_26302_, _26301_, _26187_);
  nand _77522_ (_26303_, _26302_, _12344_);
  nor _77523_ (_26304_, _12344_, _06173_);
  nor _77524_ (_26305_, _26304_, _06445_);
  nand _77525_ (_26306_, _26305_, _26303_);
  and _77526_ (_26307_, _06445_, _06150_);
  nor _77527_ (_26308_, _26307_, _25285_);
  nand _77528_ (_26309_, _26308_, _26306_);
  and _77529_ (_26310_, _06595_, _25285_);
  nor _77530_ (_26312_, _26310_, _06444_);
  nand _77531_ (_26313_, _26312_, _26309_);
  and _77532_ (_26314_, _06444_, _06150_);
  nor _77533_ (_26315_, _26314_, _12671_);
  and _77534_ (_26316_, _26315_, _26313_);
  nor _77535_ (_26317_, _12339_, _06173_);
  or _77536_ (_26318_, _26317_, _26316_);
  nand _77537_ (_26319_, _26318_, _12336_);
  nor _77538_ (_26320_, _12336_, _06150_);
  nor _77539_ (_26321_, _26320_, _06042_);
  nand _77540_ (_26323_, _26321_, _26319_);
  and _77541_ (_26324_, _06042_, _06173_);
  nor _77542_ (_26325_, _26324_, _06339_);
  and _77543_ (_26326_, _26325_, _26323_);
  and _77544_ (_26327_, _06339_, _06521_);
  or _77545_ (_26328_, _26327_, _26326_);
  nand _77546_ (_26329_, _26328_, _07745_);
  and _77547_ (_26330_, _06595_, _06039_);
  nor _77548_ (_26331_, _26330_, _06486_);
  nand _77549_ (_26332_, _26331_, _26329_);
  and _77550_ (_26334_, _12436_, _06486_);
  nor _77551_ (_26335_, _26334_, _14022_);
  nand _77552_ (_26336_, _26335_, _26332_);
  nor _77553_ (_26337_, _06334_, _06150_);
  nor _77554_ (_26338_, _26337_, _06037_);
  nand _77555_ (_26339_, _26338_, _26336_);
  and _77556_ (_26340_, _12436_, _06037_);
  nor _77557_ (_26341_, _26340_, _12700_);
  nand _77558_ (_26342_, _26341_, _26339_);
  nor _77559_ (_26343_, _12694_, _06173_);
  nor _77560_ (_26345_, _26343_, _06401_);
  nand _77561_ (_26346_, _26345_, _26342_);
  and _77562_ (_26347_, _06401_, _06150_);
  nor _77563_ (_26348_, _26347_, _12696_);
  nand _77564_ (_26349_, _26348_, _26346_);
  and _77565_ (_26350_, _06595_, _12696_);
  nor _77566_ (_26351_, _26350_, _12704_);
  nand _77567_ (_26352_, _26351_, _26349_);
  and _77568_ (_26353_, _26203_, _12704_);
  nor _77569_ (_26354_, _26353_, _08848_);
  and _77570_ (_26356_, _26354_, _26352_);
  nor _77571_ (_26357_, _06277_, _06521_);
  nor _77572_ (_26358_, _26357_, _08627_);
  or _77573_ (_26359_, _26358_, _26356_);
  and _77574_ (_26360_, _12436_, _06277_);
  nor _77575_ (_26361_, _26360_, _11028_);
  and _77576_ (_26362_, _26361_, _26359_);
  and _77577_ (_26363_, _11028_, _06521_);
  or _77578_ (_26364_, _26363_, _26362_);
  nand _77579_ (_26365_, _26364_, _12719_);
  and _77580_ (_26367_, _12718_, _06171_);
  nor _77581_ (_26368_, _26367_, _06400_);
  nand _77582_ (_26369_, _26368_, _26365_);
  and _77583_ (_26370_, _06400_, _06150_);
  nor _77584_ (_26371_, _26370_, _06275_);
  nand _77585_ (_26372_, _26371_, _26369_);
  and _77586_ (_26373_, _06595_, _06275_);
  nor _77587_ (_26374_, _26373_, _12763_);
  nand _77588_ (_26375_, _26374_, _26372_);
  nor _77589_ (_26376_, _26203_, _11389_);
  and _77590_ (_26378_, _11389_, _06521_);
  nor _77591_ (_26379_, _26378_, _12764_);
  not _77592_ (_26380_, _26379_);
  nor _77593_ (_26381_, _26380_, _26376_);
  nor _77594_ (_26382_, _26381_, _12768_);
  and _77595_ (_26383_, _26382_, _26375_);
  or _77596_ (_26384_, _26383_, _26186_);
  nand _77597_ (_26385_, _26384_, _12330_);
  nor _77598_ (_26386_, _12330_, _06150_);
  nor _77599_ (_26387_, _26386_, _06502_);
  nand _77600_ (_26388_, _26387_, _26385_);
  and _77601_ (_26389_, _12436_, _06502_);
  nor _77602_ (_26390_, _26389_, _06615_);
  and _77603_ (_26391_, _26390_, _26388_);
  and _77604_ (_26392_, _06615_, _06521_);
  or _77605_ (_26393_, _26392_, _26391_);
  nand _77606_ (_26394_, _26393_, _06012_);
  and _77607_ (_26395_, _06595_, _12782_);
  nor _77608_ (_26396_, _26395_, _12787_);
  nand _77609_ (_26397_, _26396_, _26394_);
  nor _77610_ (_26400_, _11389_, _06521_);
  and _77611_ (_26401_, _26203_, _11389_);
  or _77612_ (_26402_, _26401_, _26400_);
  and _77613_ (_26403_, _26402_, _12787_);
  nor _77614_ (_26404_, _26403_, _12792_);
  and _77615_ (_26405_, _26404_, _26397_);
  or _77616_ (_26406_, _26405_, _26185_);
  nand _77617_ (_26407_, _26406_, _12322_);
  nor _77618_ (_26408_, _12322_, _06150_);
  nor _77619_ (_26409_, _26408_, _06507_);
  nand _77620_ (_26411_, _26409_, _26407_);
  and _77621_ (_26412_, _12436_, _06507_);
  nor _77622_ (_26413_, _26412_, _06610_);
  and _77623_ (_26414_, _26413_, _26411_);
  and _77624_ (_26415_, _06610_, _06521_);
  or _77625_ (_26416_, _26415_, _26414_);
  nand _77626_ (_26417_, _26416_, _06018_);
  and _77627_ (_26418_, _06595_, _07330_);
  nor _77628_ (_26419_, _26418_, _12809_);
  nand _77629_ (_26420_, _26419_, _26417_);
  and _77630_ (_26422_, _06150_, \oc8051_golden_model_1.PSW [7]);
  and _77631_ (_26423_, _26203_, _10967_);
  or _77632_ (_26424_, _26423_, _26422_);
  and _77633_ (_26425_, _26424_, _12809_);
  nor _77634_ (_26426_, _26425_, _12814_);
  and _77635_ (_26427_, _26426_, _26420_);
  or _77636_ (_26428_, _26427_, _26184_);
  nand _77637_ (_26429_, _26428_, _12314_);
  nor _77638_ (_26430_, _12314_, _06150_);
  nor _77639_ (_26431_, _26430_, _06509_);
  nand _77640_ (_26433_, _26431_, _26429_);
  and _77641_ (_26434_, _12436_, _06509_);
  nor _77642_ (_26435_, _26434_, _06602_);
  and _77643_ (_26436_, _26435_, _26433_);
  and _77644_ (_26437_, _06602_, _06521_);
  or _77645_ (_26438_, _26437_, _26436_);
  nand _77646_ (_26439_, _26438_, _06023_);
  and _77647_ (_26440_, _06595_, _12827_);
  nor _77648_ (_26441_, _26440_, _12310_);
  nand _77649_ (_26442_, _26441_, _26439_);
  and _77650_ (_26444_, _06150_, _10967_);
  and _77651_ (_26445_, _26203_, \oc8051_golden_model_1.PSW [7]);
  or _77652_ (_26446_, _26445_, _26444_);
  and _77653_ (_26447_, _26446_, _12310_);
  nor _77654_ (_26448_, _26447_, _12839_);
  and _77655_ (_26449_, _26448_, _26442_);
  or _77656_ (_26450_, _26449_, _26183_);
  nand _77657_ (_26451_, _26450_, _11187_);
  nor _77658_ (_26452_, _11187_, _06150_);
  nor _77659_ (_26453_, _26452_, _11216_);
  nand _77660_ (_26455_, _26453_, _26451_);
  and _77661_ (_26456_, _11216_, _06173_);
  nor _77662_ (_26457_, _26456_, _06621_);
  and _77663_ (_26458_, _26457_, _26455_);
  nor _77664_ (_26459_, _09310_, _14116_);
  or _77665_ (_26460_, _26459_, _26458_);
  nand _77666_ (_26461_, _26460_, _06016_);
  and _77667_ (_26462_, _06595_, _07350_);
  nor _77668_ (_26463_, _26462_, _06512_);
  nand _77669_ (_26464_, _26463_, _26461_);
  and _77670_ (_26466_, _26266_, _13037_);
  nor _77671_ (_26467_, _12436_, _13037_);
  or _77672_ (_26468_, _26467_, _06629_);
  or _77673_ (_26469_, _26468_, _26466_);
  and _77674_ (_26470_, _26469_, _12201_);
  and _77675_ (_26471_, _26470_, _26464_);
  or _77676_ (_26472_, _26471_, _26182_);
  nand _77677_ (_26473_, _26472_, _13046_);
  nor _77678_ (_26474_, _13046_, _06150_);
  nor _77679_ (_26475_, _26474_, _10564_);
  nand _77680_ (_26477_, _26475_, _26473_);
  and _77681_ (_26478_, _10564_, _06173_);
  nor _77682_ (_26479_, _26478_, _06361_);
  and _77683_ (_26480_, _26479_, _26477_);
  nor _77684_ (_26481_, _09310_, _06362_);
  or _77685_ (_26482_, _26481_, _26480_);
  nand _77686_ (_26483_, _26482_, _06021_);
  and _77687_ (_26484_, _06595_, _12187_);
  nor _77688_ (_26485_, _26484_, _06496_);
  nand _77689_ (_26486_, _26485_, _26483_);
  nor _77690_ (_26488_, _26194_, _13037_);
  and _77691_ (_26489_, _12437_, _13037_);
  nor _77692_ (_26490_, _26489_, _26488_);
  and _77693_ (_26491_, _26490_, _06496_);
  nor _77694_ (_26492_, _26491_, _13062_);
  nand _77695_ (_26493_, _26492_, _26486_);
  nor _77696_ (_26494_, _09123_, _06173_);
  nor _77697_ (_26495_, _26494_, _06639_);
  and _77698_ (_26496_, _26495_, _26493_);
  or _77699_ (_26497_, _26496_, _26181_);
  nand _77700_ (_26499_, _26497_, _13072_);
  nor _77701_ (_26500_, _13072_, _06155_);
  nor _77702_ (_26501_, _26500_, _07783_);
  nand _77703_ (_26502_, _26501_, _26499_);
  and _77704_ (_26503_, _07783_, _06595_);
  nor _77705_ (_26504_, _26503_, _05989_);
  nand _77706_ (_26505_, _26504_, _26502_);
  and _77707_ (_26506_, _26490_, _05989_);
  nor _77708_ (_26507_, _26506_, _13088_);
  nand _77709_ (_26508_, _26507_, _26505_);
  nor _77710_ (_26510_, _13087_, _06173_);
  nor _77711_ (_26511_, _26510_, _06646_);
  and _77712_ (_26512_, _26511_, _26508_);
  or _77713_ (_26513_, _26512_, _26180_);
  nand _77714_ (_26514_, _26513_, _13095_);
  nor _77715_ (_26515_, _13095_, _06155_);
  nor _77716_ (_26516_, _26515_, _25414_);
  nand _77717_ (_26517_, _26516_, _26514_);
  and _77718_ (_26518_, _25414_, _06595_);
  nor _77719_ (_26519_, _26518_, _13105_);
  and _77720_ (_26521_, _26519_, _26517_);
  and _77721_ (_26522_, _13105_, _06173_);
  or _77722_ (_26523_, _26522_, _26521_);
  or _77723_ (_26524_, _26523_, _01446_);
  or _77724_ (_26525_, _01442_, \oc8051_golden_model_1.PC [3]);
  and _77725_ (_26526_, _26525_, _43634_);
  and _77726_ (_44210_, _26526_, _26524_);
  nor _77727_ (_26527_, _12254_, _11389_);
  and _77728_ (_26528_, _12274_, _12271_);
  nor _77729_ (_26529_, _26528_, _12275_);
  and _77730_ (_26531_, _26529_, _11389_);
  or _77731_ (_26532_, _26531_, _26527_);
  and _77732_ (_26533_, _26532_, _12787_);
  and _77733_ (_26534_, _08986_, _25285_);
  nor _77734_ (_26535_, _25555_, _12253_);
  not _77735_ (_26536_, \oc8051_golden_model_1.PC [4]);
  nor _77736_ (_26537_, _05685_, _26536_);
  and _77737_ (_26538_, _05685_, _26536_);
  nor _77738_ (_26539_, _26538_, _26537_);
  not _77739_ (_26540_, _26539_);
  and _77740_ (_26542_, _26540_, _12347_);
  and _77741_ (_26543_, _12253_, _06351_);
  and _77742_ (_26544_, _12254_, _06352_);
  and _77743_ (_26545_, _12460_, _12457_);
  nor _77744_ (_26546_, _26545_, _12461_);
  or _77745_ (_26547_, _26546_, _12512_);
  or _77746_ (_26548_, _12510_, _12432_);
  and _77747_ (_26549_, _26548_, _26547_);
  or _77748_ (_26550_, _26549_, _07275_);
  nand _77749_ (_26551_, _26529_, _12537_);
  or _77750_ (_26553_, _12537_, _12254_);
  and _77751_ (_26554_, _26553_, _26551_);
  nand _77752_ (_26555_, _26554_, _08687_);
  and _77753_ (_26556_, _08986_, _06816_);
  nand _77754_ (_26557_, _12518_, \oc8051_golden_model_1.PC [4]);
  and _77755_ (_26558_, _26557_, _07260_);
  and _77756_ (_26559_, _12254_, _07259_);
  or _77757_ (_26560_, _26559_, _06855_);
  or _77758_ (_26561_, _26560_, _26558_);
  or _77759_ (_26562_, _26540_, _12519_);
  and _77760_ (_26564_, _26562_, _07564_);
  and _77761_ (_26565_, _26564_, _26561_);
  nor _77762_ (_26566_, _26565_, _25207_);
  not _77763_ (_26567_, _26566_);
  nor _77764_ (_26568_, _26567_, _26556_);
  nor _77765_ (_26569_, _26540_, _12516_);
  nor _77766_ (_26570_, _26569_, _08687_);
  not _77767_ (_26571_, _26570_);
  nor _77768_ (_26572_, _26571_, _26568_);
  nor _77769_ (_26573_, _26572_, _07269_);
  and _77770_ (_26575_, _26573_, _26555_);
  and _77771_ (_26576_, _26539_, _07269_);
  or _77772_ (_26577_, _26576_, _06474_);
  or _77773_ (_26578_, _26577_, _26575_);
  and _77774_ (_26579_, _26578_, _12502_);
  and _77775_ (_26580_, _26579_, _26550_);
  nor _77776_ (_26581_, _26540_, _12502_);
  or _77777_ (_26582_, _26581_, _06356_);
  or _77778_ (_26583_, _26582_, _26580_);
  and _77779_ (_26584_, _12254_, _06356_);
  nor _77780_ (_26586_, _26584_, _07692_);
  nand _77781_ (_26587_, _26586_, _26583_);
  nor _77782_ (_26588_, _08986_, _06052_);
  nor _77783_ (_26589_, _26588_, _06410_);
  and _77784_ (_26590_, _26589_, _26587_);
  and _77785_ (_26591_, _12254_, _06410_);
  or _77786_ (_26592_, _26591_, _26590_);
  and _77787_ (_26593_, _26592_, _12551_);
  nor _77788_ (_26594_, _26539_, _12551_);
  or _77789_ (_26595_, _26594_, _26593_);
  nand _77790_ (_26597_, _26595_, _06426_);
  and _77791_ (_26598_, _12254_, _06417_);
  nor _77792_ (_26599_, _26598_, _12563_);
  nand _77793_ (_26600_, _26599_, _26597_);
  nor _77794_ (_26601_, _26540_, _12561_);
  nor _77795_ (_26602_, _26601_, _06352_);
  and _77796_ (_26603_, _26602_, _26600_);
  or _77797_ (_26604_, _26603_, _26544_);
  nand _77798_ (_26605_, _26604_, _06057_);
  and _77799_ (_26606_, _08986_, _12565_);
  nor _77800_ (_26608_, _26606_, _06351_);
  nand _77801_ (_26609_, _26608_, _26605_);
  nand _77802_ (_26610_, _26609_, _12573_);
  nor _77803_ (_26611_, _26610_, _26543_);
  and _77804_ (_26612_, _12609_, _12433_);
  nor _77805_ (_26613_, _26546_, _12609_);
  nor _77806_ (_26614_, _26613_, _26612_);
  and _77807_ (_26615_, _26614_, _12571_);
  nor _77808_ (_26616_, _26615_, _12574_);
  or _77809_ (_26617_, _26616_, _26611_);
  and _77810_ (_26618_, _26614_, _06469_);
  nor _77811_ (_26619_, _26618_, _06472_);
  nand _77812_ (_26620_, _26619_, _26617_);
  nor _77813_ (_26621_, _12433_, _12379_);
  and _77814_ (_26622_, _26546_, _12379_);
  or _77815_ (_26623_, _26622_, _06473_);
  nor _77816_ (_26624_, _26623_, _26621_);
  nor _77817_ (_26625_, _26624_, _06431_);
  nand _77818_ (_26626_, _26625_, _26620_);
  and _77819_ (_26627_, _12630_, _12433_);
  nor _77820_ (_26630_, _26546_, _12630_);
  or _77821_ (_26631_, _26630_, _06500_);
  or _77822_ (_26632_, _26631_, _26627_);
  nand _77823_ (_26633_, _26632_, _26626_);
  nand _77824_ (_26634_, _26633_, _12349_);
  and _77825_ (_26635_, _12648_, _12432_);
  not _77826_ (_26636_, _12648_);
  and _77827_ (_26637_, _26546_, _26636_);
  or _77828_ (_26638_, _26637_, _26635_);
  and _77829_ (_26639_, _26638_, _06490_);
  nor _77830_ (_26641_, _26639_, _12347_);
  and _77831_ (_26642_, _26641_, _26634_);
  or _77832_ (_26643_, _26642_, _26542_);
  nand _77833_ (_26644_, _26643_, _06346_);
  and _77834_ (_26645_, _12254_, _06345_);
  nor _77835_ (_26646_, _26645_, _07596_);
  nand _77836_ (_26647_, _26646_, _26644_);
  nor _77837_ (_26648_, _08986_, _06049_);
  nor _77838_ (_26649_, _26648_, _25556_);
  and _77839_ (_26650_, _26649_, _26647_);
  or _77840_ (_26652_, _26650_, _26535_);
  nand _77841_ (_26653_, _26652_, _12344_);
  nor _77842_ (_26654_, _26539_, _12344_);
  nor _77843_ (_26655_, _26654_, _06445_);
  nand _77844_ (_26656_, _26655_, _26653_);
  and _77845_ (_26657_, _12253_, _06445_);
  nor _77846_ (_26658_, _26657_, _25285_);
  and _77847_ (_26659_, _26658_, _26656_);
  or _77848_ (_26660_, _26659_, _26534_);
  nand _77849_ (_26661_, _26660_, _14251_);
  and _77850_ (_26663_, _12254_, _06444_);
  nor _77851_ (_26664_, _26663_, _12671_);
  nand _77852_ (_26665_, _26664_, _26661_);
  nor _77853_ (_26666_, _26540_, _12339_);
  nor _77854_ (_26667_, _26666_, _12337_);
  nand _77855_ (_26668_, _26667_, _26665_);
  nor _77856_ (_26669_, _12253_, _12336_);
  nor _77857_ (_26670_, _26669_, _06042_);
  nand _77858_ (_26671_, _26670_, _26668_);
  and _77859_ (_26672_, _26539_, _06042_);
  nor _77860_ (_26674_, _26672_, _06339_);
  and _77861_ (_26675_, _26674_, _26671_);
  and _77862_ (_26676_, _12254_, _06339_);
  or _77863_ (_26677_, _26676_, _26675_);
  nand _77864_ (_26678_, _26677_, _07745_);
  and _77865_ (_26679_, _08986_, _06039_);
  nor _77866_ (_26680_, _26679_, _06486_);
  nand _77867_ (_26681_, _26680_, _26678_);
  and _77868_ (_26682_, _12432_, _06486_);
  nor _77869_ (_26683_, _26682_, _14022_);
  and _77870_ (_26685_, _26683_, _26681_);
  nor _77871_ (_26686_, _12253_, _06334_);
  or _77872_ (_26687_, _26686_, _26685_);
  nand _77873_ (_26688_, _26687_, _06313_);
  and _77874_ (_26689_, _12433_, _06037_);
  nor _77875_ (_26690_, _26689_, _12700_);
  nand _77876_ (_26691_, _26690_, _26688_);
  nor _77877_ (_26692_, _26540_, _12694_);
  nor _77878_ (_26693_, _26692_, _06401_);
  and _77879_ (_26694_, _26693_, _26691_);
  and _77880_ (_26696_, _12254_, _06401_);
  or _77881_ (_26697_, _26696_, _26694_);
  nand _77882_ (_26698_, _26697_, _06004_);
  and _77883_ (_26699_, _08986_, _12696_);
  nor _77884_ (_26700_, _26699_, _12704_);
  nand _77885_ (_26701_, _26700_, _26698_);
  and _77886_ (_26702_, _26529_, _12704_);
  nor _77887_ (_26703_, _26702_, _08848_);
  and _77888_ (_26704_, _26703_, _26701_);
  nor _77889_ (_26705_, _12254_, _06277_);
  nor _77890_ (_26707_, _26705_, _08627_);
  or _77891_ (_26708_, _26707_, _26704_);
  and _77892_ (_26709_, _12432_, _06277_);
  nor _77893_ (_26710_, _26709_, _11028_);
  nand _77894_ (_26711_, _26710_, _26708_);
  and _77895_ (_26712_, _12254_, _11028_);
  nor _77896_ (_26713_, _26712_, _12718_);
  nand _77897_ (_26714_, _26713_, _26711_);
  and _77898_ (_26715_, _12741_, _12738_);
  nor _77899_ (_26716_, _26715_, _12742_);
  and _77900_ (_26718_, _26716_, _12718_);
  nor _77901_ (_26719_, _26718_, _06400_);
  and _77902_ (_26720_, _26719_, _26714_);
  and _77903_ (_26721_, _12254_, _06400_);
  or _77904_ (_26722_, _26721_, _26720_);
  nand _77905_ (_26723_, _26722_, _06009_);
  and _77906_ (_26724_, _08986_, _06275_);
  nor _77907_ (_26725_, _26724_, _12763_);
  nand _77908_ (_26726_, _26725_, _26723_);
  nand _77909_ (_26727_, _12253_, _11389_);
  nand _77910_ (_26729_, _26529_, _12770_);
  and _77911_ (_26730_, _26729_, _26727_);
  or _77912_ (_26731_, _26730_, _12764_);
  nand _77913_ (_26732_, _26731_, _26726_);
  nand _77914_ (_26733_, _26732_, _12333_);
  nor _77915_ (_26734_, _26540_, _12333_);
  nor _77916_ (_26735_, _26734_, _12331_);
  nand _77917_ (_26736_, _26735_, _26733_);
  nor _77918_ (_26737_, _12253_, _12330_);
  nor _77919_ (_26738_, _26737_, _06502_);
  nand _77920_ (_26740_, _26738_, _26736_);
  and _77921_ (_26741_, _12432_, _06502_);
  nor _77922_ (_26742_, _26741_, _06615_);
  and _77923_ (_26743_, _26742_, _26740_);
  and _77924_ (_26744_, _12254_, _06615_);
  or _77925_ (_26745_, _26744_, _26743_);
  nand _77926_ (_26746_, _26745_, _06012_);
  and _77927_ (_26747_, _08986_, _12782_);
  nor _77928_ (_26748_, _26747_, _12787_);
  and _77929_ (_26749_, _26748_, _26746_);
  or _77930_ (_26751_, _26749_, _26533_);
  nand _77931_ (_26752_, _26751_, _12328_);
  nor _77932_ (_26753_, _26540_, _12328_);
  nor _77933_ (_26754_, _26753_, _12323_);
  nand _77934_ (_26755_, _26754_, _26752_);
  nor _77935_ (_26756_, _12253_, _12322_);
  nor _77936_ (_26757_, _26756_, _06507_);
  nand _77937_ (_26758_, _26757_, _26755_);
  and _77938_ (_26759_, _12432_, _06507_);
  nor _77939_ (_26760_, _26759_, _06610_);
  and _77940_ (_26762_, _26760_, _26758_);
  and _77941_ (_26763_, _12254_, _06610_);
  or _77942_ (_26764_, _26763_, _26762_);
  nand _77943_ (_26765_, _26764_, _06018_);
  and _77944_ (_26766_, _08986_, _07330_);
  nor _77945_ (_26767_, _26766_, _12809_);
  nand _77946_ (_26768_, _26767_, _26765_);
  nand _77947_ (_26769_, _12253_, \oc8051_golden_model_1.PSW [7]);
  nand _77948_ (_26770_, _26529_, _10967_);
  and _77949_ (_26771_, _26770_, _26769_);
  or _77950_ (_26773_, _26771_, _12810_);
  nand _77951_ (_26774_, _26773_, _26768_);
  nand _77952_ (_26775_, _26774_, _12320_);
  nor _77953_ (_26776_, _26540_, _12320_);
  nor _77954_ (_26777_, _26776_, _12315_);
  nand _77955_ (_26778_, _26777_, _26775_);
  nor _77956_ (_26779_, _12253_, _12314_);
  nor _77957_ (_26780_, _26779_, _06509_);
  nand _77958_ (_26781_, _26780_, _26778_);
  and _77959_ (_26782_, _12432_, _06509_);
  nor _77960_ (_26784_, _26782_, _06602_);
  and _77961_ (_26785_, _26784_, _26781_);
  and _77962_ (_26786_, _12254_, _06602_);
  or _77963_ (_26787_, _26786_, _26785_);
  nand _77964_ (_26788_, _26787_, _06023_);
  and _77965_ (_26789_, _08986_, _12827_);
  nor _77966_ (_26790_, _26789_, _12310_);
  nand _77967_ (_26791_, _26790_, _26788_);
  nand _77968_ (_26792_, _12253_, _10967_);
  nand _77969_ (_26793_, _26529_, \oc8051_golden_model_1.PSW [7]);
  and _77970_ (_26795_, _26793_, _26792_);
  or _77971_ (_26796_, _26795_, _12832_);
  nand _77972_ (_26797_, _26796_, _26791_);
  nand _77973_ (_26798_, _26797_, _12837_);
  nor _77974_ (_26799_, _26540_, _12837_);
  nor _77975_ (_26800_, _26799_, _11188_);
  nand _77976_ (_26801_, _26800_, _26798_);
  nor _77977_ (_26802_, _12253_, _11187_);
  nor _77978_ (_26803_, _26802_, _11216_);
  nand _77979_ (_26804_, _26803_, _26801_);
  and _77980_ (_26806_, _26539_, _11216_);
  nor _77981_ (_26807_, _26806_, _06621_);
  and _77982_ (_26808_, _26807_, _26804_);
  nor _77983_ (_26809_, _09264_, _14116_);
  or _77984_ (_26810_, _26809_, _26808_);
  nand _77985_ (_26811_, _26810_, _06016_);
  and _77986_ (_26812_, _08986_, _07350_);
  nor _77987_ (_26813_, _26812_, _06512_);
  and _77988_ (_26814_, _26813_, _26811_);
  nor _77989_ (_26815_, _12433_, _13037_);
  and _77990_ (_26817_, _26546_, _13037_);
  nor _77991_ (_26818_, _26817_, _26815_);
  nor _77992_ (_26819_, _26818_, _06629_);
  or _77993_ (_26820_, _26819_, _26814_);
  nand _77994_ (_26821_, _26820_, _12201_);
  nor _77995_ (_26822_, _26540_, _12201_);
  nor _77996_ (_26823_, _26822_, _13047_);
  nand _77997_ (_26824_, _26823_, _26821_);
  nor _77998_ (_26825_, _13046_, _12253_);
  nor _77999_ (_26826_, _26825_, _10564_);
  nand _78000_ (_26828_, _26826_, _26824_);
  and _78001_ (_26829_, _26539_, _10564_);
  nor _78002_ (_26830_, _26829_, _06361_);
  nand _78003_ (_26831_, _26830_, _26828_);
  nor _78004_ (_26832_, _09264_, _06362_);
  nor _78005_ (_26833_, _26832_, _12187_);
  nand _78006_ (_26834_, _26833_, _26831_);
  nor _78007_ (_26835_, _08986_, _06021_);
  nor _78008_ (_26836_, _26835_, _06496_);
  nand _78009_ (_26837_, _26836_, _26834_);
  and _78010_ (_26839_, _12433_, _13037_);
  nor _78011_ (_26840_, _26546_, _13037_);
  nor _78012_ (_26841_, _26840_, _26839_);
  nor _78013_ (_26842_, _26841_, _07035_);
  nor _78014_ (_26843_, _26842_, _13062_);
  nand _78015_ (_26844_, _26843_, _26837_);
  nor _78016_ (_26845_, _26540_, _09123_);
  nor _78017_ (_26846_, _26845_, _06639_);
  nand _78018_ (_26847_, _26846_, _26844_);
  not _78019_ (_26848_, _13072_);
  and _78020_ (_26850_, _12254_, _06639_);
  nor _78021_ (_26851_, _26850_, _26848_);
  nand _78022_ (_26852_, _26851_, _26847_);
  nor _78023_ (_26853_, _26540_, _13072_);
  nor _78024_ (_26854_, _26853_, _07783_);
  nand _78025_ (_26855_, _26854_, _26852_);
  and _78026_ (_26856_, _08986_, _07783_);
  nor _78027_ (_26857_, _26856_, _05989_);
  nand _78028_ (_26858_, _26857_, _26855_);
  and _78029_ (_26859_, _26841_, _05989_);
  nor _78030_ (_26861_, _26859_, _13088_);
  and _78031_ (_26862_, _26861_, _26858_);
  nor _78032_ (_26863_, _26539_, _13087_);
  or _78033_ (_26864_, _26863_, _26862_);
  nand _78034_ (_26865_, _26864_, _06651_);
  not _78035_ (_26866_, _13095_);
  and _78036_ (_26867_, _12254_, _06646_);
  nor _78037_ (_26868_, _26867_, _26866_);
  nand _78038_ (_26869_, _26868_, _26865_);
  nor _78039_ (_26870_, _26540_, _13095_);
  nor _78040_ (_26872_, _26870_, _25414_);
  nand _78041_ (_26873_, _26872_, _26869_);
  and _78042_ (_26874_, _25414_, _08986_);
  nor _78043_ (_26875_, _26874_, _13105_);
  and _78044_ (_26876_, _26875_, _26873_);
  and _78045_ (_26877_, _26539_, _13105_);
  or _78046_ (_26878_, _26877_, _26876_);
  or _78047_ (_26879_, _26878_, _01446_);
  or _78048_ (_26880_, _01442_, \oc8051_golden_model_1.PC [4]);
  and _78049_ (_26881_, _26880_, _43634_);
  and _78050_ (_44211_, _26881_, _26879_);
  and _78051_ (_26883_, _12248_, _06646_);
  nor _78052_ (_26884_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _78053_ (_26885_, _12248_, _05701_);
  nor _78054_ (_26886_, _26885_, _26884_);
  nor _78055_ (_26887_, _26886_, _12201_);
  nor _78056_ (_26888_, _26886_, _12837_);
  nor _78057_ (_26889_, _26886_, _12320_);
  nor _78058_ (_26890_, _26886_, _12328_);
  nor _78059_ (_26891_, _26886_, _12333_);
  and _78060_ (_26893_, _12249_, _06400_);
  nor _78061_ (_26894_, _25555_, _12248_);
  or _78062_ (_26895_, _12428_, _12379_);
  or _78063_ (_26896_, _12430_, _12429_);
  not _78064_ (_26897_, _26896_);
  nor _78065_ (_26898_, _26897_, _12462_);
  and _78066_ (_26899_, _26897_, _12462_);
  nor _78067_ (_26900_, _26899_, _26898_);
  not _78068_ (_26901_, _26900_);
  nand _78069_ (_26902_, _26901_, _12379_);
  and _78070_ (_26904_, _26902_, _06472_);
  nand _78071_ (_26905_, _26904_, _26895_);
  and _78072_ (_26906_, _12609_, _12428_);
  nor _78073_ (_26907_, _26901_, _12609_);
  nor _78074_ (_26908_, _26907_, _26906_);
  and _78075_ (_26909_, _26908_, _06469_);
  and _78076_ (_26910_, _12248_, _06351_);
  or _78077_ (_26911_, _12510_, _12427_);
  or _78078_ (_26912_, _26901_, _12512_);
  and _78079_ (_26913_, _26912_, _26911_);
  or _78080_ (_26915_, _26913_, _07275_);
  and _78081_ (_26916_, _12539_, _12248_);
  or _78082_ (_26917_, _12251_, _12250_);
  not _78083_ (_26918_, _26917_);
  nor _78084_ (_26919_, _26918_, _12276_);
  and _78085_ (_26920_, _26918_, _12276_);
  nor _78086_ (_26921_, _26920_, _26919_);
  nor _78087_ (_26922_, _26921_, _12539_);
  nor _78088_ (_26923_, _26922_, _26916_);
  nand _78089_ (_26924_, _26923_, _08687_);
  nor _78090_ (_26926_, _26886_, _12516_);
  not _78091_ (_26927_, _12518_);
  nor _78092_ (_26928_, _26927_, \oc8051_golden_model_1.PC [5]);
  nor _78093_ (_26929_, _26928_, _07259_);
  and _78094_ (_26930_, _12248_, _07259_);
  nor _78095_ (_26931_, _26930_, _06855_);
  not _78096_ (_26932_, _26931_);
  nor _78097_ (_26933_, _26932_, _26929_);
  nor _78098_ (_26934_, _26886_, _12519_);
  nor _78099_ (_26935_, _26934_, _06816_);
  not _78100_ (_26937_, _26935_);
  nor _78101_ (_26938_, _26937_, _26933_);
  nor _78102_ (_26939_, _08953_, _07564_);
  or _78103_ (_26940_, _26939_, _25207_);
  nor _78104_ (_26941_, _26940_, _26938_);
  nor _78105_ (_26942_, _26941_, _26926_);
  nor _78106_ (_26943_, _26942_, _08687_);
  nor _78107_ (_26944_, _26943_, _07269_);
  and _78108_ (_26945_, _26944_, _26924_);
  and _78109_ (_26946_, _26886_, _07269_);
  or _78110_ (_26948_, _26946_, _06474_);
  or _78111_ (_26949_, _26948_, _26945_);
  nand _78112_ (_26950_, _26949_, _26915_);
  nand _78113_ (_26951_, _26950_, _12502_);
  nor _78114_ (_26952_, _26886_, _12502_);
  nor _78115_ (_26953_, _26952_, _06356_);
  nand _78116_ (_26954_, _26953_, _26951_);
  and _78117_ (_26955_, _12248_, _06356_);
  nor _78118_ (_26956_, _26955_, _07692_);
  nand _78119_ (_26957_, _26956_, _26954_);
  and _78120_ (_26959_, _08953_, _07692_);
  nor _78121_ (_26960_, _26959_, _06410_);
  nand _78122_ (_26961_, _26960_, _26957_);
  and _78123_ (_26962_, _12248_, _06410_);
  nor _78124_ (_26963_, _26962_, _12552_);
  nand _78125_ (_26964_, _26963_, _26961_);
  nor _78126_ (_26965_, _26886_, _12551_);
  nor _78127_ (_26966_, _26965_, _06417_);
  nand _78128_ (_26967_, _26966_, _26964_);
  and _78129_ (_26968_, _12248_, _06417_);
  nor _78130_ (_26970_, _26968_, _12563_);
  nand _78131_ (_26971_, _26970_, _26967_);
  nor _78132_ (_26972_, _26886_, _12561_);
  nor _78133_ (_26973_, _26972_, _06352_);
  nand _78134_ (_26974_, _26973_, _26971_);
  and _78135_ (_26975_, _12248_, _06352_);
  nor _78136_ (_26976_, _26975_, _12565_);
  nand _78137_ (_26977_, _26976_, _26974_);
  and _78138_ (_26978_, _08953_, _12565_);
  nor _78139_ (_26979_, _26978_, _06351_);
  nand _78140_ (_26981_, _26979_, _26977_);
  nand _78141_ (_26982_, _26981_, _12573_);
  or _78142_ (_26983_, _26982_, _26910_);
  nor _78143_ (_26984_, _26983_, _26909_);
  nor _78144_ (_26985_, _26908_, _12574_);
  or _78145_ (_26986_, _26985_, _26984_);
  nand _78146_ (_26987_, _26986_, _06473_);
  and _78147_ (_26988_, _26987_, _26905_);
  or _78148_ (_26989_, _26988_, _06431_);
  and _78149_ (_26990_, _12630_, _12427_);
  nor _78150_ (_26992_, _26900_, _12630_);
  or _78151_ (_26993_, _26992_, _06500_);
  or _78152_ (_26994_, _26993_, _26990_);
  and _78153_ (_26995_, _26994_, _12349_);
  nand _78154_ (_26996_, _26995_, _26989_);
  nand _78155_ (_26997_, _12648_, _12427_);
  or _78156_ (_26998_, _26900_, _12648_);
  and _78157_ (_26999_, _26998_, _26997_);
  or _78158_ (_27000_, _26999_, _12349_);
  and _78159_ (_27001_, _27000_, _26996_);
  or _78160_ (_27003_, _27001_, _12347_);
  nand _78161_ (_27004_, _26886_, _12347_);
  and _78162_ (_27005_, _27004_, _27003_);
  nand _78163_ (_27006_, _27005_, _06346_);
  and _78164_ (_27007_, _12249_, _06345_);
  nor _78165_ (_27008_, _27007_, _07596_);
  nand _78166_ (_27009_, _27008_, _27006_);
  nor _78167_ (_27010_, _08953_, _06049_);
  nor _78168_ (_27011_, _27010_, _25556_);
  and _78169_ (_27012_, _27011_, _27009_);
  or _78170_ (_27014_, _27012_, _26894_);
  nand _78171_ (_27015_, _27014_, _12344_);
  nor _78172_ (_27016_, _26886_, _12344_);
  nor _78173_ (_27017_, _27016_, _06445_);
  nand _78174_ (_27018_, _27017_, _27015_);
  and _78175_ (_27019_, _12248_, _06445_);
  nor _78176_ (_27020_, _27019_, _25285_);
  nand _78177_ (_27021_, _27020_, _27018_);
  and _78178_ (_27022_, _08953_, _25285_);
  nor _78179_ (_27023_, _27022_, _06444_);
  nand _78180_ (_27025_, _27023_, _27021_);
  and _78181_ (_27026_, _12248_, _06444_);
  nor _78182_ (_27027_, _27026_, _12671_);
  and _78183_ (_27028_, _27027_, _27025_);
  nor _78184_ (_27029_, _26886_, _12339_);
  or _78185_ (_27030_, _27029_, _27028_);
  nand _78186_ (_27031_, _27030_, _12336_);
  nor _78187_ (_27032_, _12248_, _12336_);
  nor _78188_ (_27033_, _27032_, _06042_);
  nand _78189_ (_27034_, _27033_, _27031_);
  and _78190_ (_27036_, _26886_, _06042_);
  nor _78191_ (_27037_, _27036_, _06339_);
  and _78192_ (_27038_, _27037_, _27034_);
  and _78193_ (_27039_, _12249_, _06339_);
  or _78194_ (_27040_, _27039_, _27038_);
  nand _78195_ (_27041_, _27040_, _07745_);
  and _78196_ (_27042_, _08953_, _06039_);
  nor _78197_ (_27043_, _27042_, _06486_);
  nand _78198_ (_27044_, _27043_, _27041_);
  and _78199_ (_27045_, _12427_, _06486_);
  nor _78200_ (_27047_, _27045_, _14022_);
  nand _78201_ (_27048_, _27047_, _27044_);
  nor _78202_ (_27049_, _12248_, _06334_);
  nor _78203_ (_27050_, _27049_, _06037_);
  nand _78204_ (_27051_, _27050_, _27048_);
  and _78205_ (_27052_, _12427_, _06037_);
  nor _78206_ (_27053_, _27052_, _12700_);
  nand _78207_ (_27054_, _27053_, _27051_);
  nor _78208_ (_27055_, _26886_, _12694_);
  nor _78209_ (_27056_, _27055_, _06401_);
  nand _78210_ (_27058_, _27056_, _27054_);
  and _78211_ (_27059_, _12248_, _06401_);
  nor _78212_ (_27060_, _27059_, _12696_);
  nand _78213_ (_27061_, _27060_, _27058_);
  and _78214_ (_27062_, _08953_, _12696_);
  nor _78215_ (_27063_, _27062_, _12704_);
  nand _78216_ (_27064_, _27063_, _27061_);
  nor _78217_ (_27065_, _26921_, _12705_);
  nor _78218_ (_27066_, _27065_, _08848_);
  and _78219_ (_27067_, _27066_, _27064_);
  nor _78220_ (_27069_, _12249_, _06277_);
  nor _78221_ (_27070_, _27069_, _08627_);
  or _78222_ (_27071_, _27070_, _27067_);
  and _78223_ (_27072_, _12427_, _06277_);
  nor _78224_ (_27073_, _27072_, _11028_);
  nand _78225_ (_27074_, _27073_, _27071_);
  and _78226_ (_27075_, _12249_, _11028_);
  nor _78227_ (_27076_, _27075_, _12718_);
  nand _78228_ (_27077_, _27076_, _27074_);
  and _78229_ (_27078_, _12743_, _12736_);
  not _78230_ (_27080_, _27078_);
  nor _78231_ (_27081_, _12744_, _12719_);
  and _78232_ (_27082_, _27081_, _27080_);
  nor _78233_ (_27083_, _27082_, _06400_);
  and _78234_ (_27084_, _27083_, _27077_);
  or _78235_ (_27085_, _27084_, _26893_);
  nand _78236_ (_27086_, _27085_, _06009_);
  and _78237_ (_27087_, _08953_, _06275_);
  nor _78238_ (_27088_, _27087_, _12763_);
  nand _78239_ (_27089_, _27088_, _27086_);
  and _78240_ (_27091_, _26921_, _12770_);
  and _78241_ (_27092_, _12249_, _11389_);
  nor _78242_ (_27093_, _27092_, _12764_);
  not _78243_ (_27094_, _27093_);
  nor _78244_ (_27095_, _27094_, _27091_);
  nor _78245_ (_27096_, _27095_, _12768_);
  and _78246_ (_27097_, _27096_, _27089_);
  or _78247_ (_27098_, _27097_, _26891_);
  nand _78248_ (_27099_, _27098_, _12330_);
  nor _78249_ (_27100_, _12248_, _12330_);
  nor _78250_ (_27102_, _27100_, _06502_);
  nand _78251_ (_27103_, _27102_, _27099_);
  and _78252_ (_27104_, _12427_, _06502_);
  nor _78253_ (_27105_, _27104_, _06615_);
  and _78254_ (_27106_, _27105_, _27103_);
  and _78255_ (_27107_, _12249_, _06615_);
  or _78256_ (_27108_, _27107_, _27106_);
  nand _78257_ (_27109_, _27108_, _06012_);
  and _78258_ (_27110_, _08953_, _12782_);
  nor _78259_ (_27111_, _27110_, _12787_);
  nand _78260_ (_27113_, _27111_, _27109_);
  and _78261_ (_27114_, _26921_, _11389_);
  nor _78262_ (_27115_, _12248_, _11389_);
  nor _78263_ (_27116_, _27115_, _12788_);
  not _78264_ (_27117_, _27116_);
  nor _78265_ (_27118_, _27117_, _27114_);
  nor _78266_ (_27119_, _27118_, _12792_);
  and _78267_ (_27120_, _27119_, _27113_);
  or _78268_ (_27121_, _27120_, _26890_);
  nand _78269_ (_27122_, _27121_, _12322_);
  nor _78270_ (_27124_, _12248_, _12322_);
  nor _78271_ (_27125_, _27124_, _06507_);
  nand _78272_ (_27126_, _27125_, _27122_);
  and _78273_ (_27127_, _12427_, _06507_);
  nor _78274_ (_27128_, _27127_, _06610_);
  and _78275_ (_27129_, _27128_, _27126_);
  and _78276_ (_27130_, _12249_, _06610_);
  or _78277_ (_27131_, _27130_, _27129_);
  nand _78278_ (_27132_, _27131_, _06018_);
  and _78279_ (_27133_, _08953_, _07330_);
  nor _78280_ (_27135_, _27133_, _12809_);
  nand _78281_ (_27136_, _27135_, _27132_);
  and _78282_ (_27137_, _12248_, \oc8051_golden_model_1.PSW [7]);
  nor _78283_ (_27138_, _26921_, \oc8051_golden_model_1.PSW [7]);
  or _78284_ (_27139_, _27138_, _27137_);
  and _78285_ (_27140_, _27139_, _12809_);
  nor _78286_ (_27141_, _27140_, _12814_);
  and _78287_ (_27142_, _27141_, _27136_);
  or _78288_ (_27143_, _27142_, _26889_);
  nand _78289_ (_27144_, _27143_, _12314_);
  nor _78290_ (_27145_, _12248_, _12314_);
  nor _78291_ (_27146_, _27145_, _06509_);
  nand _78292_ (_27147_, _27146_, _27144_);
  and _78293_ (_27148_, _12427_, _06509_);
  nor _78294_ (_27149_, _27148_, _06602_);
  and _78295_ (_27150_, _27149_, _27147_);
  and _78296_ (_27151_, _12249_, _06602_);
  or _78297_ (_27152_, _27151_, _27150_);
  nand _78298_ (_27153_, _27152_, _06023_);
  and _78299_ (_27154_, _08953_, _12827_);
  nor _78300_ (_27156_, _27154_, _12310_);
  nand _78301_ (_27157_, _27156_, _27153_);
  nand _78302_ (_27158_, _26921_, \oc8051_golden_model_1.PSW [7]);
  or _78303_ (_27159_, _12248_, \oc8051_golden_model_1.PSW [7]);
  and _78304_ (_27160_, _27159_, _12310_);
  and _78305_ (_27161_, _27160_, _27158_);
  nor _78306_ (_27162_, _27161_, _12839_);
  and _78307_ (_27163_, _27162_, _27157_);
  or _78308_ (_27164_, _27163_, _26888_);
  nand _78309_ (_27165_, _27164_, _11187_);
  nor _78310_ (_27167_, _12248_, _11187_);
  nor _78311_ (_27168_, _27167_, _11216_);
  nand _78312_ (_27169_, _27168_, _27165_);
  and _78313_ (_27170_, _26886_, _11216_);
  nor _78314_ (_27171_, _27170_, _06621_);
  and _78315_ (_27172_, _27171_, _27169_);
  nor _78316_ (_27173_, _09218_, _14116_);
  or _78317_ (_27174_, _27173_, _27172_);
  nand _78318_ (_27175_, _27174_, _06016_);
  and _78319_ (_27176_, _08953_, _07350_);
  nor _78320_ (_27177_, _27176_, _06512_);
  nand _78321_ (_27178_, _27177_, _27175_);
  and _78322_ (_27179_, _26900_, _13037_);
  nor _78323_ (_27180_, _12427_, _13037_);
  or _78324_ (_27181_, _27180_, _06629_);
  or _78325_ (_27182_, _27181_, _27179_);
  and _78326_ (_27183_, _27182_, _12201_);
  and _78327_ (_27184_, _27183_, _27178_);
  or _78328_ (_27185_, _27184_, _26887_);
  nand _78329_ (_27186_, _27185_, _13046_);
  nor _78330_ (_27187_, _13046_, _12248_);
  nor _78331_ (_27188_, _27187_, _10564_);
  nand _78332_ (_27189_, _27188_, _27186_);
  and _78333_ (_27190_, _26886_, _10564_);
  nor _78334_ (_27191_, _27190_, _06361_);
  and _78335_ (_27192_, _27191_, _27189_);
  nor _78336_ (_27193_, _09218_, _06362_);
  or _78337_ (_27194_, _27193_, _27192_);
  nand _78338_ (_27195_, _27194_, _06021_);
  and _78339_ (_27196_, _08953_, _12187_);
  nor _78340_ (_27197_, _27196_, _06496_);
  nand _78341_ (_27198_, _27197_, _27195_);
  and _78342_ (_27199_, _12428_, _13037_);
  nor _78343_ (_27200_, _26901_, _13037_);
  nor _78344_ (_27201_, _27200_, _27199_);
  and _78345_ (_27202_, _27201_, _06496_);
  nor _78346_ (_27203_, _27202_, _13062_);
  nand _78347_ (_27204_, _27203_, _27198_);
  nor _78348_ (_27205_, _26886_, _09123_);
  nor _78349_ (_27206_, _27205_, _06639_);
  nand _78350_ (_27207_, _27206_, _27204_);
  and _78351_ (_27208_, _12248_, _06639_);
  nor _78352_ (_27209_, _27208_, _26848_);
  and _78353_ (_27210_, _27209_, _27207_);
  nor _78354_ (_27211_, _26886_, _13072_);
  or _78355_ (_27212_, _27211_, _27210_);
  nand _78356_ (_27213_, _27212_, _07367_);
  and _78357_ (_27214_, _08953_, _07783_);
  nor _78358_ (_27215_, _27214_, _05989_);
  nand _78359_ (_27216_, _27215_, _27213_);
  and _78360_ (_27217_, _27201_, _05989_);
  nor _78361_ (_27218_, _27217_, _13088_);
  nand _78362_ (_27219_, _27218_, _27216_);
  nor _78363_ (_27220_, _26886_, _13087_);
  nor _78364_ (_27221_, _27220_, _06646_);
  and _78365_ (_27222_, _27221_, _27219_);
  or _78366_ (_27223_, _27222_, _26883_);
  nand _78367_ (_27224_, _27223_, _13095_);
  and _78368_ (_27225_, _26886_, _26866_);
  nor _78369_ (_27226_, _27225_, _25414_);
  nand _78370_ (_27228_, _27226_, _27224_);
  and _78371_ (_27229_, _25414_, _08953_);
  nor _78372_ (_27230_, _27229_, _13105_);
  and _78373_ (_27231_, _27230_, _27228_);
  and _78374_ (_27232_, _26886_, _13105_);
  or _78375_ (_27233_, _27232_, _27231_);
  or _78376_ (_27234_, _27233_, _01446_);
  or _78377_ (_27235_, _01442_, \oc8051_golden_model_1.PC [5]);
  and _78378_ (_27236_, _27235_, _43634_);
  and _78379_ (_44212_, _27236_, _27234_);
  and _78380_ (_27238_, _08918_, _07783_);
  and _78381_ (_27239_, _08607_, _12188_);
  nor _78382_ (_27240_, _27239_, \oc8051_golden_model_1.PC [6]);
  nor _78383_ (_27241_, _27240_, _12189_);
  not _78384_ (_27242_, _27241_);
  and _78385_ (_27243_, _27242_, _10564_);
  and _78386_ (_27244_, _12278_, _12245_);
  or _78387_ (_27245_, _27244_, _12279_);
  or _78388_ (_27246_, _27245_, _12705_);
  and _78389_ (_27247_, _27242_, _12347_);
  and _78390_ (_27248_, _12241_, _06352_);
  and _78391_ (_27249_, _27242_, _07269_);
  or _78392_ (_27250_, _27249_, _06474_);
  or _78393_ (_27251_, _27245_, _12539_);
  or _78394_ (_27252_, _12537_, _12241_);
  and _78395_ (_27253_, _27252_, _27251_);
  and _78396_ (_27254_, _27253_, _08687_);
  and _78397_ (_27255_, _08918_, _06816_);
  nor _78398_ (_27256_, _27241_, _12518_);
  nor _78399_ (_27257_, _26927_, \oc8051_golden_model_1.PC [6]);
  or _78400_ (_27259_, _27257_, _27256_);
  and _78401_ (_27260_, _27259_, _07260_);
  and _78402_ (_27261_, _12241_, _07259_);
  or _78403_ (_27262_, _27261_, _06855_);
  or _78404_ (_27263_, _27262_, _27260_);
  nand _78405_ (_27264_, _27241_, _06855_);
  and _78406_ (_27265_, _27264_, _07564_);
  and _78407_ (_27266_, _27265_, _27263_);
  or _78408_ (_27267_, _27266_, _25207_);
  or _78409_ (_27268_, _27267_, _27255_);
  or _78410_ (_27270_, _27242_, _12516_);
  and _78411_ (_27271_, _27270_, _08685_);
  and _78412_ (_27272_, _27271_, _27268_);
  or _78413_ (_27273_, _27272_, _27254_);
  and _78414_ (_27274_, _27273_, _07270_);
  or _78415_ (_27275_, _27274_, _27250_);
  and _78416_ (_27276_, _12464_, _12424_);
  nor _78417_ (_27277_, _27276_, _12465_);
  not _78418_ (_27278_, _27277_);
  or _78419_ (_27279_, _27278_, _12512_);
  or _78420_ (_27281_, _12510_, _12420_);
  and _78421_ (_27282_, _27281_, _27279_);
  or _78422_ (_27283_, _27282_, _07275_);
  and _78423_ (_27284_, _27283_, _27275_);
  or _78424_ (_27285_, _27284_, _25228_);
  or _78425_ (_27286_, _27242_, _12502_);
  and _78426_ (_27287_, _27286_, _06357_);
  and _78427_ (_27288_, _27287_, _27285_);
  and _78428_ (_27289_, _12241_, _06356_);
  or _78429_ (_27290_, _27289_, _07692_);
  or _78430_ (_27292_, _27290_, _27288_);
  or _78431_ (_27293_, _08918_, _06052_);
  and _78432_ (_27294_, _27293_, _06772_);
  and _78433_ (_27295_, _27294_, _27292_);
  nand _78434_ (_27296_, _12241_, _06410_);
  nand _78435_ (_27297_, _27296_, _12551_);
  or _78436_ (_27298_, _27297_, _27295_);
  or _78437_ (_27299_, _27242_, _12551_);
  and _78438_ (_27300_, _27299_, _06426_);
  and _78439_ (_27301_, _27300_, _27298_);
  nand _78440_ (_27302_, _12241_, _06417_);
  nand _78441_ (_27303_, _27302_, _12561_);
  or _78442_ (_27304_, _27303_, _27301_);
  or _78443_ (_27305_, _27242_, _12561_);
  and _78444_ (_27306_, _27305_, _06353_);
  and _78445_ (_27307_, _27306_, _27304_);
  or _78446_ (_27308_, _27307_, _27248_);
  and _78447_ (_27309_, _27308_, _06057_);
  and _78448_ (_27310_, _08918_, _12565_);
  or _78449_ (_27311_, _27310_, _06351_);
  or _78450_ (_27313_, _27311_, _27309_);
  nand _78451_ (_27314_, _12240_, _06351_);
  and _78452_ (_27315_, _27314_, _12574_);
  and _78453_ (_27316_, _27315_, _27313_);
  or _78454_ (_27317_, _27278_, _12609_);
  nand _78455_ (_27318_, _12609_, _12419_);
  and _78456_ (_27319_, _27318_, _12611_);
  and _78457_ (_27320_, _27319_, _27317_);
  or _78458_ (_27321_, _27320_, _27316_);
  and _78459_ (_27322_, _27321_, _06473_);
  or _78460_ (_27324_, _12420_, _12379_);
  nand _78461_ (_27325_, _27277_, _12379_);
  and _78462_ (_27326_, _27325_, _27324_);
  and _78463_ (_27327_, _27326_, _06472_);
  or _78464_ (_27328_, _27327_, _06431_);
  or _78465_ (_27329_, _27328_, _27322_);
  nand _78466_ (_27330_, _12630_, _12419_);
  or _78467_ (_27331_, _27278_, _12630_);
  and _78468_ (_27332_, _27331_, _27330_);
  or _78469_ (_27333_, _27332_, _06500_);
  and _78470_ (_27335_, _27333_, _27329_);
  or _78471_ (_27336_, _27335_, _06490_);
  nor _78472_ (_27337_, _27277_, _12648_);
  and _78473_ (_27338_, _12648_, _12420_);
  or _78474_ (_27339_, _27338_, _12349_);
  or _78475_ (_27340_, _27339_, _27337_);
  and _78476_ (_27341_, _27340_, _12348_);
  and _78477_ (_27342_, _27341_, _27336_);
  or _78478_ (_27343_, _27342_, _27247_);
  and _78479_ (_27344_, _27343_, _06346_);
  and _78480_ (_27346_, _12241_, _06345_);
  or _78481_ (_27347_, _27346_, _07596_);
  or _78482_ (_27348_, _27347_, _27344_);
  or _78483_ (_27349_, _08918_, _06049_);
  and _78484_ (_27350_, _27349_, _25555_);
  and _78485_ (_27351_, _27350_, _27348_);
  nor _78486_ (_27352_, _25555_, _12240_);
  or _78487_ (_27353_, _27352_, _27351_);
  and _78488_ (_27354_, _27353_, _12344_);
  nor _78489_ (_27355_, _27241_, _12344_);
  or _78490_ (_27357_, _27355_, _06445_);
  or _78491_ (_27358_, _27357_, _27354_);
  nand _78492_ (_27359_, _12240_, _06445_);
  and _78493_ (_27360_, _27359_, _06055_);
  and _78494_ (_27361_, _27360_, _27358_);
  and _78495_ (_27362_, _08918_, _25285_);
  or _78496_ (_27363_, _27362_, _06444_);
  or _78497_ (_27364_, _27363_, _27361_);
  nand _78498_ (_27365_, _12240_, _06444_);
  and _78499_ (_27366_, _27365_, _12339_);
  and _78500_ (_27367_, _27366_, _27364_);
  nor _78501_ (_27368_, _27241_, _12339_);
  or _78502_ (_27369_, _27368_, _12337_);
  or _78503_ (_27370_, _27369_, _27367_);
  or _78504_ (_27371_, _12241_, _12336_);
  and _78505_ (_27372_, _27371_, _06043_);
  and _78506_ (_27373_, _27372_, _27370_);
  and _78507_ (_27374_, _27242_, _06042_);
  or _78508_ (_27375_, _27374_, _27373_);
  and _78509_ (_27376_, _27375_, _06340_);
  and _78510_ (_27378_, _12241_, _06339_);
  or _78511_ (_27379_, _27378_, _06039_);
  or _78512_ (_27380_, _27379_, _27376_);
  or _78513_ (_27381_, _08918_, _07745_);
  and _78514_ (_27382_, _27381_, _06487_);
  and _78515_ (_27383_, _27382_, _27380_);
  nand _78516_ (_27384_, _12420_, _06486_);
  nand _78517_ (_27385_, _27384_, _06334_);
  or _78518_ (_27386_, _27385_, _27383_);
  or _78519_ (_27387_, _12241_, _06334_);
  and _78520_ (_27389_, _27387_, _06313_);
  and _78521_ (_27390_, _27389_, _27386_);
  nand _78522_ (_27391_, _12420_, _06037_);
  nand _78523_ (_27392_, _27391_, _12694_);
  or _78524_ (_27393_, _27392_, _27390_);
  or _78525_ (_27394_, _27242_, _12694_);
  and _78526_ (_27395_, _27394_, _25604_);
  and _78527_ (_27396_, _27395_, _27393_);
  and _78528_ (_27397_, _12241_, _06401_);
  or _78529_ (_27398_, _27397_, _12696_);
  or _78530_ (_27400_, _27398_, _27396_);
  or _78531_ (_27401_, _08918_, _06004_);
  and _78532_ (_27402_, _27401_, _27400_);
  or _78533_ (_27403_, _27402_, _12704_);
  and _78534_ (_27404_, _27403_, _27246_);
  or _78535_ (_27405_, _27404_, _08848_);
  or _78536_ (_27406_, _12241_, _08626_);
  and _78537_ (_27407_, _27406_, _06278_);
  and _78538_ (_27408_, _27407_, _27405_);
  and _78539_ (_27409_, _12420_, _06277_);
  or _78540_ (_27411_, _27409_, _11028_);
  or _78541_ (_27412_, _27411_, _27408_);
  nand _78542_ (_27413_, _12240_, _11028_);
  and _78543_ (_27414_, _27413_, _12719_);
  and _78544_ (_27415_, _27414_, _27412_);
  and _78545_ (_27416_, _12745_, _12732_);
  or _78546_ (_27417_, _27416_, _12746_);
  and _78547_ (_27418_, _27417_, _12718_);
  or _78548_ (_27419_, _27418_, _06400_);
  or _78549_ (_27420_, _27419_, _27415_);
  nand _78550_ (_27422_, _12240_, _06400_);
  and _78551_ (_27423_, _27422_, _06009_);
  and _78552_ (_27424_, _27423_, _27420_);
  and _78553_ (_27425_, _08918_, _06275_);
  or _78554_ (_27426_, _27425_, _12763_);
  or _78555_ (_27427_, _27426_, _27424_);
  and _78556_ (_27428_, _27245_, _12770_);
  nand _78557_ (_27429_, _12241_, _11389_);
  nand _78558_ (_27430_, _27429_, _12763_);
  or _78559_ (_27431_, _27430_, _27428_);
  and _78560_ (_27432_, _27431_, _12333_);
  and _78561_ (_27433_, _27432_, _27427_);
  nor _78562_ (_27434_, _27241_, _12333_);
  or _78563_ (_27435_, _27434_, _12331_);
  or _78564_ (_27436_, _27435_, _27433_);
  or _78565_ (_27437_, _12241_, _12330_);
  and _78566_ (_27438_, _27437_, _07334_);
  and _78567_ (_27439_, _27438_, _27436_);
  and _78568_ (_27440_, _12420_, _06502_);
  or _78569_ (_27441_, _27440_, _27439_);
  and _78570_ (_27443_, _27441_, _07337_);
  and _78571_ (_27444_, _12241_, _06615_);
  or _78572_ (_27445_, _27444_, _12782_);
  or _78573_ (_27446_, _27445_, _27443_);
  or _78574_ (_27447_, _08918_, _06012_);
  and _78575_ (_27448_, _27447_, _27446_);
  or _78576_ (_27449_, _27448_, _12787_);
  and _78577_ (_27450_, _27245_, _11389_);
  or _78578_ (_27451_, _12240_, _11389_);
  nand _78579_ (_27452_, _27451_, _12787_);
  or _78580_ (_27454_, _27452_, _27450_);
  and _78581_ (_27455_, _27454_, _12328_);
  and _78582_ (_27456_, _27455_, _27449_);
  nor _78583_ (_27457_, _27241_, _12328_);
  or _78584_ (_27458_, _27457_, _12323_);
  or _78585_ (_27459_, _27458_, _27456_);
  or _78586_ (_27460_, _12241_, _12322_);
  and _78587_ (_27461_, _27460_, _07339_);
  and _78588_ (_27462_, _27461_, _27459_);
  and _78589_ (_27463_, _12420_, _06507_);
  or _78590_ (_27465_, _27463_, _27462_);
  and _78591_ (_27466_, _27465_, _07331_);
  and _78592_ (_27467_, _12241_, _06610_);
  or _78593_ (_27468_, _27467_, _07330_);
  or _78594_ (_27469_, _27468_, _27466_);
  or _78595_ (_27470_, _08918_, _06018_);
  and _78596_ (_27471_, _27470_, _27469_);
  or _78597_ (_27472_, _27471_, _12809_);
  and _78598_ (_27473_, _27245_, _10967_);
  or _78599_ (_27474_, _12240_, _10967_);
  nand _78600_ (_27476_, _27474_, _12809_);
  or _78601_ (_27477_, _27476_, _27473_);
  and _78602_ (_27478_, _27477_, _12320_);
  and _78603_ (_27479_, _27478_, _27472_);
  nor _78604_ (_27480_, _27241_, _12320_);
  or _78605_ (_27481_, _27480_, _12315_);
  or _78606_ (_27482_, _27481_, _27479_);
  or _78607_ (_27483_, _12241_, _12314_);
  and _78608_ (_27484_, _27483_, _09107_);
  and _78609_ (_27485_, _27484_, _27482_);
  and _78610_ (_27487_, _12420_, _06509_);
  or _78611_ (_27488_, _27487_, _27485_);
  and _78612_ (_27489_, _27488_, _09112_);
  and _78613_ (_27490_, _12241_, _06602_);
  or _78614_ (_27491_, _27490_, _12827_);
  or _78615_ (_27492_, _27491_, _27489_);
  or _78616_ (_27493_, _08918_, _06023_);
  and _78617_ (_27494_, _27493_, _27492_);
  or _78618_ (_27495_, _27494_, _12310_);
  and _78619_ (_27496_, _27245_, \oc8051_golden_model_1.PSW [7]);
  or _78620_ (_27497_, _12240_, \oc8051_golden_model_1.PSW [7]);
  nand _78621_ (_27498_, _27497_, _12310_);
  or _78622_ (_27499_, _27498_, _27496_);
  and _78623_ (_27500_, _27499_, _12837_);
  and _78624_ (_27501_, _27500_, _27495_);
  nor _78625_ (_27502_, _27241_, _12837_);
  or _78626_ (_27503_, _27502_, _11188_);
  or _78627_ (_27504_, _27503_, _27501_);
  or _78628_ (_27505_, _12241_, _11187_);
  and _78629_ (_27506_, _27505_, _11217_);
  and _78630_ (_27508_, _27506_, _27504_);
  and _78631_ (_27509_, _27242_, _11216_);
  or _78632_ (_27510_, _27509_, _06621_);
  or _78633_ (_27511_, _27510_, _27508_);
  nand _78634_ (_27512_, _09172_, _06621_);
  and _78635_ (_27513_, _27512_, _06016_);
  and _78636_ (_27514_, _27513_, _27511_);
  and _78637_ (_27515_, _08918_, _07350_);
  or _78638_ (_27516_, _27515_, _06512_);
  or _78639_ (_27517_, _27516_, _27514_);
  and _78640_ (_27519_, _27278_, _13037_);
  nor _78641_ (_27520_, _12419_, _13037_);
  or _78642_ (_27521_, _27520_, _06629_);
  or _78643_ (_27522_, _27521_, _27519_);
  and _78644_ (_27523_, _27522_, _12201_);
  and _78645_ (_27524_, _27523_, _27517_);
  nor _78646_ (_27525_, _27241_, _12201_);
  or _78647_ (_27526_, _27525_, _13047_);
  or _78648_ (_27527_, _27526_, _27524_);
  or _78649_ (_27528_, _13046_, _12241_);
  and _78650_ (_27530_, _27528_, _13049_);
  and _78651_ (_27531_, _27530_, _27527_);
  or _78652_ (_27532_, _27531_, _27243_);
  and _78653_ (_27533_, _27532_, _06362_);
  nor _78654_ (_27534_, _09172_, _06362_);
  or _78655_ (_27535_, _27534_, _12187_);
  or _78656_ (_27536_, _27535_, _27533_);
  or _78657_ (_27537_, _08918_, _06021_);
  and _78658_ (_27538_, _27537_, _07035_);
  and _78659_ (_27539_, _27538_, _27536_);
  nor _78660_ (_27541_, _27277_, _13037_);
  and _78661_ (_27542_, _12420_, _13037_);
  or _78662_ (_27543_, _27542_, _27541_);
  and _78663_ (_27544_, _27543_, _06496_);
  or _78664_ (_27545_, _27544_, _27539_);
  and _78665_ (_27546_, _27545_, _09123_);
  nor _78666_ (_27547_, _27241_, _09123_);
  or _78667_ (_27548_, _27547_, _27546_);
  and _78668_ (_27549_, _27548_, _07048_);
  nand _78669_ (_27550_, _12241_, _06639_);
  nand _78670_ (_27552_, _27550_, _13072_);
  or _78671_ (_27553_, _27552_, _27549_);
  or _78672_ (_27554_, _27242_, _13072_);
  and _78673_ (_27555_, _27554_, _07367_);
  and _78674_ (_27556_, _27555_, _27553_);
  or _78675_ (_27557_, _27556_, _27238_);
  and _78676_ (_27558_, _27557_, _05990_);
  and _78677_ (_27559_, _27543_, _05989_);
  or _78678_ (_27560_, _27559_, _13088_);
  or _78679_ (_27561_, _27560_, _27558_);
  nor _78680_ (_27562_, _27242_, _13087_);
  nor _78681_ (_27563_, _27562_, _06646_);
  nand _78682_ (_27564_, _27563_, _27561_);
  and _78683_ (_27565_, _12241_, _06646_);
  nor _78684_ (_27566_, _27565_, _26866_);
  nand _78685_ (_27567_, _27566_, _27564_);
  nor _78686_ (_27568_, _27242_, _13095_);
  nor _78687_ (_27569_, _27568_, _25414_);
  and _78688_ (_27570_, _27569_, _27567_);
  and _78689_ (_27571_, _25414_, _08918_);
  or _78690_ (_27573_, _27571_, _13105_);
  nor _78691_ (_27574_, _27573_, _27570_);
  and _78692_ (_27575_, _27241_, _13105_);
  or _78693_ (_27576_, _27575_, _27574_);
  or _78694_ (_27577_, _27576_, _01446_);
  or _78695_ (_27578_, _01442_, \oc8051_golden_model_1.PC [6]);
  and _78696_ (_27579_, _27578_, _43634_);
  and _78697_ (_44213_, _27579_, _27577_);
  nor _78698_ (_27580_, _12189_, \oc8051_golden_model_1.PC [7]);
  nor _78699_ (_27581_, _27580_, _12190_);
  and _78700_ (_27583_, _27581_, _13105_);
  and _78701_ (_27584_, _08620_, _06646_);
  and _78702_ (_27585_, _08620_, _06639_);
  nor _78703_ (_27586_, _27581_, _12201_);
  nor _78704_ (_27587_, _27581_, _12837_);
  nor _78705_ (_27588_, _27581_, _12320_);
  nor _78706_ (_27589_, _27581_, _12328_);
  nor _78707_ (_27590_, _27581_, _12333_);
  nor _78708_ (_27591_, _25555_, _08620_);
  not _78709_ (_27592_, _27581_);
  and _78710_ (_27594_, _27592_, _12347_);
  nor _78711_ (_27595_, _08879_, _06052_);
  nor _78712_ (_27596_, _27581_, _12503_);
  or _78713_ (_27597_, _12510_, _08615_);
  or _78714_ (_27598_, _12415_, _12416_);
  and _78715_ (_27599_, _27598_, _12466_);
  nor _78716_ (_27600_, _27598_, _12466_);
  nor _78717_ (_27601_, _27600_, _27599_);
  not _78718_ (_27602_, _27601_);
  or _78719_ (_27603_, _27602_, _12512_);
  and _78720_ (_27605_, _27603_, _06474_);
  nand _78721_ (_27606_, _27605_, _27597_);
  or _78722_ (_27607_, _12236_, _12237_);
  and _78723_ (_27608_, _27607_, _12280_);
  nor _78724_ (_27609_, _27607_, _12280_);
  nor _78725_ (_27610_, _27609_, _27608_);
  nand _78726_ (_27611_, _27610_, _12537_);
  or _78727_ (_27612_, _12537_, _08814_);
  nand _78728_ (_27613_, _27612_, _27611_);
  nand _78729_ (_27614_, _27613_, _08687_);
  not _78730_ (_27616_, _12544_);
  nor _78731_ (_27617_, _26927_, \oc8051_golden_model_1.PC [7]);
  nor _78732_ (_27618_, _27617_, _07259_);
  and _78733_ (_27619_, _08620_, _07259_);
  nor _78734_ (_27620_, _27619_, _06855_);
  not _78735_ (_27621_, _27620_);
  nor _78736_ (_27622_, _27621_, _27618_);
  nor _78737_ (_27623_, _27581_, _12519_);
  nor _78738_ (_27624_, _27623_, _06816_);
  not _78739_ (_27625_, _27624_);
  nor _78740_ (_27627_, _27625_, _27622_);
  nor _78741_ (_27628_, _08879_, _07564_);
  or _78742_ (_27629_, _27628_, _25207_);
  nor _78743_ (_27630_, _27629_, _27627_);
  nor _78744_ (_27631_, _27581_, _12516_);
  or _78745_ (_27632_, _27631_, _08687_);
  nor _78746_ (_27633_, _27632_, _27630_);
  nor _78747_ (_27634_, _27633_, _27616_);
  nand _78748_ (_27635_, _27634_, _27614_);
  nand _78749_ (_27636_, _27635_, _27606_);
  and _78750_ (_27638_, _27636_, _12502_);
  or _78751_ (_27639_, _27638_, _27596_);
  nand _78752_ (_27640_, _27639_, _06357_);
  and _78753_ (_27641_, _08814_, _06356_);
  nor _78754_ (_27642_, _27641_, _07692_);
  and _78755_ (_27643_, _27642_, _27640_);
  or _78756_ (_27644_, _27643_, _27595_);
  nand _78757_ (_27645_, _27644_, _06772_);
  and _78758_ (_27646_, _08620_, _06410_);
  nor _78759_ (_27647_, _27646_, _12552_);
  nand _78760_ (_27648_, _27647_, _27645_);
  nor _78761_ (_27649_, _27581_, _12551_);
  nor _78762_ (_27650_, _27649_, _06417_);
  nand _78763_ (_27651_, _27650_, _27648_);
  and _78764_ (_27652_, _08620_, _06417_);
  nor _78765_ (_27653_, _27652_, _12563_);
  nand _78766_ (_27654_, _27653_, _27651_);
  nor _78767_ (_27655_, _27581_, _12561_);
  nor _78768_ (_27656_, _27655_, _06352_);
  nand _78769_ (_27657_, _27656_, _27654_);
  and _78770_ (_27659_, _08620_, _06352_);
  nor _78771_ (_27660_, _27659_, _12565_);
  nand _78772_ (_27661_, _27660_, _27657_);
  and _78773_ (_27662_, _08879_, _12565_);
  nor _78774_ (_27663_, _27662_, _06351_);
  nand _78775_ (_27664_, _27663_, _27661_);
  and _78776_ (_27665_, _08620_, _06351_);
  nor _78777_ (_27666_, _27665_, _12611_);
  and _78778_ (_27667_, _27666_, _27664_);
  and _78779_ (_27668_, _12609_, _08614_);
  nor _78780_ (_27670_, _27602_, _12609_);
  or _78781_ (_27671_, _27670_, _12574_);
  nor _78782_ (_27672_, _27671_, _27668_);
  nor _78783_ (_27673_, _27672_, _27667_);
  or _78784_ (_27674_, _27673_, _06472_);
  nand _78785_ (_27675_, _27601_, _12379_);
  or _78786_ (_27676_, _12379_, _08615_);
  and _78787_ (_27677_, _27676_, _06472_);
  nand _78788_ (_27678_, _27677_, _27675_);
  and _78789_ (_27679_, _27678_, _27674_);
  or _78790_ (_27681_, _27679_, _06431_);
  and _78791_ (_27682_, _12630_, _08614_);
  nor _78792_ (_27683_, _27602_, _12630_);
  or _78793_ (_27684_, _27683_, _06500_);
  or _78794_ (_27685_, _27684_, _27682_);
  and _78795_ (_27686_, _27685_, _12349_);
  nand _78796_ (_27687_, _27686_, _27681_);
  and _78797_ (_27688_, _12648_, _08614_);
  and _78798_ (_27689_, _27601_, _26636_);
  or _78799_ (_27690_, _27689_, _27688_);
  and _78800_ (_27692_, _27690_, _06490_);
  nor _78801_ (_27693_, _27692_, _12347_);
  and _78802_ (_27694_, _27693_, _27687_);
  or _78803_ (_27695_, _27694_, _27594_);
  nand _78804_ (_27696_, _27695_, _06346_);
  and _78805_ (_27697_, _08814_, _06345_);
  nor _78806_ (_27698_, _27697_, _07596_);
  nand _78807_ (_27699_, _27698_, _27696_);
  nor _78808_ (_27700_, _08879_, _06049_);
  nor _78809_ (_27701_, _27700_, _25556_);
  and _78810_ (_27703_, _27701_, _27699_);
  or _78811_ (_27704_, _27703_, _27591_);
  nand _78812_ (_27705_, _27704_, _12344_);
  nor _78813_ (_27706_, _27581_, _12344_);
  nor _78814_ (_27707_, _27706_, _06445_);
  nand _78815_ (_27708_, _27707_, _27705_);
  and _78816_ (_27709_, _08620_, _06445_);
  nor _78817_ (_27710_, _27709_, _25285_);
  nand _78818_ (_27711_, _27710_, _27708_);
  and _78819_ (_27712_, _08879_, _25285_);
  nor _78820_ (_27713_, _27712_, _06444_);
  nand _78821_ (_27714_, _27713_, _27711_);
  and _78822_ (_27715_, _08620_, _06444_);
  nor _78823_ (_27716_, _27715_, _12671_);
  and _78824_ (_27717_, _27716_, _27714_);
  nor _78825_ (_27718_, _27581_, _12339_);
  or _78826_ (_27719_, _27718_, _27717_);
  nand _78827_ (_27720_, _27719_, _12336_);
  nor _78828_ (_27721_, _12336_, _08620_);
  nor _78829_ (_27722_, _27721_, _06042_);
  nand _78830_ (_27724_, _27722_, _27720_);
  and _78831_ (_27725_, _27581_, _06042_);
  nor _78832_ (_27726_, _27725_, _06339_);
  and _78833_ (_27727_, _27726_, _27724_);
  and _78834_ (_27728_, _08814_, _06339_);
  or _78835_ (_27729_, _27728_, _27727_);
  nand _78836_ (_27730_, _27729_, _07745_);
  and _78837_ (_27731_, _08879_, _06039_);
  nor _78838_ (_27732_, _27731_, _06486_);
  nand _78839_ (_27733_, _27732_, _27730_);
  and _78840_ (_27735_, _08614_, _06486_);
  nor _78841_ (_27736_, _27735_, _14022_);
  nand _78842_ (_27737_, _27736_, _27733_);
  nor _78843_ (_27738_, _08620_, _06334_);
  nor _78844_ (_27739_, _27738_, _06037_);
  nand _78845_ (_27740_, _27739_, _27737_);
  and _78846_ (_27741_, _08614_, _06037_);
  nor _78847_ (_27742_, _27741_, _12700_);
  nand _78848_ (_27743_, _27742_, _27740_);
  nor _78849_ (_27744_, _27581_, _12694_);
  nor _78850_ (_27746_, _27744_, _06401_);
  nand _78851_ (_27747_, _27746_, _27743_);
  and _78852_ (_27748_, _08620_, _06401_);
  nor _78853_ (_27749_, _27748_, _12696_);
  nand _78854_ (_27750_, _27749_, _27747_);
  and _78855_ (_27751_, _08879_, _12696_);
  nor _78856_ (_27752_, _27751_, _12704_);
  nand _78857_ (_27753_, _27752_, _27750_);
  and _78858_ (_27754_, _27610_, _12704_);
  nor _78859_ (_27755_, _27754_, _08848_);
  and _78860_ (_27757_, _27755_, _27753_);
  nor _78861_ (_27758_, _08814_, _06277_);
  nor _78862_ (_27759_, _27758_, _08627_);
  or _78863_ (_27760_, _27759_, _27757_);
  and _78864_ (_27761_, _08614_, _06277_);
  nor _78865_ (_27762_, _27761_, _11028_);
  nand _78866_ (_27763_, _27762_, _27760_);
  and _78867_ (_27764_, _11028_, _08814_);
  nor _78868_ (_27765_, _27764_, _12718_);
  nand _78869_ (_27766_, _27765_, _27763_);
  or _78870_ (_27768_, _12728_, _12727_);
  nor _78871_ (_27769_, _27768_, _12747_);
  and _78872_ (_27770_, _27768_, _12747_);
  nor _78873_ (_27771_, _27770_, _27769_);
  and _78874_ (_27772_, _27771_, _12718_);
  nor _78875_ (_27773_, _27772_, _06400_);
  and _78876_ (_27774_, _27773_, _27766_);
  and _78877_ (_27775_, _08814_, _06400_);
  or _78878_ (_27776_, _27775_, _27774_);
  nand _78879_ (_27777_, _27776_, _06009_);
  and _78880_ (_27779_, _08879_, _06275_);
  nor _78881_ (_27780_, _27779_, _12763_);
  nand _78882_ (_27781_, _27780_, _27777_);
  nor _78883_ (_27782_, _27610_, _11389_);
  and _78884_ (_27783_, _11389_, _08814_);
  nor _78885_ (_27784_, _27783_, _12764_);
  not _78886_ (_27785_, _27784_);
  nor _78887_ (_27786_, _27785_, _27782_);
  nor _78888_ (_27787_, _27786_, _12768_);
  and _78889_ (_27788_, _27787_, _27781_);
  or _78890_ (_27790_, _27788_, _27590_);
  nand _78891_ (_27791_, _27790_, _12330_);
  nor _78892_ (_27792_, _12330_, _08620_);
  nor _78893_ (_27793_, _27792_, _06502_);
  nand _78894_ (_27794_, _27793_, _27791_);
  and _78895_ (_27795_, _08614_, _06502_);
  nor _78896_ (_27796_, _27795_, _06615_);
  and _78897_ (_27797_, _27796_, _27794_);
  and _78898_ (_27798_, _08814_, _06615_);
  or _78899_ (_27799_, _27798_, _27797_);
  nand _78900_ (_27801_, _27799_, _06012_);
  and _78901_ (_27802_, _08879_, _12782_);
  nor _78902_ (_27803_, _27802_, _12787_);
  nand _78903_ (_27804_, _27803_, _27801_);
  nor _78904_ (_27805_, _27610_, _12770_);
  nor _78905_ (_27806_, _11389_, _08620_);
  nor _78906_ (_27807_, _27806_, _12788_);
  not _78907_ (_27808_, _27807_);
  nor _78908_ (_27809_, _27808_, _27805_);
  nor _78909_ (_27810_, _27809_, _12792_);
  and _78910_ (_27812_, _27810_, _27804_);
  or _78911_ (_27813_, _27812_, _27589_);
  nand _78912_ (_27814_, _27813_, _12322_);
  nor _78913_ (_27815_, _12322_, _08620_);
  nor _78914_ (_27816_, _27815_, _06507_);
  nand _78915_ (_27817_, _27816_, _27814_);
  and _78916_ (_27818_, _08614_, _06507_);
  nor _78917_ (_27819_, _27818_, _06610_);
  and _78918_ (_27820_, _27819_, _27817_);
  and _78919_ (_27821_, _08814_, _06610_);
  or _78920_ (_27822_, _27821_, _27820_);
  nand _78921_ (_27823_, _27822_, _06018_);
  and _78922_ (_27824_, _08879_, _07330_);
  nor _78923_ (_27825_, _27824_, _12809_);
  nand _78924_ (_27826_, _27825_, _27823_);
  nor _78925_ (_27827_, _27610_, \oc8051_golden_model_1.PSW [7]);
  nor _78926_ (_27828_, _08620_, _10967_);
  nor _78927_ (_27829_, _27828_, _12810_);
  not _78928_ (_27830_, _27829_);
  nor _78929_ (_27831_, _27830_, _27827_);
  nor _78930_ (_27834_, _27831_, _12814_);
  and _78931_ (_27835_, _27834_, _27826_);
  or _78932_ (_27836_, _27835_, _27588_);
  nand _78933_ (_27837_, _27836_, _12314_);
  nor _78934_ (_27838_, _12314_, _08620_);
  nor _78935_ (_27839_, _27838_, _06509_);
  nand _78936_ (_27840_, _27839_, _27837_);
  and _78937_ (_27841_, _08614_, _06509_);
  nor _78938_ (_27842_, _27841_, _06602_);
  and _78939_ (_27843_, _27842_, _27840_);
  and _78940_ (_27845_, _08814_, _06602_);
  or _78941_ (_27846_, _27845_, _27843_);
  nand _78942_ (_27847_, _27846_, _06023_);
  and _78943_ (_27848_, _08879_, _12827_);
  nor _78944_ (_27849_, _27848_, _12310_);
  nand _78945_ (_27850_, _27849_, _27847_);
  and _78946_ (_27851_, _08620_, _10967_);
  and _78947_ (_27852_, _27610_, \oc8051_golden_model_1.PSW [7]);
  or _78948_ (_27853_, _27852_, _27851_);
  and _78949_ (_27854_, _27853_, _12310_);
  nor _78950_ (_27856_, _27854_, _12839_);
  and _78951_ (_27857_, _27856_, _27850_);
  or _78952_ (_27858_, _27857_, _27587_);
  nand _78953_ (_27859_, _27858_, _11187_);
  nor _78954_ (_27860_, _11187_, _08620_);
  nor _78955_ (_27861_, _27860_, _11216_);
  nand _78956_ (_27862_, _27861_, _27859_);
  and _78957_ (_27863_, _27581_, _11216_);
  nor _78958_ (_27864_, _27863_, _06621_);
  and _78959_ (_27865_, _27864_, _27862_);
  nor _78960_ (_27867_, _08778_, _14116_);
  or _78961_ (_27868_, _27867_, _27865_);
  nand _78962_ (_27869_, _27868_, _06016_);
  and _78963_ (_27870_, _08879_, _07350_);
  nor _78964_ (_27871_, _27870_, _06512_);
  nand _78965_ (_27872_, _27871_, _27869_);
  and _78966_ (_27873_, _27602_, _13037_);
  nor _78967_ (_27874_, _13037_, _08614_);
  or _78968_ (_27875_, _27874_, _06629_);
  or _78969_ (_27876_, _27875_, _27873_);
  and _78970_ (_27878_, _27876_, _12201_);
  and _78971_ (_27879_, _27878_, _27872_);
  or _78972_ (_27880_, _27879_, _27586_);
  nand _78973_ (_27881_, _27880_, _13046_);
  nor _78974_ (_27882_, _13046_, _08620_);
  nor _78975_ (_27883_, _27882_, _10564_);
  nand _78976_ (_27884_, _27883_, _27881_);
  and _78977_ (_27885_, _27581_, _10564_);
  nor _78978_ (_27886_, _27885_, _06361_);
  and _78979_ (_27887_, _27886_, _27884_);
  nor _78980_ (_27889_, _08778_, _06362_);
  or _78981_ (_27890_, _27889_, _27887_);
  nand _78982_ (_27891_, _27890_, _06021_);
  and _78983_ (_27892_, _08879_, _12187_);
  nor _78984_ (_27893_, _27892_, _06496_);
  nand _78985_ (_27894_, _27893_, _27891_);
  and _78986_ (_27895_, _13037_, _08615_);
  nor _78987_ (_27896_, _27601_, _13037_);
  nor _78988_ (_27897_, _27896_, _27895_);
  and _78989_ (_27898_, _27897_, _06496_);
  nor _78990_ (_27900_, _27898_, _13062_);
  nand _78991_ (_27901_, _27900_, _27894_);
  nor _78992_ (_27902_, _27581_, _09123_);
  nor _78993_ (_27903_, _27902_, _06639_);
  and _78994_ (_27904_, _27903_, _27901_);
  or _78995_ (_27905_, _27904_, _27585_);
  nand _78996_ (_27906_, _27905_, _13072_);
  nor _78997_ (_27907_, _27592_, _13072_);
  nor _78998_ (_27908_, _27907_, _07783_);
  nand _78999_ (_27909_, _27908_, _27906_);
  and _79000_ (_27911_, _08879_, _07783_);
  nor _79001_ (_27912_, _27911_, _05989_);
  nand _79002_ (_27913_, _27912_, _27909_);
  and _79003_ (_27914_, _27897_, _05989_);
  nor _79004_ (_27915_, _27914_, _13088_);
  nand _79005_ (_27916_, _27915_, _27913_);
  nor _79006_ (_27917_, _27581_, _13087_);
  nor _79007_ (_27918_, _27917_, _06646_);
  and _79008_ (_27919_, _27918_, _27916_);
  or _79009_ (_27920_, _27919_, _27584_);
  nand _79010_ (_27922_, _27920_, _13095_);
  nor _79011_ (_27923_, _27592_, _13095_);
  nor _79012_ (_27924_, _27923_, _25414_);
  nand _79013_ (_27925_, _27924_, _27922_);
  and _79014_ (_27926_, _25414_, _08879_);
  nor _79015_ (_27927_, _27926_, _13105_);
  and _79016_ (_27928_, _27927_, _27925_);
  or _79017_ (_27929_, _27928_, _27583_);
  or _79018_ (_27930_, _27929_, _01446_);
  or _79019_ (_27931_, _01442_, \oc8051_golden_model_1.PC [7]);
  and _79020_ (_27933_, _27931_, _43634_);
  and _79021_ (_44214_, _27933_, _27930_);
  nor _79022_ (_27934_, _13098_, _06310_);
  nor _79023_ (_27935_, _09534_, _06310_);
  nor _79024_ (_27936_, _12190_, \oc8051_golden_model_1.PC [8]);
  nor _79025_ (_27937_, _27936_, _12191_);
  nor _79026_ (_27938_, _27937_, _12201_);
  nor _79027_ (_27939_, _27937_, _12837_);
  nor _79028_ (_27940_, _27937_, _12320_);
  nor _79029_ (_27941_, _27937_, _12328_);
  and _79030_ (_27943_, _12412_, _06502_);
  nor _79031_ (_27944_, _27937_, _12333_);
  nor _79032_ (_27945_, _12704_, _12696_);
  nor _79033_ (_27946_, _25555_, _12234_);
  nor _79034_ (_27947_, _12470_, _12468_);
  nor _79035_ (_27948_, _27947_, _12471_);
  not _79036_ (_27949_, _27948_);
  and _79037_ (_27950_, _27949_, _12379_);
  nor _79038_ (_27951_, _12412_, _12379_);
  nor _79039_ (_27952_, _27951_, _27950_);
  nor _79040_ (_27954_, _27952_, _06473_);
  and _79041_ (_27955_, _12234_, _06352_);
  and _79042_ (_27956_, _12234_, _06410_);
  and _79043_ (_27957_, _12234_, _06356_);
  and _79044_ (_27958_, _27949_, _12510_);
  and _79045_ (_27959_, _12512_, _12413_);
  nor _79046_ (_27960_, _27959_, _27958_);
  or _79047_ (_27961_, _27960_, _07275_);
  and _79048_ (_27962_, _12539_, _12234_);
  nor _79049_ (_27963_, _12284_, _12282_);
  nor _79050_ (_27965_, _27963_, _12285_);
  and _79051_ (_27966_, _27965_, _12537_);
  or _79052_ (_27967_, _27966_, _27962_);
  nor _79053_ (_27968_, _27967_, _08685_);
  nand _79054_ (_27969_, _12234_, _07259_);
  not _79055_ (_27970_, \oc8051_golden_model_1.PC [8]);
  nor _79056_ (_27971_, _07259_, _27970_);
  nand _79057_ (_27972_, _27971_, _12518_);
  and _79058_ (_27973_, _27972_, _27969_);
  or _79059_ (_27974_, _27973_, _06855_);
  and _79060_ (_27976_, _27974_, _07564_);
  or _79061_ (_27977_, _27976_, _25207_);
  not _79062_ (_27978_, _27937_);
  or _79063_ (_27979_, _27978_, _12520_);
  and _79064_ (_27980_, _27979_, _08685_);
  and _79065_ (_27981_, _27980_, _27977_);
  or _79066_ (_27982_, _27981_, _07269_);
  nor _79067_ (_27983_, _27982_, _27968_);
  and _79068_ (_27984_, _27937_, _07269_);
  or _79069_ (_27985_, _27984_, _06474_);
  or _79070_ (_27987_, _27985_, _27983_);
  and _79071_ (_27988_, _27987_, _27961_);
  nor _79072_ (_27989_, _27988_, _25228_);
  nor _79073_ (_27990_, _27937_, _12502_);
  nor _79074_ (_27991_, _27990_, _06356_);
  not _79075_ (_27992_, _27991_);
  nor _79076_ (_27993_, _27992_, _27989_);
  nor _79077_ (_27994_, _27993_, _27957_);
  nor _79078_ (_27995_, _27994_, _07692_);
  and _79079_ (_27996_, _27995_, _06772_);
  or _79080_ (_27998_, _27996_, _12552_);
  or _79081_ (_27999_, _27998_, _27956_);
  nor _79082_ (_28000_, _27937_, _12551_);
  nor _79083_ (_28001_, _28000_, _06417_);
  nand _79084_ (_28002_, _28001_, _27999_);
  and _79085_ (_28003_, _12234_, _06417_);
  nor _79086_ (_28004_, _28003_, _12563_);
  nand _79087_ (_28005_, _28004_, _28002_);
  nor _79088_ (_28006_, _27937_, _12561_);
  nor _79089_ (_28007_, _28006_, _06352_);
  and _79090_ (_28009_, _28007_, _28005_);
  or _79091_ (_28010_, _28009_, _27955_);
  nand _79092_ (_28011_, _28010_, _12566_);
  and _79093_ (_28012_, _12234_, _06351_);
  nor _79094_ (_28013_, _28012_, _12611_);
  and _79095_ (_28014_, _28013_, _28011_);
  and _79096_ (_28015_, _12609_, _12412_);
  nor _79097_ (_28016_, _27949_, _12609_);
  or _79098_ (_28017_, _28016_, _28015_);
  nor _79099_ (_28018_, _28017_, _12574_);
  or _79100_ (_28020_, _28018_, _28014_);
  and _79101_ (_28021_, _28020_, _06473_);
  or _79102_ (_28022_, _28021_, _27954_);
  or _79103_ (_28023_, _28022_, _06431_);
  nor _79104_ (_28024_, _27949_, _12630_);
  and _79105_ (_28025_, _12630_, _12412_);
  nor _79106_ (_28026_, _28025_, _28024_);
  or _79107_ (_28027_, _28026_, _06500_);
  and _79108_ (_28028_, _28027_, _28023_);
  or _79109_ (_28029_, _28028_, _06490_);
  and _79110_ (_28031_, _12648_, _12412_);
  and _79111_ (_28032_, _27948_, _26636_);
  or _79112_ (_28033_, _28032_, _28031_);
  and _79113_ (_28034_, _28033_, _06490_);
  nor _79114_ (_28035_, _28034_, _12347_);
  nand _79115_ (_28036_, _28035_, _28029_);
  and _79116_ (_28037_, _27978_, _12347_);
  nor _79117_ (_28038_, _28037_, _06345_);
  nand _79118_ (_28039_, _28038_, _28036_);
  and _79119_ (_28040_, _12234_, _06345_);
  not _79120_ (_28042_, _28040_);
  and _79121_ (_28043_, _25555_, _06049_);
  and _79122_ (_28044_, _28043_, _28042_);
  and _79123_ (_28045_, _28044_, _28039_);
  or _79124_ (_28046_, _28045_, _27946_);
  nand _79125_ (_28047_, _28046_, _12344_);
  nor _79126_ (_28048_, _27937_, _12344_);
  nor _79127_ (_28049_, _28048_, _06445_);
  nand _79128_ (_28050_, _28049_, _28047_);
  and _79129_ (_28051_, _12234_, _06445_);
  nor _79130_ (_28053_, _28051_, _25285_);
  nand _79131_ (_28054_, _28053_, _28050_);
  nand _79132_ (_28055_, _28054_, _14251_);
  and _79133_ (_28056_, _12234_, _06444_);
  nor _79134_ (_28057_, _28056_, _12671_);
  and _79135_ (_28058_, _28057_, _28055_);
  nor _79136_ (_28059_, _27937_, _12339_);
  or _79137_ (_28060_, _28059_, _28058_);
  nand _79138_ (_28061_, _28060_, _12336_);
  nor _79139_ (_28062_, _12234_, _12336_);
  nor _79140_ (_28064_, _28062_, _06042_);
  nand _79141_ (_28065_, _28064_, _28061_);
  and _79142_ (_28066_, _27937_, _06042_);
  nor _79143_ (_28067_, _28066_, _06339_);
  nand _79144_ (_28068_, _28067_, _28065_);
  nor _79145_ (_28069_, _06486_, _06039_);
  not _79146_ (_28070_, _28069_);
  and _79147_ (_28071_, _14737_, _06339_);
  nor _79148_ (_28072_, _28071_, _28070_);
  nand _79149_ (_28073_, _28072_, _28068_);
  and _79150_ (_28075_, _12412_, _06486_);
  nor _79151_ (_28076_, _28075_, _14022_);
  nand _79152_ (_28077_, _28076_, _28073_);
  nor _79153_ (_28078_, _12234_, _06334_);
  nor _79154_ (_28079_, _28078_, _06037_);
  nand _79155_ (_28080_, _28079_, _28077_);
  and _79156_ (_28081_, _12412_, _06037_);
  nor _79157_ (_28082_, _28081_, _12700_);
  nand _79158_ (_28083_, _28082_, _28080_);
  nor _79159_ (_28084_, _27937_, _12694_);
  nor _79160_ (_28086_, _28084_, _06401_);
  and _79161_ (_28087_, _28086_, _28083_);
  and _79162_ (_28088_, _12234_, _06401_);
  or _79163_ (_28089_, _28088_, _28087_);
  nand _79164_ (_28090_, _28089_, _27945_);
  and _79165_ (_28091_, _27965_, _12704_);
  nor _79166_ (_28092_, _28091_, _08848_);
  nand _79167_ (_28093_, _28092_, _28090_);
  nor _79168_ (_28094_, _12234_, _08626_);
  nor _79169_ (_28095_, _28094_, _06277_);
  nand _79170_ (_28097_, _28095_, _28093_);
  and _79171_ (_28098_, _12412_, _06277_);
  nor _79172_ (_28099_, _28098_, _11028_);
  nand _79173_ (_28100_, _28099_, _28097_);
  and _79174_ (_28101_, _14737_, _11028_);
  nor _79175_ (_28102_, _28101_, _12718_);
  and _79176_ (_28103_, _28102_, _28100_);
  and _79177_ (_28104_, _12749_, _12726_);
  not _79178_ (_28105_, _28104_);
  nor _79179_ (_28106_, _12750_, _12719_);
  and _79180_ (_28108_, _28106_, _28105_);
  or _79181_ (_28109_, _28108_, _28103_);
  nand _79182_ (_28110_, _28109_, _06958_);
  and _79183_ (_28111_, _12234_, _06400_);
  nor _79184_ (_28112_, _28111_, _06275_);
  nand _79185_ (_28113_, _28112_, _28110_);
  nand _79186_ (_28114_, _28113_, _12764_);
  nor _79187_ (_28115_, _27965_, _11389_);
  and _79188_ (_28116_, _14737_, _11389_);
  nor _79189_ (_28117_, _28116_, _12764_);
  not _79190_ (_28119_, _28117_);
  nor _79191_ (_28120_, _28119_, _28115_);
  nor _79192_ (_28121_, _28120_, _12768_);
  and _79193_ (_28122_, _28121_, _28114_);
  or _79194_ (_28123_, _28122_, _27944_);
  nand _79195_ (_28124_, _28123_, _12330_);
  nor _79196_ (_28125_, _12234_, _12330_);
  nor _79197_ (_28126_, _28125_, _06502_);
  and _79198_ (_28127_, _28126_, _28124_);
  or _79199_ (_28128_, _28127_, _27943_);
  nand _79200_ (_28129_, _28128_, _07337_);
  and _79201_ (_28130_, _12234_, _06615_);
  nor _79202_ (_28131_, _28130_, _12782_);
  nand _79203_ (_28132_, _28131_, _28129_);
  nand _79204_ (_28133_, _28132_, _12788_);
  nor _79205_ (_28134_, _14737_, _11389_);
  and _79206_ (_28135_, _27965_, _11389_);
  or _79207_ (_28136_, _28135_, _28134_);
  and _79208_ (_28137_, _28136_, _12787_);
  nor _79209_ (_28138_, _28137_, _12792_);
  and _79210_ (_28141_, _28138_, _28133_);
  or _79211_ (_28142_, _28141_, _27941_);
  nand _79212_ (_28143_, _28142_, _12322_);
  nor _79213_ (_28144_, _12234_, _12322_);
  nor _79214_ (_28145_, _28144_, _06507_);
  nand _79215_ (_28146_, _28145_, _28143_);
  and _79216_ (_28147_, _12412_, _06507_);
  nor _79217_ (_28148_, _28147_, _06610_);
  nand _79218_ (_28149_, _28148_, _28146_);
  nor _79219_ (_28150_, _12809_, _07330_);
  and _79220_ (_28152_, _14737_, _06610_);
  not _79221_ (_28153_, _28152_);
  and _79222_ (_28154_, _28153_, _28150_);
  nand _79223_ (_28155_, _28154_, _28149_);
  and _79224_ (_28156_, _12234_, \oc8051_golden_model_1.PSW [7]);
  and _79225_ (_28157_, _27965_, _10967_);
  or _79226_ (_28158_, _28157_, _28156_);
  and _79227_ (_28159_, _28158_, _12809_);
  nor _79228_ (_28160_, _28159_, _12814_);
  and _79229_ (_28161_, _28160_, _28155_);
  or _79230_ (_28163_, _28161_, _27940_);
  nand _79231_ (_28164_, _28163_, _12314_);
  nor _79232_ (_28165_, _12234_, _12314_);
  nor _79233_ (_28166_, _28165_, _06509_);
  nand _79234_ (_28167_, _28166_, _28164_);
  and _79235_ (_28168_, _12412_, _06509_);
  nor _79236_ (_28169_, _28168_, _06602_);
  nand _79237_ (_28170_, _28169_, _28167_);
  nor _79238_ (_28171_, _12310_, _12827_);
  and _79239_ (_28172_, _14737_, _06602_);
  not _79240_ (_28174_, _28172_);
  and _79241_ (_28175_, _28174_, _28171_);
  nand _79242_ (_28176_, _28175_, _28170_);
  and _79243_ (_28177_, _12234_, _10967_);
  and _79244_ (_28178_, _27965_, \oc8051_golden_model_1.PSW [7]);
  or _79245_ (_28179_, _28178_, _28177_);
  and _79246_ (_28180_, _28179_, _12310_);
  nor _79247_ (_28181_, _28180_, _12839_);
  and _79248_ (_28182_, _28181_, _28176_);
  or _79249_ (_28183_, _28182_, _27939_);
  nand _79250_ (_28185_, _28183_, _11187_);
  nor _79251_ (_28186_, _12234_, _11187_);
  nor _79252_ (_28187_, _28186_, _11216_);
  and _79253_ (_28188_, _28187_, _28185_);
  and _79254_ (_28189_, _27937_, _11216_);
  or _79255_ (_28190_, _28189_, _28188_);
  nand _79256_ (_28191_, _28190_, _14116_);
  and _79257_ (_28192_, _07250_, _06621_);
  nor _79258_ (_28193_, _28192_, _07350_);
  nand _79259_ (_28194_, _28193_, _28191_);
  nand _79260_ (_28196_, _28194_, _06629_);
  nor _79261_ (_28197_, _12412_, _13037_);
  and _79262_ (_28198_, _27949_, _13037_);
  or _79263_ (_28199_, _28198_, _06629_);
  or _79264_ (_28200_, _28199_, _28197_);
  and _79265_ (_28201_, _28200_, _12201_);
  and _79266_ (_28202_, _28201_, _28196_);
  or _79267_ (_28203_, _28202_, _27938_);
  nand _79268_ (_28204_, _28203_, _13046_);
  nor _79269_ (_28205_, _13046_, _12234_);
  nor _79270_ (_28207_, _28205_, _10564_);
  and _79271_ (_28208_, _28207_, _28204_);
  and _79272_ (_28209_, _27937_, _10564_);
  or _79273_ (_28210_, _28209_, _28208_);
  nand _79274_ (_28211_, _28210_, _06362_);
  and _79275_ (_28212_, _07250_, _06361_);
  nor _79276_ (_28213_, _28212_, _12187_);
  nand _79277_ (_28214_, _28213_, _28211_);
  nand _79278_ (_28215_, _28214_, _07035_);
  and _79279_ (_28216_, _12413_, _13037_);
  nor _79280_ (_28218_, _27948_, _13037_);
  nor _79281_ (_28219_, _28218_, _28216_);
  and _79282_ (_28220_, _28219_, _06496_);
  nor _79283_ (_28221_, _28220_, _13062_);
  nand _79284_ (_28222_, _28221_, _28215_);
  nor _79285_ (_28223_, _27937_, _09123_);
  nor _79286_ (_28224_, _28223_, _06639_);
  nand _79287_ (_28225_, _28224_, _28222_);
  and _79288_ (_28226_, _12234_, _06639_);
  nor _79289_ (_28227_, _28226_, _26848_);
  nand _79290_ (_28229_, _28227_, _28225_);
  nor _79291_ (_28230_, _27937_, _13072_);
  nor _79292_ (_28231_, _28230_, _06503_);
  and _79293_ (_28232_, _28231_, _28229_);
  or _79294_ (_28233_, _28232_, _27935_);
  nor _79295_ (_28234_, _05998_, _05989_);
  nand _79296_ (_28235_, _28234_, _28233_);
  and _79297_ (_28236_, _28219_, _05989_);
  nor _79298_ (_28237_, _28236_, _13088_);
  nand _79299_ (_28238_, _28237_, _28235_);
  nor _79300_ (_28240_, _27937_, _13087_);
  nor _79301_ (_28241_, _28240_, _06646_);
  nand _79302_ (_28242_, _28241_, _28238_);
  and _79303_ (_28243_, _12234_, _06646_);
  nor _79304_ (_28244_, _28243_, _26866_);
  nand _79305_ (_28245_, _28244_, _28242_);
  nor _79306_ (_28246_, _27937_, _13095_);
  nor _79307_ (_28247_, _28246_, _06488_);
  and _79308_ (_28248_, _28247_, _28245_);
  or _79309_ (_28249_, _28248_, _27934_);
  nor _79310_ (_28251_, _13105_, _05997_);
  and _79311_ (_28252_, _28251_, _28249_);
  and _79312_ (_28253_, _27937_, _13105_);
  or _79313_ (_28254_, _28253_, _28252_);
  or _79314_ (_28255_, _28254_, _01446_);
  or _79315_ (_28256_, _01442_, \oc8051_golden_model_1.PC [8]);
  and _79316_ (_28257_, _28256_, _43634_);
  and _79317_ (_44215_, _28257_, _28255_);
  nor _79318_ (_28258_, _07127_, _13098_);
  nor _79319_ (_28259_, _07127_, _09534_);
  nor _79320_ (_28261_, _12191_, \oc8051_golden_model_1.PC [9]);
  nor _79321_ (_28262_, _28261_, _12192_);
  nor _79322_ (_28263_, _28262_, _12201_);
  nor _79323_ (_28264_, _28262_, _12837_);
  and _79324_ (_28265_, _12407_, _06509_);
  nor _79325_ (_28266_, _28262_, _12320_);
  and _79326_ (_28267_, _12407_, _06507_);
  nor _79327_ (_28268_, _28262_, _12328_);
  and _79328_ (_28269_, _12407_, _06502_);
  nor _79329_ (_28270_, _28262_, _12333_);
  and _79330_ (_28272_, _12230_, _06444_);
  nor _79331_ (_28273_, _06444_, _25285_);
  not _79332_ (_28274_, _28262_);
  and _79333_ (_28275_, _28274_, _12347_);
  nand _79334_ (_28276_, _12230_, _07259_);
  not _79335_ (_28277_, \oc8051_golden_model_1.PC [9]);
  nor _79336_ (_28278_, _07259_, _28277_);
  nand _79337_ (_28279_, _28278_, _12518_);
  and _79338_ (_28280_, _28279_, _28276_);
  or _79339_ (_28281_, _28280_, _06855_);
  and _79340_ (_28283_, _28281_, _07564_);
  or _79341_ (_28284_, _28283_, _25207_);
  or _79342_ (_28285_, _28274_, _12520_);
  and _79343_ (_28286_, _28285_, _08685_);
  and _79344_ (_28287_, _28286_, _28284_);
  and _79345_ (_28288_, _12539_, _12230_);
  or _79346_ (_28289_, _12232_, _12231_);
  not _79347_ (_28290_, _28289_);
  nor _79348_ (_28291_, _28290_, _12286_);
  and _79349_ (_28292_, _28290_, _12286_);
  nor _79350_ (_28294_, _28292_, _28291_);
  nor _79351_ (_28295_, _28294_, _12539_);
  or _79352_ (_28296_, _28295_, _28288_);
  nor _79353_ (_28297_, _28296_, _08685_);
  nor _79354_ (_28298_, _28297_, _28287_);
  nor _79355_ (_28299_, _28298_, _07269_);
  and _79356_ (_28300_, _28274_, _07269_);
  nor _79357_ (_28301_, _28300_, _28299_);
  and _79358_ (_28302_, _28301_, _07275_);
  and _79359_ (_28303_, _12512_, _12408_);
  or _79360_ (_28305_, _12410_, _12409_);
  not _79361_ (_28306_, _28305_);
  nor _79362_ (_28307_, _28306_, _12472_);
  and _79363_ (_28308_, _28306_, _12472_);
  nor _79364_ (_28309_, _28308_, _28307_);
  and _79365_ (_28310_, _28309_, _12510_);
  nor _79366_ (_28311_, _28310_, _28303_);
  and _79367_ (_28312_, _28311_, _06474_);
  or _79368_ (_28313_, _28312_, _28302_);
  nor _79369_ (_28314_, _28313_, _25228_);
  nor _79370_ (_28316_, _28262_, _12502_);
  nor _79371_ (_28317_, _28316_, _06356_);
  not _79372_ (_28318_, _28317_);
  or _79373_ (_28319_, _28318_, _28314_);
  and _79374_ (_28320_, _12230_, _06356_);
  nor _79375_ (_28321_, _28320_, _07692_);
  nand _79376_ (_28322_, _28321_, _28319_);
  nand _79377_ (_28323_, _28322_, _06772_);
  and _79378_ (_28324_, _12230_, _06410_);
  nor _79379_ (_28325_, _28324_, _12552_);
  nand _79380_ (_28327_, _28325_, _28323_);
  nor _79381_ (_28328_, _28262_, _12551_);
  nor _79382_ (_28329_, _28328_, _06417_);
  nand _79383_ (_28330_, _28329_, _28327_);
  and _79384_ (_28331_, _12230_, _06417_);
  nor _79385_ (_28332_, _28331_, _12563_);
  nand _79386_ (_28333_, _28332_, _28330_);
  nor _79387_ (_28334_, _28262_, _12561_);
  nor _79388_ (_28335_, _28334_, _06352_);
  nand _79389_ (_28336_, _28335_, _28333_);
  and _79390_ (_28338_, _12230_, _06352_);
  nor _79391_ (_28339_, _28338_, _12565_);
  nand _79392_ (_28340_, _28339_, _28336_);
  nand _79393_ (_28341_, _28340_, _07394_);
  and _79394_ (_28342_, _12230_, _06351_);
  nor _79395_ (_28343_, _28342_, _12611_);
  and _79396_ (_28344_, _28343_, _28341_);
  and _79397_ (_28345_, _12609_, _12407_);
  nor _79398_ (_28346_, _28309_, _12609_);
  or _79399_ (_28347_, _28346_, _28345_);
  nor _79400_ (_28349_, _28347_, _12574_);
  or _79401_ (_28350_, _28349_, _28344_);
  nand _79402_ (_28351_, _28350_, _06473_);
  nor _79403_ (_28352_, _12408_, _12379_);
  not _79404_ (_28353_, _28309_);
  and _79405_ (_28354_, _28353_, _12379_);
  or _79406_ (_28355_, _28354_, _28352_);
  nor _79407_ (_28356_, _28355_, _06473_);
  nor _79408_ (_28357_, _28356_, _06431_);
  nand _79409_ (_28358_, _28357_, _28351_);
  and _79410_ (_28360_, _12630_, _12408_);
  nor _79411_ (_28361_, _28353_, _12630_);
  or _79412_ (_28362_, _28361_, _06500_);
  or _79413_ (_28363_, _28362_, _28360_);
  nand _79414_ (_28364_, _28363_, _28358_);
  nand _79415_ (_28365_, _28364_, _12349_);
  and _79416_ (_28366_, _12648_, _12407_);
  nor _79417_ (_28367_, _28309_, _12648_);
  or _79418_ (_28368_, _28367_, _28366_);
  and _79419_ (_28369_, _28368_, _06490_);
  nor _79420_ (_28371_, _28369_, _12347_);
  and _79421_ (_28372_, _28371_, _28365_);
  or _79422_ (_28373_, _28372_, _28275_);
  nand _79423_ (_28374_, _28373_, _06346_);
  and _79424_ (_28375_, _14934_, _06345_);
  not _79425_ (_28376_, _28375_);
  and _79426_ (_28377_, _28376_, _28043_);
  nand _79427_ (_28378_, _28377_, _28374_);
  nor _79428_ (_28379_, _25555_, _14934_);
  nor _79429_ (_28380_, _28379_, _12345_);
  nand _79430_ (_28382_, _28380_, _28378_);
  nor _79431_ (_28383_, _28262_, _12344_);
  nor _79432_ (_28384_, _28383_, _06445_);
  and _79433_ (_28385_, _28384_, _28382_);
  and _79434_ (_28386_, _12230_, _06445_);
  or _79435_ (_28387_, _28386_, _28385_);
  and _79436_ (_28388_, _28387_, _28273_);
  or _79437_ (_28389_, _28388_, _28272_);
  nand _79438_ (_28390_, _28389_, _12339_);
  nor _79439_ (_28391_, _28274_, _12339_);
  nor _79440_ (_28393_, _28391_, _12337_);
  nand _79441_ (_28394_, _28393_, _28390_);
  nor _79442_ (_28395_, _12230_, _12336_);
  nor _79443_ (_28396_, _28395_, _06042_);
  nand _79444_ (_28397_, _28396_, _28394_);
  and _79445_ (_28398_, _28262_, _06042_);
  nor _79446_ (_28399_, _28398_, _06339_);
  nand _79447_ (_28400_, _28399_, _28397_);
  and _79448_ (_28401_, _14934_, _06339_);
  nor _79449_ (_28402_, _28401_, _28070_);
  nand _79450_ (_28404_, _28402_, _28400_);
  and _79451_ (_28405_, _12407_, _06486_);
  nor _79452_ (_28406_, _28405_, _14022_);
  nand _79453_ (_28407_, _28406_, _28404_);
  nor _79454_ (_28408_, _12230_, _06334_);
  nor _79455_ (_28409_, _28408_, _06037_);
  nand _79456_ (_28410_, _28409_, _28407_);
  and _79457_ (_28411_, _12407_, _06037_);
  nor _79458_ (_28412_, _28411_, _12700_);
  nand _79459_ (_28413_, _28412_, _28410_);
  nor _79460_ (_28415_, _28262_, _12694_);
  nor _79461_ (_28416_, _28415_, _06401_);
  and _79462_ (_28417_, _28416_, _28413_);
  and _79463_ (_28418_, _12230_, _06401_);
  or _79464_ (_28419_, _28418_, _28417_);
  nand _79465_ (_28420_, _28419_, _27945_);
  nor _79466_ (_28421_, _28294_, _12705_);
  nor _79467_ (_28422_, _28421_, _08848_);
  and _79468_ (_28423_, _28422_, _28420_);
  nor _79469_ (_28424_, _14934_, _06277_);
  nor _79470_ (_28426_, _28424_, _08627_);
  or _79471_ (_28427_, _28426_, _28423_);
  and _79472_ (_28428_, _12407_, _06277_);
  nor _79473_ (_28429_, _28428_, _11028_);
  nand _79474_ (_28430_, _28429_, _28427_);
  and _79475_ (_28431_, _14934_, _11028_);
  nor _79476_ (_28432_, _28431_, _12718_);
  and _79477_ (_28433_, _28432_, _28430_);
  nor _79478_ (_28434_, _12750_, \oc8051_golden_model_1.DPH [1]);
  not _79479_ (_28435_, _28434_);
  nor _79480_ (_28437_, _12751_, _12719_);
  and _79481_ (_28438_, _28437_, _28435_);
  or _79482_ (_28439_, _28438_, _28433_);
  nand _79483_ (_28440_, _28439_, _06958_);
  and _79484_ (_28441_, _12230_, _06400_);
  nor _79485_ (_28442_, _28441_, _06275_);
  nand _79486_ (_28443_, _28442_, _28440_);
  nand _79487_ (_28444_, _28443_, _12764_);
  and _79488_ (_28445_, _28294_, _12770_);
  and _79489_ (_28446_, _14934_, _11389_);
  nor _79490_ (_28448_, _28446_, _12764_);
  not _79491_ (_28449_, _28448_);
  nor _79492_ (_28450_, _28449_, _28445_);
  nor _79493_ (_28451_, _28450_, _12768_);
  and _79494_ (_28452_, _28451_, _28444_);
  or _79495_ (_28453_, _28452_, _28270_);
  nand _79496_ (_28454_, _28453_, _12330_);
  nor _79497_ (_28455_, _12230_, _12330_);
  nor _79498_ (_28456_, _28455_, _06502_);
  and _79499_ (_28457_, _28456_, _28454_);
  or _79500_ (_28459_, _28457_, _28269_);
  nand _79501_ (_28460_, _28459_, _07337_);
  and _79502_ (_28461_, _12230_, _06615_);
  nor _79503_ (_28462_, _28461_, _12782_);
  nand _79504_ (_28463_, _28462_, _28460_);
  nand _79505_ (_28464_, _28463_, _12788_);
  and _79506_ (_28465_, _12230_, _12770_);
  nor _79507_ (_28466_, _28294_, _12770_);
  or _79508_ (_28467_, _28466_, _28465_);
  and _79509_ (_28468_, _28467_, _12787_);
  nor _79510_ (_28470_, _28468_, _12792_);
  and _79511_ (_28471_, _28470_, _28464_);
  or _79512_ (_28472_, _28471_, _28268_);
  nand _79513_ (_28473_, _28472_, _12322_);
  nor _79514_ (_28474_, _12230_, _12322_);
  nor _79515_ (_28475_, _28474_, _06507_);
  and _79516_ (_28476_, _28475_, _28473_);
  or _79517_ (_28477_, _28476_, _28267_);
  nand _79518_ (_28478_, _28477_, _07331_);
  and _79519_ (_28479_, _12230_, _06610_);
  nor _79520_ (_28480_, _28479_, _07330_);
  nand _79521_ (_28481_, _28480_, _28478_);
  nand _79522_ (_28482_, _28481_, _12810_);
  and _79523_ (_28483_, _28294_, _10967_);
  nor _79524_ (_28484_, _12230_, _10967_);
  nor _79525_ (_28485_, _28484_, _12810_);
  not _79526_ (_28486_, _28485_);
  nor _79527_ (_28487_, _28486_, _28483_);
  nor _79528_ (_28488_, _28487_, _12814_);
  and _79529_ (_28489_, _28488_, _28482_);
  or _79530_ (_28492_, _28489_, _28266_);
  nand _79531_ (_28493_, _28492_, _12314_);
  nor _79532_ (_28494_, _12230_, _12314_);
  nor _79533_ (_28495_, _28494_, _06509_);
  and _79534_ (_28496_, _28495_, _28493_);
  or _79535_ (_28497_, _28496_, _28265_);
  nand _79536_ (_28498_, _28497_, _09112_);
  and _79537_ (_28499_, _12230_, _06602_);
  nor _79538_ (_28500_, _28499_, _12827_);
  nand _79539_ (_28501_, _28500_, _28498_);
  nand _79540_ (_28503_, _28501_, _12832_);
  and _79541_ (_28504_, _12230_, _10967_);
  nor _79542_ (_28505_, _28294_, _10967_);
  or _79543_ (_28506_, _28505_, _28504_);
  and _79544_ (_28507_, _28506_, _12310_);
  nor _79545_ (_28508_, _28507_, _12839_);
  and _79546_ (_28509_, _28508_, _28503_);
  or _79547_ (_28510_, _28509_, _28264_);
  nand _79548_ (_28511_, _28510_, _11187_);
  nor _79549_ (_28512_, _12230_, _11187_);
  nor _79550_ (_28514_, _28512_, _11216_);
  nand _79551_ (_28515_, _28514_, _28511_);
  and _79552_ (_28516_, _28262_, _11216_);
  nor _79553_ (_28517_, _28516_, _06621_);
  nand _79554_ (_28518_, _28517_, _28515_);
  nor _79555_ (_28519_, _06512_, _07350_);
  not _79556_ (_28520_, _28519_);
  and _79557_ (_28521_, _07448_, _06621_);
  nor _79558_ (_28522_, _28521_, _28520_);
  nand _79559_ (_28523_, _28522_, _28518_);
  and _79560_ (_28525_, _28309_, _13037_);
  nor _79561_ (_28526_, _12407_, _13037_);
  or _79562_ (_28527_, _28526_, _06629_);
  or _79563_ (_28528_, _28527_, _28525_);
  and _79564_ (_28529_, _28528_, _12201_);
  and _79565_ (_28530_, _28529_, _28523_);
  or _79566_ (_28531_, _28530_, _28263_);
  nand _79567_ (_28532_, _28531_, _13046_);
  nor _79568_ (_28533_, _13046_, _12230_);
  nor _79569_ (_28534_, _28533_, _10564_);
  nand _79570_ (_28536_, _28534_, _28532_);
  and _79571_ (_28537_, _28262_, _10564_);
  nor _79572_ (_28538_, _28537_, _06361_);
  nand _79573_ (_28539_, _28538_, _28536_);
  nor _79574_ (_28540_, _06496_, _12187_);
  not _79575_ (_28541_, _28540_);
  and _79576_ (_28542_, _07448_, _06361_);
  nor _79577_ (_28543_, _28542_, _28541_);
  nand _79578_ (_28544_, _28543_, _28539_);
  and _79579_ (_28545_, _12408_, _13037_);
  nor _79580_ (_28547_, _28353_, _13037_);
  nor _79581_ (_28548_, _28547_, _28545_);
  and _79582_ (_28549_, _28548_, _06496_);
  nor _79583_ (_28550_, _28549_, _13062_);
  nand _79584_ (_28551_, _28550_, _28544_);
  nor _79585_ (_28552_, _28262_, _09123_);
  nor _79586_ (_28553_, _28552_, _06639_);
  nand _79587_ (_28554_, _28553_, _28551_);
  and _79588_ (_28555_, _12230_, _06639_);
  nor _79589_ (_28556_, _28555_, _26848_);
  nand _79590_ (_28558_, _28556_, _28554_);
  nor _79591_ (_28559_, _28262_, _13072_);
  nor _79592_ (_28560_, _28559_, _06503_);
  and _79593_ (_28561_, _28560_, _28558_);
  or _79594_ (_28562_, _28561_, _28259_);
  nand _79595_ (_28563_, _28562_, _28234_);
  and _79596_ (_28564_, _28548_, _05989_);
  nor _79597_ (_28565_, _28564_, _13088_);
  nand _79598_ (_28566_, _28565_, _28563_);
  nor _79599_ (_28567_, _28262_, _13087_);
  nor _79600_ (_28569_, _28567_, _06646_);
  nand _79601_ (_28570_, _28569_, _28566_);
  and _79602_ (_28571_, _12230_, _06646_);
  nor _79603_ (_28572_, _28571_, _26866_);
  nand _79604_ (_28573_, _28572_, _28570_);
  nor _79605_ (_28574_, _28262_, _13095_);
  nor _79606_ (_28575_, _28574_, _06488_);
  and _79607_ (_28576_, _28575_, _28573_);
  or _79608_ (_28577_, _28576_, _28258_);
  and _79609_ (_28578_, _28577_, _28251_);
  and _79610_ (_28580_, _28262_, _13105_);
  or _79611_ (_28581_, _28580_, _28578_);
  or _79612_ (_28582_, _28581_, _01446_);
  or _79613_ (_28583_, _01442_, \oc8051_golden_model_1.PC [9]);
  and _79614_ (_28584_, _28583_, _43634_);
  and _79615_ (_44216_, _28584_, _28582_);
  nand _79616_ (_28585_, _12401_, _06507_);
  nor _79617_ (_28586_, _12192_, \oc8051_golden_model_1.PC [10]);
  nor _79618_ (_28587_, _28586_, _12193_);
  not _79619_ (_28588_, _28587_);
  nor _79620_ (_28590_, _28588_, _12694_);
  or _79621_ (_28591_, _28587_, _12551_);
  nor _79622_ (_28592_, _12475_, _12404_);
  nor _79623_ (_28593_, _28592_, _12476_);
  or _79624_ (_28594_, _28593_, _12512_);
  or _79625_ (_28595_, _12510_, _12400_);
  and _79626_ (_28596_, _28595_, _28594_);
  or _79627_ (_28597_, _28596_, _07275_);
  and _79628_ (_28598_, _12539_, _12224_);
  nor _79629_ (_28599_, _12289_, _12227_);
  nor _79630_ (_28601_, _28599_, _12290_);
  and _79631_ (_28602_, _28601_, _12537_);
  or _79632_ (_28603_, _28602_, _28598_);
  or _79633_ (_28604_, _28603_, _08685_);
  and _79634_ (_28605_, _12224_, _07259_);
  and _79635_ (_28606_, _07260_, \oc8051_golden_model_1.PC [10]);
  and _79636_ (_28607_, _28606_, _12518_);
  or _79637_ (_28608_, _28607_, _28605_);
  and _79638_ (_28609_, _28608_, _12517_);
  or _79639_ (_28610_, _28609_, _06816_);
  and _79640_ (_28612_, _28610_, _12516_);
  nor _79641_ (_28613_, _28588_, _12520_);
  or _79642_ (_28614_, _28613_, _08687_);
  or _79643_ (_28615_, _28614_, _28612_);
  and _79644_ (_28616_, _28615_, _07270_);
  and _79645_ (_28617_, _28616_, _28604_);
  and _79646_ (_28618_, _28587_, _07269_);
  or _79647_ (_28619_, _28618_, _06474_);
  or _79648_ (_28620_, _28619_, _28617_);
  and _79649_ (_28621_, _28620_, _28597_);
  or _79650_ (_28623_, _28621_, _25228_);
  or _79651_ (_28624_, _28587_, _12502_);
  and _79652_ (_28625_, _28624_, _06357_);
  and _79653_ (_28626_, _28625_, _28623_);
  or _79654_ (_28627_, _28626_, _07692_);
  and _79655_ (_28628_, _28627_, _06772_);
  and _79656_ (_28629_, _12224_, _14297_);
  or _79657_ (_28630_, _28629_, _12552_);
  or _79658_ (_28631_, _28630_, _28628_);
  and _79659_ (_28632_, _28631_, _28591_);
  or _79660_ (_28634_, _28632_, _06417_);
  or _79661_ (_28635_, _12224_, _06426_);
  and _79662_ (_28636_, _28635_, _12561_);
  and _79663_ (_28637_, _28636_, _28634_);
  nor _79664_ (_28638_, _28588_, _12561_);
  or _79665_ (_28639_, _28638_, _28637_);
  and _79666_ (_28640_, _28639_, _06353_);
  and _79667_ (_28641_, _12224_, _06352_);
  or _79668_ (_28642_, _28641_, _12565_);
  or _79669_ (_28643_, _28642_, _28640_);
  and _79670_ (_28645_, _28643_, _07394_);
  nand _79671_ (_28646_, _12224_, _06351_);
  nand _79672_ (_28647_, _28646_, _12574_);
  or _79673_ (_28648_, _28647_, _28645_);
  or _79674_ (_28649_, _28593_, _12609_);
  nand _79675_ (_28650_, _12609_, _12401_);
  and _79676_ (_28651_, _28650_, _28649_);
  or _79677_ (_28652_, _28651_, _12574_);
  and _79678_ (_28653_, _28652_, _28648_);
  or _79679_ (_28654_, _28653_, _06472_);
  and _79680_ (_28656_, _28593_, _12379_);
  nor _79681_ (_28657_, _12401_, _12379_);
  or _79682_ (_28658_, _28657_, _28656_);
  or _79683_ (_28659_, _28658_, _06473_);
  and _79684_ (_28660_, _28659_, _06500_);
  and _79685_ (_28661_, _28660_, _28654_);
  and _79686_ (_28662_, _12630_, _12400_);
  and _79687_ (_28663_, _28593_, _12632_);
  or _79688_ (_28664_, _28663_, _28662_);
  and _79689_ (_28665_, _28664_, _06431_);
  or _79690_ (_28667_, _28665_, _28661_);
  and _79691_ (_28668_, _28667_, _12349_);
  or _79692_ (_28669_, _28593_, _12648_);
  nand _79693_ (_28670_, _12648_, _12401_);
  and _79694_ (_28671_, _28670_, _06490_);
  and _79695_ (_28672_, _28671_, _28669_);
  or _79696_ (_28673_, _28672_, _12347_);
  or _79697_ (_28674_, _28673_, _28668_);
  nand _79698_ (_28675_, _28588_, _12347_);
  and _79699_ (_28676_, _28675_, _06346_);
  and _79700_ (_28678_, _28676_, _28674_);
  or _79701_ (_28679_, _28678_, _07596_);
  and _79702_ (_28680_, _28679_, _25555_);
  nand _79703_ (_28681_, _25555_, _06346_);
  and _79704_ (_28682_, _28681_, _12224_);
  or _79705_ (_28683_, _28682_, _12345_);
  or _79706_ (_28684_, _28683_, _28680_);
  or _79707_ (_28685_, _28587_, _12344_);
  and _79708_ (_28686_, _28685_, _06446_);
  and _79709_ (_28687_, _28686_, _28684_);
  and _79710_ (_28689_, _12224_, _06447_);
  or _79711_ (_28690_, _28689_, _25285_);
  or _79712_ (_28691_, _28690_, _12671_);
  or _79713_ (_28692_, _28691_, _28687_);
  or _79714_ (_28693_, _28587_, _12339_);
  and _79715_ (_28694_, _28693_, _12336_);
  and _79716_ (_28695_, _28694_, _28692_);
  and _79717_ (_28696_, _12224_, _12337_);
  or _79718_ (_28697_, _28696_, _06042_);
  or _79719_ (_28698_, _28697_, _28695_);
  nand _79720_ (_28700_, _28588_, _06042_);
  and _79721_ (_28701_, _28700_, _06340_);
  and _79722_ (_28702_, _28701_, _28698_);
  nand _79723_ (_28703_, _12224_, _06339_);
  nand _79724_ (_28704_, _28703_, _28069_);
  or _79725_ (_28705_, _28704_, _28702_);
  nand _79726_ (_28706_, _12401_, _06486_);
  and _79727_ (_28707_, _28706_, _06334_);
  and _79728_ (_28708_, _28707_, _28705_);
  and _79729_ (_28709_, _12224_, _14022_);
  or _79730_ (_28711_, _28709_, _06037_);
  or _79731_ (_28712_, _28711_, _28708_);
  nand _79732_ (_28713_, _12401_, _06037_);
  and _79733_ (_28714_, _28713_, _12694_);
  and _79734_ (_28715_, _28714_, _28712_);
  or _79735_ (_28716_, _28715_, _28590_);
  and _79736_ (_28717_, _28716_, _25604_);
  nand _79737_ (_28718_, _12224_, _06401_);
  nand _79738_ (_28719_, _28718_, _27945_);
  or _79739_ (_28720_, _28719_, _28717_);
  or _79740_ (_28722_, _28601_, _12705_);
  and _79741_ (_28723_, _28722_, _08626_);
  and _79742_ (_28724_, _28723_, _28720_);
  and _79743_ (_28725_, _12224_, _08848_);
  or _79744_ (_28726_, _28725_, _06277_);
  or _79745_ (_28727_, _28726_, _28724_);
  nand _79746_ (_28728_, _12401_, _06277_);
  and _79747_ (_28729_, _28728_, _11029_);
  and _79748_ (_28730_, _28729_, _28727_);
  and _79749_ (_28731_, _12224_, _11028_);
  or _79750_ (_28733_, _28731_, _12718_);
  or _79751_ (_28734_, _28733_, _28730_);
  nor _79752_ (_28735_, _12751_, \oc8051_golden_model_1.DPH [2]);
  nor _79753_ (_28736_, _28735_, _12752_);
  or _79754_ (_28737_, _28736_, _12719_);
  and _79755_ (_28738_, _28737_, _06958_);
  and _79756_ (_28739_, _28738_, _28734_);
  and _79757_ (_28740_, _12224_, _06400_);
  or _79758_ (_28741_, _28740_, _28739_);
  nor _79759_ (_28742_, _12763_, _06275_);
  and _79760_ (_28744_, _28742_, _28741_);
  or _79761_ (_28745_, _28601_, _11389_);
  or _79762_ (_28746_, _12224_, _12770_);
  and _79763_ (_28747_, _28746_, _12763_);
  and _79764_ (_28748_, _28747_, _28745_);
  or _79765_ (_28749_, _28748_, _12768_);
  or _79766_ (_28750_, _28749_, _28744_);
  or _79767_ (_28751_, _28587_, _12333_);
  and _79768_ (_28752_, _28751_, _12330_);
  and _79769_ (_28753_, _28752_, _28750_);
  and _79770_ (_28755_, _12224_, _12331_);
  or _79771_ (_28756_, _28755_, _06502_);
  or _79772_ (_28757_, _28756_, _28753_);
  nand _79773_ (_28758_, _12401_, _06502_);
  and _79774_ (_28759_, _28758_, _28757_);
  or _79775_ (_28760_, _28759_, _06615_);
  or _79776_ (_28761_, _12224_, _07337_);
  nor _79777_ (_28762_, _12787_, _12782_);
  and _79778_ (_28763_, _28762_, _28761_);
  and _79779_ (_28764_, _28763_, _28760_);
  or _79780_ (_28766_, _28601_, _12770_);
  or _79781_ (_28767_, _12224_, _11389_);
  and _79782_ (_28768_, _28767_, _12787_);
  and _79783_ (_28769_, _28768_, _28766_);
  or _79784_ (_28770_, _28769_, _12792_);
  or _79785_ (_28771_, _28770_, _28764_);
  or _79786_ (_28772_, _28587_, _12328_);
  and _79787_ (_28773_, _28772_, _12322_);
  and _79788_ (_28774_, _28773_, _28771_);
  and _79789_ (_28775_, _12224_, _12323_);
  or _79790_ (_28777_, _28775_, _06507_);
  or _79791_ (_28778_, _28777_, _28774_);
  and _79792_ (_28779_, _28778_, _28585_);
  or _79793_ (_28780_, _28779_, _06610_);
  or _79794_ (_28781_, _12224_, _07331_);
  and _79795_ (_28782_, _28781_, _28150_);
  and _79796_ (_28783_, _28782_, _28780_);
  or _79797_ (_28784_, _28601_, \oc8051_golden_model_1.PSW [7]);
  or _79798_ (_28785_, _12224_, _10967_);
  and _79799_ (_28786_, _28785_, _12809_);
  and _79800_ (_28788_, _28786_, _28784_);
  or _79801_ (_28789_, _28788_, _12814_);
  or _79802_ (_28790_, _28789_, _28783_);
  or _79803_ (_28791_, _28587_, _12320_);
  and _79804_ (_28792_, _28791_, _12314_);
  and _79805_ (_28793_, _28792_, _28790_);
  and _79806_ (_28794_, _12224_, _12315_);
  or _79807_ (_28795_, _28794_, _06509_);
  or _79808_ (_28796_, _28795_, _28793_);
  nand _79809_ (_28797_, _12401_, _06509_);
  and _79810_ (_28799_, _28797_, _28796_);
  or _79811_ (_28800_, _28799_, _06602_);
  or _79812_ (_28801_, _12224_, _09112_);
  and _79813_ (_28802_, _28801_, _28171_);
  and _79814_ (_28803_, _28802_, _28800_);
  or _79815_ (_28804_, _28601_, _10967_);
  or _79816_ (_28805_, _12224_, \oc8051_golden_model_1.PSW [7]);
  and _79817_ (_28806_, _28805_, _12310_);
  and _79818_ (_28807_, _28806_, _28804_);
  or _79819_ (_28808_, _28807_, _12839_);
  or _79820_ (_28810_, _28808_, _28803_);
  or _79821_ (_28811_, _28587_, _12837_);
  and _79822_ (_28812_, _28811_, _11187_);
  and _79823_ (_28813_, _28812_, _28810_);
  and _79824_ (_28814_, _12224_, _11188_);
  or _79825_ (_28815_, _28814_, _11216_);
  or _79826_ (_28816_, _28815_, _28813_);
  nand _79827_ (_28817_, _28588_, _11216_);
  and _79828_ (_28818_, _28817_, _28816_);
  or _79829_ (_28819_, _28818_, _06621_);
  nand _79830_ (_28821_, _07854_, _06621_);
  and _79831_ (_28822_, _28821_, _28519_);
  and _79832_ (_28823_, _28822_, _28819_);
  or _79833_ (_28824_, _28593_, _13038_);
  or _79834_ (_28825_, _12400_, _13037_);
  and _79835_ (_28826_, _28825_, _06512_);
  and _79836_ (_28827_, _28826_, _28824_);
  or _79837_ (_28828_, _28827_, _12854_);
  or _79838_ (_28829_, _28828_, _28823_);
  or _79839_ (_28830_, _28587_, _12201_);
  and _79840_ (_28832_, _28830_, _13046_);
  and _79841_ (_28833_, _28832_, _28829_);
  and _79842_ (_28834_, _13047_, _12224_);
  or _79843_ (_28835_, _28834_, _10564_);
  or _79844_ (_28836_, _28835_, _28833_);
  nand _79845_ (_28837_, _28588_, _10564_);
  and _79846_ (_28838_, _28837_, _28836_);
  or _79847_ (_28839_, _28838_, _06361_);
  nand _79848_ (_28840_, _07854_, _06361_);
  and _79849_ (_28841_, _28840_, _28540_);
  and _79850_ (_28843_, _28841_, _28839_);
  or _79851_ (_28844_, _28593_, _13037_);
  nand _79852_ (_28845_, _12401_, _13037_);
  and _79853_ (_28846_, _28845_, _28844_);
  and _79854_ (_28847_, _28846_, _06496_);
  or _79855_ (_28848_, _28847_, _13062_);
  or _79856_ (_28849_, _28848_, _28843_);
  or _79857_ (_28850_, _28587_, _09123_);
  and _79858_ (_28851_, _28850_, _28849_);
  or _79859_ (_28852_, _28851_, _06639_);
  or _79860_ (_28853_, _12224_, _07048_);
  and _79861_ (_28854_, _28853_, _13072_);
  and _79862_ (_28855_, _28854_, _28852_);
  nor _79863_ (_28856_, _28588_, _13072_);
  or _79864_ (_28857_, _28856_, _06503_);
  or _79865_ (_28858_, _28857_, _28855_);
  nand _79866_ (_28859_, _06727_, _06503_);
  and _79867_ (_28860_, _28859_, _28234_);
  and _79868_ (_28861_, _28860_, _28858_);
  and _79869_ (_28862_, _28846_, _05989_);
  or _79870_ (_28865_, _28862_, _13088_);
  or _79871_ (_28866_, _28865_, _28861_);
  or _79872_ (_28867_, _28587_, _13087_);
  and _79873_ (_28868_, _28867_, _28866_);
  or _79874_ (_28869_, _28868_, _06646_);
  or _79875_ (_28870_, _12224_, _06651_);
  and _79876_ (_28871_, _28870_, _13095_);
  and _79877_ (_28872_, _28871_, _28869_);
  nor _79878_ (_28873_, _28588_, _13095_);
  or _79879_ (_28874_, _28873_, _06488_);
  or _79880_ (_28876_, _28874_, _28872_);
  nand _79881_ (_28877_, _06727_, _06488_);
  and _79882_ (_28878_, _28877_, _28251_);
  and _79883_ (_28879_, _28878_, _28876_);
  and _79884_ (_28880_, _28587_, _13105_);
  or _79885_ (_28881_, _28880_, _28879_);
  or _79886_ (_28882_, _28881_, _01446_);
  or _79887_ (_28883_, _01442_, \oc8051_golden_model_1.PC [10]);
  and _79888_ (_28884_, _28883_, _43634_);
  and _79889_ (_44217_, _28884_, _28882_);
  nor _79890_ (_28886_, _12193_, \oc8051_golden_model_1.PC [11]);
  nor _79891_ (_28887_, _28886_, _12194_);
  or _79892_ (_28888_, _28887_, _12201_);
  or _79893_ (_28889_, _28887_, _12320_);
  or _79894_ (_28890_, _28887_, _12328_);
  or _79895_ (_28891_, _28887_, _12333_);
  or _79896_ (_28892_, _12220_, _08626_);
  and _79897_ (_28893_, _12395_, _06037_);
  or _79898_ (_28894_, _12397_, _12398_);
  nand _79899_ (_28895_, _28894_, _12477_);
  or _79900_ (_28897_, _28894_, _12477_);
  and _79901_ (_28898_, _28897_, _28895_);
  or _79902_ (_28899_, _28898_, _12648_);
  nand _79903_ (_28900_, _12648_, _12396_);
  and _79904_ (_28901_, _28900_, _06490_);
  and _79905_ (_28902_, _28901_, _28899_);
  nor _79906_ (_28903_, _12396_, _12379_);
  and _79907_ (_28904_, _28898_, _12379_);
  or _79908_ (_28905_, _28904_, _28903_);
  or _79909_ (_28906_, _28905_, _06473_);
  and _79910_ (_28908_, _12220_, _06417_);
  or _79911_ (_28909_, _28887_, _07270_);
  or _79912_ (_28910_, _12221_, _12222_);
  nand _79913_ (_28911_, _28910_, _12291_);
  or _79914_ (_28912_, _28910_, _12291_);
  and _79915_ (_28913_, _28912_, _28911_);
  and _79916_ (_28914_, _28913_, _12537_);
  and _79917_ (_28915_, _12539_, _12220_);
  or _79918_ (_28916_, _28915_, _28914_);
  and _79919_ (_28917_, _28916_, _08687_);
  or _79920_ (_28919_, _28887_, _12520_);
  and _79921_ (_28920_, _12523_, _15329_);
  nor _79922_ (_28921_, _06816_, \oc8051_golden_model_1.PC [11]);
  and _79923_ (_28922_, _28921_, _12525_);
  and _79924_ (_28923_, _28922_, _12518_);
  or _79925_ (_28924_, _28923_, _28920_);
  nand _79926_ (_28925_, _28924_, _12516_);
  and _79927_ (_28926_, _28925_, _08685_);
  and _79928_ (_28927_, _28926_, _28919_);
  or _79929_ (_28928_, _28927_, _07269_);
  or _79930_ (_28930_, _28928_, _28917_);
  and _79931_ (_28931_, _28930_, _28909_);
  and _79932_ (_28932_, _28931_, _07275_);
  and _79933_ (_28933_, _12512_, _12395_);
  and _79934_ (_28934_, _28898_, _12510_);
  or _79935_ (_28935_, _28934_, _28933_);
  and _79936_ (_28936_, _28935_, _06474_);
  or _79937_ (_28937_, _28936_, _28932_);
  or _79938_ (_28938_, _28937_, _25228_);
  or _79939_ (_28939_, _28887_, _12502_);
  and _79940_ (_28941_, _28939_, _12549_);
  and _79941_ (_28942_, _28941_, _28938_);
  nor _79942_ (_28943_, _12549_, _15329_);
  or _79943_ (_28944_, _28943_, _12552_);
  or _79944_ (_28945_, _28944_, _28942_);
  or _79945_ (_28946_, _28887_, _12551_);
  and _79946_ (_28947_, _28946_, _06426_);
  and _79947_ (_28948_, _28947_, _28945_);
  or _79948_ (_28949_, _28948_, _28908_);
  and _79949_ (_28950_, _28949_, _12561_);
  and _79950_ (_28952_, _28887_, _12563_);
  or _79951_ (_28953_, _28952_, _12568_);
  or _79952_ (_28954_, _28953_, _28950_);
  or _79953_ (_28955_, _12567_, _12220_);
  and _79954_ (_28956_, _28955_, _12574_);
  and _79955_ (_28957_, _28956_, _28954_);
  nand _79956_ (_28958_, _12609_, _12396_);
  or _79957_ (_28959_, _28898_, _12609_);
  and _79958_ (_28960_, _28959_, _12611_);
  and _79959_ (_28961_, _28960_, _28958_);
  or _79960_ (_28963_, _28961_, _06472_);
  or _79961_ (_28964_, _28963_, _28957_);
  and _79962_ (_28965_, _28964_, _28906_);
  or _79963_ (_28966_, _28965_, _06431_);
  and _79964_ (_28967_, _12630_, _12395_);
  and _79965_ (_28968_, _28898_, _12632_);
  or _79966_ (_28969_, _28968_, _06500_);
  or _79967_ (_28970_, _28969_, _28967_);
  and _79968_ (_28971_, _28970_, _12349_);
  and _79969_ (_28972_, _28971_, _28966_);
  or _79970_ (_28974_, _28972_, _28902_);
  and _79971_ (_28975_, _28974_, _12348_);
  nand _79972_ (_28976_, _28887_, _12347_);
  nand _79973_ (_28977_, _28976_, _12662_);
  or _79974_ (_28978_, _28977_, _28975_);
  or _79975_ (_28979_, _12662_, _12220_);
  and _79976_ (_28980_, _28979_, _12344_);
  and _79977_ (_28981_, _28980_, _28978_);
  not _79978_ (_28982_, _12669_);
  and _79979_ (_28983_, _28887_, _12345_);
  or _79980_ (_28985_, _28983_, _28982_);
  or _79981_ (_28986_, _28985_, _28981_);
  or _79982_ (_28987_, _12669_, _12220_);
  and _79983_ (_28988_, _28987_, _12339_);
  and _79984_ (_28989_, _28988_, _28986_);
  and _79985_ (_28990_, _28887_, _12671_);
  or _79986_ (_28991_, _28990_, _12337_);
  or _79987_ (_28992_, _28991_, _28989_);
  or _79988_ (_28993_, _12220_, _12336_);
  and _79989_ (_28994_, _28993_, _06043_);
  and _79990_ (_28996_, _28994_, _28992_);
  nand _79991_ (_28997_, _28887_, _06042_);
  nand _79992_ (_28998_, _28997_, _12681_);
  or _79993_ (_28999_, _28998_, _28996_);
  or _79994_ (_29000_, _12681_, _12220_);
  and _79995_ (_29001_, _29000_, _06487_);
  and _79996_ (_29002_, _29001_, _28999_);
  nand _79997_ (_29003_, _12395_, _06486_);
  nand _79998_ (_29004_, _29003_, _06334_);
  or _79999_ (_29005_, _29004_, _29002_);
  or _80000_ (_29007_, _12220_, _06334_);
  and _80001_ (_29008_, _29007_, _06313_);
  and _80002_ (_29009_, _29008_, _29005_);
  or _80003_ (_29010_, _29009_, _28893_);
  and _80004_ (_29011_, _29010_, _12694_);
  and _80005_ (_29012_, _28887_, _12700_);
  or _80006_ (_29013_, _29012_, _12698_);
  or _80007_ (_29014_, _29013_, _29011_);
  or _80008_ (_29015_, _12697_, _12220_);
  and _80009_ (_29016_, _29015_, _12705_);
  and _80010_ (_29018_, _29016_, _29014_);
  and _80011_ (_29019_, _28913_, _12704_);
  or _80012_ (_29020_, _29019_, _08848_);
  or _80013_ (_29021_, _29020_, _29018_);
  and _80014_ (_29022_, _29021_, _28892_);
  or _80015_ (_29023_, _29022_, _06277_);
  nand _80016_ (_29024_, _12396_, _06277_);
  and _80017_ (_29025_, _29024_, _11029_);
  and _80018_ (_29026_, _29025_, _29023_);
  and _80019_ (_29027_, _12220_, _11028_);
  or _80020_ (_29029_, _29027_, _29026_);
  and _80021_ (_29030_, _29029_, _12719_);
  or _80022_ (_29031_, _12752_, \oc8051_golden_model_1.DPH [3]);
  nor _80023_ (_29032_, _12753_, _12719_);
  and _80024_ (_29033_, _29032_, _29031_);
  or _80025_ (_29034_, _29033_, _12725_);
  or _80026_ (_29035_, _29034_, _29030_);
  or _80027_ (_29036_, _12724_, _12220_);
  and _80028_ (_29037_, _29036_, _12764_);
  and _80029_ (_29038_, _29037_, _29035_);
  or _80030_ (_29040_, _28913_, _11389_);
  or _80031_ (_29041_, _12220_, _12770_);
  and _80032_ (_29042_, _29041_, _12763_);
  and _80033_ (_29043_, _29042_, _29040_);
  or _80034_ (_29044_, _29043_, _12768_);
  or _80035_ (_29045_, _29044_, _29038_);
  and _80036_ (_29046_, _29045_, _28891_);
  or _80037_ (_29047_, _29046_, _12331_);
  or _80038_ (_29048_, _12220_, _12330_);
  and _80039_ (_29049_, _29048_, _07334_);
  and _80040_ (_29051_, _29049_, _29047_);
  nand _80041_ (_29052_, _12395_, _06502_);
  nand _80042_ (_29053_, _29052_, _12783_);
  or _80043_ (_29054_, _29053_, _29051_);
  or _80044_ (_29055_, _12783_, _12220_);
  and _80045_ (_29056_, _29055_, _12788_);
  and _80046_ (_29057_, _29056_, _29054_);
  or _80047_ (_29058_, _28913_, _12770_);
  or _80048_ (_29059_, _12220_, _11389_);
  and _80049_ (_29060_, _29059_, _12787_);
  and _80050_ (_29062_, _29060_, _29058_);
  or _80051_ (_29063_, _29062_, _12792_);
  or _80052_ (_29064_, _29063_, _29057_);
  and _80053_ (_29065_, _29064_, _28890_);
  or _80054_ (_29066_, _29065_, _12323_);
  or _80055_ (_29067_, _12220_, _12322_);
  and _80056_ (_29068_, _29067_, _07339_);
  and _80057_ (_29069_, _29068_, _29066_);
  nand _80058_ (_29070_, _12395_, _06507_);
  nand _80059_ (_29071_, _29070_, _12805_);
  or _80060_ (_29073_, _29071_, _29069_);
  or _80061_ (_29074_, _12805_, _12220_);
  and _80062_ (_29075_, _29074_, _12810_);
  and _80063_ (_29076_, _29075_, _29073_);
  or _80064_ (_29077_, _28913_, \oc8051_golden_model_1.PSW [7]);
  or _80065_ (_29078_, _12220_, _10967_);
  and _80066_ (_29079_, _29078_, _12809_);
  and _80067_ (_29080_, _29079_, _29077_);
  or _80068_ (_29081_, _29080_, _12814_);
  or _80069_ (_29082_, _29081_, _29076_);
  and _80070_ (_29084_, _29082_, _28889_);
  or _80071_ (_29085_, _29084_, _12315_);
  or _80072_ (_29086_, _12220_, _12314_);
  and _80073_ (_29087_, _29086_, _09107_);
  and _80074_ (_29088_, _29087_, _29085_);
  nand _80075_ (_29089_, _12395_, _06509_);
  nand _80076_ (_29090_, _29089_, _12828_);
  or _80077_ (_29091_, _29090_, _29088_);
  or _80078_ (_29092_, _12828_, _12220_);
  and _80079_ (_29093_, _29092_, _12832_);
  and _80080_ (_29095_, _29093_, _29091_);
  or _80081_ (_29096_, _28913_, _10967_);
  or _80082_ (_29097_, _12220_, \oc8051_golden_model_1.PSW [7]);
  and _80083_ (_29098_, _29097_, _12310_);
  and _80084_ (_29099_, _29098_, _29096_);
  or _80085_ (_29100_, _29099_, _29095_);
  and _80086_ (_29101_, _29100_, _12837_);
  and _80087_ (_29102_, _28887_, _12839_);
  or _80088_ (_29103_, _29102_, _11188_);
  or _80089_ (_29104_, _29103_, _29101_);
  or _80090_ (_29106_, _12220_, _11187_);
  and _80091_ (_29107_, _29106_, _11217_);
  and _80092_ (_29108_, _29107_, _29104_);
  and _80093_ (_29109_, _28887_, _11216_);
  or _80094_ (_29110_, _29109_, _06621_);
  or _80095_ (_29111_, _29110_, _29108_);
  nand _80096_ (_29112_, _07680_, _06621_);
  and _80097_ (_29113_, _29112_, _29111_);
  or _80098_ (_29114_, _29113_, _07350_);
  nor _80099_ (_29115_, _12220_, _06016_);
  nor _80100_ (_29117_, _29115_, _06512_);
  and _80101_ (_29118_, _29117_, _29114_);
  or _80102_ (_29119_, _28898_, _13038_);
  or _80103_ (_29120_, _12395_, _13037_);
  and _80104_ (_29121_, _29120_, _06512_);
  and _80105_ (_29122_, _29121_, _29119_);
  or _80106_ (_29123_, _29122_, _12854_);
  or _80107_ (_29124_, _29123_, _29118_);
  and _80108_ (_29125_, _29124_, _28888_);
  or _80109_ (_29126_, _29125_, _13047_);
  or _80110_ (_29128_, _13046_, _12220_);
  and _80111_ (_29129_, _29128_, _13049_);
  and _80112_ (_29130_, _29129_, _29126_);
  and _80113_ (_29131_, _28887_, _10564_);
  or _80114_ (_29132_, _29131_, _06361_);
  or _80115_ (_29133_, _29132_, _29130_);
  nand _80116_ (_29134_, _07680_, _06361_);
  and _80117_ (_29135_, _29134_, _29133_);
  or _80118_ (_29136_, _29135_, _12187_);
  nor _80119_ (_29137_, _12220_, _06021_);
  nor _80120_ (_29139_, _29137_, _06496_);
  and _80121_ (_29140_, _29139_, _29136_);
  nand _80122_ (_29141_, _12396_, _13037_);
  or _80123_ (_29142_, _28898_, _13037_);
  and _80124_ (_29143_, _29142_, _29141_);
  and _80125_ (_29144_, _29143_, _06496_);
  or _80126_ (_29145_, _29144_, _13062_);
  or _80127_ (_29146_, _29145_, _29140_);
  or _80128_ (_29147_, _28887_, _09123_);
  and _80129_ (_29148_, _29147_, _07048_);
  and _80130_ (_29150_, _29148_, _29146_);
  nand _80131_ (_29151_, _12220_, _06639_);
  nand _80132_ (_29152_, _29151_, _13072_);
  or _80133_ (_29153_, _29152_, _29150_);
  or _80134_ (_29154_, _28887_, _13072_);
  and _80135_ (_29155_, _29154_, _09534_);
  and _80136_ (_29156_, _29155_, _29153_);
  nor _80137_ (_29157_, _09534_, _06269_);
  or _80138_ (_29158_, _29157_, _05998_);
  or _80139_ (_29159_, _29158_, _29156_);
  nand _80140_ (_29161_, _15329_, _05998_);
  and _80141_ (_29162_, _29161_, _05990_);
  and _80142_ (_29163_, _29162_, _29159_);
  and _80143_ (_29164_, _29143_, _05989_);
  or _80144_ (_29165_, _29164_, _13088_);
  or _80145_ (_29166_, _29165_, _29163_);
  or _80146_ (_29167_, _28887_, _13087_);
  and _80147_ (_29168_, _29167_, _06651_);
  and _80148_ (_29169_, _29168_, _29166_);
  nand _80149_ (_29170_, _12220_, _06646_);
  nand _80150_ (_29172_, _29170_, _13095_);
  or _80151_ (_29173_, _29172_, _29169_);
  or _80152_ (_29174_, _28887_, _13095_);
  and _80153_ (_29175_, _29174_, _13098_);
  and _80154_ (_29176_, _29175_, _29173_);
  nor _80155_ (_29177_, _13098_, _06269_);
  or _80156_ (_29178_, _29177_, _05997_);
  or _80157_ (_29179_, _29178_, _29176_);
  nand _80158_ (_29180_, _15329_, _05997_);
  and _80159_ (_29181_, _29180_, _13106_);
  and _80160_ (_29183_, _29181_, _29179_);
  and _80161_ (_29184_, _28887_, _13105_);
  or _80162_ (_29185_, _29184_, _29183_);
  or _80163_ (_29186_, _29185_, _01446_);
  or _80164_ (_29187_, _01442_, \oc8051_golden_model_1.PC [11]);
  and _80165_ (_29188_, _29187_, _43634_);
  and _80166_ (_44218_, _29188_, _29186_);
  and _80167_ (_29189_, _12190_, _09536_);
  and _80168_ (_29190_, _29189_, \oc8051_golden_model_1.PC [11]);
  and _80169_ (_29191_, _29190_, \oc8051_golden_model_1.PC [12]);
  nor _80170_ (_29193_, _29190_, \oc8051_golden_model_1.PC [12]);
  nor _80171_ (_29194_, _29193_, _29191_);
  not _80172_ (_29195_, _29194_);
  and _80173_ (_29196_, _29195_, _10564_);
  nor _80174_ (_29197_, _12828_, _15533_);
  nor _80175_ (_29198_, _12805_, _15533_);
  nor _80176_ (_29199_, _12783_, _15533_);
  nor _80177_ (_29200_, _12481_, _12479_);
  nor _80178_ (_29201_, _29200_, _12482_);
  not _80179_ (_29202_, _29201_);
  nand _80180_ (_29204_, _29202_, _12379_);
  or _80181_ (_29205_, _12391_, _12379_);
  and _80182_ (_29206_, _29205_, _06472_);
  and _80183_ (_29207_, _29206_, _29204_);
  nor _80184_ (_29208_, _29195_, _12561_);
  or _80185_ (_29209_, _29194_, _12551_);
  or _80186_ (_29210_, _12510_, _12391_);
  or _80187_ (_29211_, _29201_, _12512_);
  and _80188_ (_29212_, _29211_, _29210_);
  or _80189_ (_29213_, _29212_, _07275_);
  nor _80190_ (_29215_, _29195_, _12520_);
  and _80191_ (_29216_, _12523_, _12215_);
  and _80192_ (_29217_, _12518_, _07564_);
  and _80193_ (_29218_, _12525_, \oc8051_golden_model_1.PC [12]);
  and _80194_ (_29219_, _29218_, _29217_);
  or _80195_ (_29220_, _29219_, _29216_);
  and _80196_ (_29221_, _29220_, _12516_);
  or _80197_ (_29222_, _29221_, _08687_);
  or _80198_ (_29223_, _29222_, _29215_);
  and _80199_ (_29224_, _12539_, _12215_);
  nor _80200_ (_29226_, _12295_, _12293_);
  nor _80201_ (_29227_, _29226_, _12296_);
  and _80202_ (_29228_, _29227_, _12537_);
  or _80203_ (_29229_, _29228_, _29224_);
  or _80204_ (_29230_, _29229_, _08685_);
  and _80205_ (_29231_, _29230_, _29223_);
  or _80206_ (_29232_, _29231_, _27616_);
  and _80207_ (_29233_, _29232_, _29213_);
  or _80208_ (_29234_, _29233_, _25228_);
  or _80209_ (_29235_, _29194_, _12503_);
  and _80210_ (_29237_, _29235_, _12549_);
  and _80211_ (_29238_, _29237_, _29234_);
  nor _80212_ (_29239_, _12549_, _15533_);
  or _80213_ (_29240_, _29239_, _12552_);
  or _80214_ (_29241_, _29240_, _29238_);
  and _80215_ (_29242_, _29241_, _29209_);
  or _80216_ (_29243_, _29242_, _06417_);
  nand _80217_ (_29244_, _15533_, _06417_);
  and _80218_ (_29245_, _29244_, _12561_);
  and _80219_ (_29246_, _29245_, _29243_);
  or _80220_ (_29248_, _29246_, _29208_);
  and _80221_ (_29249_, _29248_, _12567_);
  or _80222_ (_29250_, _12567_, _15533_);
  nand _80223_ (_29251_, _29250_, _12574_);
  or _80224_ (_29252_, _29251_, _29249_);
  nor _80225_ (_29253_, _29202_, _12609_);
  and _80226_ (_29254_, _12609_, _12391_);
  or _80227_ (_29255_, _29254_, _12574_);
  or _80228_ (_29256_, _29255_, _29253_);
  and _80229_ (_29257_, _29256_, _06473_);
  and _80230_ (_29259_, _29257_, _29252_);
  or _80231_ (_29260_, _29259_, _06431_);
  or _80232_ (_29261_, _29260_, _29207_);
  nor _80233_ (_29262_, _29202_, _12630_);
  and _80234_ (_29263_, _12630_, _12391_);
  or _80235_ (_29264_, _29263_, _29262_);
  or _80236_ (_29265_, _29264_, _06500_);
  and _80237_ (_29266_, _29265_, _12349_);
  and _80238_ (_29267_, _29266_, _29261_);
  or _80239_ (_29268_, _29201_, _12648_);
  or _80240_ (_29270_, _26636_, _12391_);
  and _80241_ (_29271_, _29270_, _06490_);
  and _80242_ (_29272_, _29271_, _29268_);
  or _80243_ (_29273_, _29272_, _12347_);
  or _80244_ (_29274_, _29273_, _29267_);
  nand _80245_ (_29275_, _29195_, _12347_);
  and _80246_ (_29276_, _29275_, _12662_);
  and _80247_ (_29277_, _29276_, _29274_);
  nor _80248_ (_29278_, _12662_, _15533_);
  or _80249_ (_29279_, _29278_, _12345_);
  or _80250_ (_29281_, _29279_, _29277_);
  or _80251_ (_29282_, _29194_, _12344_);
  and _80252_ (_29283_, _29282_, _12669_);
  and _80253_ (_29284_, _29283_, _29281_);
  nor _80254_ (_29285_, _12669_, _15533_);
  or _80255_ (_29286_, _29285_, _12671_);
  or _80256_ (_29287_, _29286_, _29284_);
  or _80257_ (_29288_, _29194_, _12339_);
  and _80258_ (_29289_, _29288_, _12336_);
  and _80259_ (_29290_, _29289_, _29287_);
  nor _80260_ (_29292_, _15533_, _12336_);
  or _80261_ (_29293_, _29292_, _06042_);
  or _80262_ (_29294_, _29293_, _29290_);
  nand _80263_ (_29295_, _29195_, _06042_);
  and _80264_ (_29296_, _29295_, _12681_);
  and _80265_ (_29297_, _29296_, _29294_);
  nor _80266_ (_29298_, _12681_, _15533_);
  or _80267_ (_29299_, _29298_, _06486_);
  or _80268_ (_29300_, _29299_, _29297_);
  or _80269_ (_29301_, _12391_, _06487_);
  and _80270_ (_29303_, _29301_, _06334_);
  and _80271_ (_29304_, _29303_, _29300_);
  nor _80272_ (_29305_, _15533_, _06334_);
  or _80273_ (_29306_, _29305_, _06037_);
  or _80274_ (_29307_, _29306_, _29304_);
  or _80275_ (_29308_, _12391_, _06313_);
  and _80276_ (_29309_, _29308_, _12694_);
  and _80277_ (_29310_, _29309_, _29307_);
  or _80278_ (_29311_, _29195_, _12694_);
  nand _80279_ (_29312_, _29311_, _12697_);
  or _80280_ (_29314_, _29312_, _29310_);
  or _80281_ (_29315_, _12697_, _12215_);
  and _80282_ (_29316_, _29315_, _12705_);
  and _80283_ (_29317_, _29316_, _29314_);
  and _80284_ (_29318_, _29227_, _12704_);
  or _80285_ (_29319_, _29318_, _29317_);
  nor _80286_ (_29320_, _29319_, _08848_);
  nor _80287_ (_29321_, _12215_, _08626_);
  nor _80288_ (_29322_, _29321_, _29320_);
  and _80289_ (_29323_, _29322_, _06278_);
  and _80290_ (_29325_, _12391_, _06277_);
  or _80291_ (_29326_, _29325_, _29323_);
  and _80292_ (_29327_, _29326_, _11029_);
  and _80293_ (_29328_, _12215_, _11028_);
  or _80294_ (_29329_, _29328_, _12718_);
  nor _80295_ (_29330_, _29329_, _29327_);
  nor _80296_ (_29331_, _12753_, \oc8051_golden_model_1.DPH [4]);
  nor _80297_ (_29332_, _29331_, _12754_);
  nor _80298_ (_29333_, _29332_, _12719_);
  nor _80299_ (_29334_, _29333_, _12725_);
  not _80300_ (_29336_, _29334_);
  nor _80301_ (_29337_, _29336_, _29330_);
  nor _80302_ (_29338_, _12724_, _15533_);
  or _80303_ (_29339_, _29338_, _29337_);
  nand _80304_ (_29340_, _29339_, _12764_);
  nor _80305_ (_29341_, _29227_, _11389_);
  nor _80306_ (_29342_, _12215_, _12770_);
  nor _80307_ (_29343_, _29342_, _12764_);
  not _80308_ (_29344_, _29343_);
  nor _80309_ (_29345_, _29344_, _29341_);
  nor _80310_ (_29347_, _29345_, _12768_);
  nand _80311_ (_29348_, _29347_, _29340_);
  nor _80312_ (_29349_, _29194_, _12333_);
  nor _80313_ (_29350_, _29349_, _12331_);
  nand _80314_ (_29351_, _29350_, _29348_);
  nor _80315_ (_29352_, _15533_, _12330_);
  nor _80316_ (_29353_, _29352_, _06502_);
  nand _80317_ (_29354_, _29353_, _29351_);
  nor _80318_ (_29355_, _12391_, _07334_);
  nor _80319_ (_29356_, _29355_, _12784_);
  and _80320_ (_29358_, _29356_, _29354_);
  or _80321_ (_29359_, _29358_, _29199_);
  nand _80322_ (_29360_, _29359_, _12788_);
  and _80323_ (_29361_, _12215_, _12770_);
  and _80324_ (_29362_, _29227_, _11389_);
  or _80325_ (_29363_, _29362_, _29361_);
  and _80326_ (_29364_, _29363_, _12787_);
  nor _80327_ (_29365_, _29364_, _12792_);
  nand _80328_ (_29366_, _29365_, _29360_);
  nor _80329_ (_29367_, _29194_, _12328_);
  nor _80330_ (_29369_, _29367_, _12323_);
  nand _80331_ (_29370_, _29369_, _29366_);
  nor _80332_ (_29371_, _15533_, _12322_);
  nor _80333_ (_29372_, _29371_, _06507_);
  nand _80334_ (_29373_, _29372_, _29370_);
  nor _80335_ (_29374_, _12391_, _07339_);
  nor _80336_ (_29375_, _29374_, _12806_);
  and _80337_ (_29376_, _29375_, _29373_);
  or _80338_ (_29377_, _29376_, _29198_);
  nand _80339_ (_29378_, _29377_, _12810_);
  nor _80340_ (_29379_, _29227_, \oc8051_golden_model_1.PSW [7]);
  nor _80341_ (_29380_, _12215_, _10967_);
  nor _80342_ (_29381_, _29380_, _12810_);
  not _80343_ (_29382_, _29381_);
  nor _80344_ (_29383_, _29382_, _29379_);
  nor _80345_ (_29384_, _29383_, _12814_);
  nand _80346_ (_29385_, _29384_, _29378_);
  nor _80347_ (_29386_, _29194_, _12320_);
  nor _80348_ (_29387_, _29386_, _12315_);
  nand _80349_ (_29388_, _29387_, _29385_);
  nor _80350_ (_29391_, _15533_, _12314_);
  nor _80351_ (_29392_, _29391_, _06509_);
  nand _80352_ (_29393_, _29392_, _29388_);
  nor _80353_ (_29394_, _12391_, _09107_);
  nor _80354_ (_29395_, _29394_, _12829_);
  and _80355_ (_29396_, _29395_, _29393_);
  or _80356_ (_29397_, _29396_, _29197_);
  nand _80357_ (_29398_, _29397_, _12832_);
  and _80358_ (_29399_, _12215_, _10967_);
  and _80359_ (_29400_, _29227_, \oc8051_golden_model_1.PSW [7]);
  or _80360_ (_29402_, _29400_, _29399_);
  and _80361_ (_29403_, _29402_, _12310_);
  nor _80362_ (_29404_, _29403_, _12839_);
  nand _80363_ (_29405_, _29404_, _29398_);
  nor _80364_ (_29406_, _29194_, _12837_);
  nor _80365_ (_29407_, _29406_, _11188_);
  nand _80366_ (_29408_, _29407_, _29405_);
  nor _80367_ (_29409_, _15533_, _11187_);
  nor _80368_ (_29410_, _29409_, _11216_);
  nand _80369_ (_29411_, _29410_, _29408_);
  and _80370_ (_29413_, _29195_, _11216_);
  nor _80371_ (_29414_, _29413_, _06621_);
  and _80372_ (_29415_, _29414_, _29411_);
  nor _80373_ (_29416_, _08596_, _14116_);
  or _80374_ (_29417_, _29416_, _07350_);
  or _80375_ (_29418_, _29417_, _29415_);
  nor _80376_ (_29419_, _12215_, _06016_);
  nor _80377_ (_29420_, _29419_, _06512_);
  nand _80378_ (_29421_, _29420_, _29418_);
  nor _80379_ (_29422_, _12391_, _13037_);
  and _80380_ (_29424_, _29202_, _13037_);
  or _80381_ (_29425_, _29424_, _06629_);
  or _80382_ (_29426_, _29425_, _29422_);
  and _80383_ (_29427_, _29426_, _12201_);
  nand _80384_ (_29428_, _29427_, _29421_);
  nor _80385_ (_29429_, _29194_, _12201_);
  nor _80386_ (_29430_, _29429_, _13047_);
  nand _80387_ (_29431_, _29430_, _29428_);
  nor _80388_ (_29432_, _13046_, _15533_);
  nor _80389_ (_29433_, _29432_, _10564_);
  and _80390_ (_29435_, _29433_, _29431_);
  or _80391_ (_29436_, _29435_, _29196_);
  nand _80392_ (_29437_, _29436_, _06362_);
  and _80393_ (_29438_, _08596_, _06361_);
  nor _80394_ (_29439_, _29438_, _12187_);
  and _80395_ (_29440_, _29439_, _29437_);
  nor _80396_ (_29441_, _15533_, _06021_);
  or _80397_ (_29442_, _29441_, _06496_);
  nor _80398_ (_29443_, _29442_, _29440_);
  and _80399_ (_29444_, _12391_, _13037_);
  nor _80400_ (_29446_, _29202_, _13037_);
  or _80401_ (_29447_, _29446_, _29444_);
  nor _80402_ (_29448_, _29447_, _07035_);
  or _80403_ (_29449_, _29448_, _29443_);
  and _80404_ (_29450_, _29449_, _09123_);
  nor _80405_ (_29451_, _29194_, _09123_);
  or _80406_ (_29452_, _29451_, _29450_);
  nand _80407_ (_29453_, _29452_, _07048_);
  nand _80408_ (_29454_, _15533_, _06639_);
  and _80409_ (_29455_, _29454_, _13072_);
  nand _80410_ (_29457_, _29455_, _29453_);
  nor _80411_ (_29458_, _29195_, _13072_);
  nor _80412_ (_29459_, _29458_, _06503_);
  nand _80413_ (_29460_, _29459_, _29457_);
  and _80414_ (_29461_, _07093_, _06503_);
  nor _80415_ (_29462_, _29461_, _05998_);
  and _80416_ (_29463_, _29462_, _29460_);
  and _80417_ (_29464_, _12215_, _05998_);
  or _80418_ (_29465_, _29464_, _05989_);
  or _80419_ (_29466_, _29465_, _29463_);
  nor _80420_ (_29468_, _29447_, _05990_);
  nor _80421_ (_29469_, _29468_, _13088_);
  nand _80422_ (_29470_, _29469_, _29466_);
  nor _80423_ (_29471_, _29195_, _13087_);
  nor _80424_ (_29472_, _29471_, _06646_);
  nand _80425_ (_29473_, _29472_, _29470_);
  and _80426_ (_29474_, _15533_, _06646_);
  nor _80427_ (_29475_, _29474_, _26866_);
  nand _80428_ (_29476_, _29475_, _29473_);
  nor _80429_ (_29477_, _29195_, _13095_);
  nor _80430_ (_29479_, _29477_, _06488_);
  and _80431_ (_29480_, _29479_, _29476_);
  and _80432_ (_29481_, _07093_, _06488_);
  or _80433_ (_29482_, _29481_, _05997_);
  nor _80434_ (_29483_, _29482_, _29480_);
  and _80435_ (_29484_, _12215_, _05997_);
  or _80436_ (_29485_, _29484_, _29483_);
  and _80437_ (_29486_, _29485_, _13106_);
  and _80438_ (_29487_, _29194_, _13105_);
  or _80439_ (_29488_, _29487_, _29486_);
  or _80440_ (_29490_, _29488_, _01446_);
  or _80441_ (_29491_, _01442_, \oc8051_golden_model_1.PC [12]);
  and _80442_ (_29492_, _29491_, _43634_);
  and _80443_ (_44219_, _29492_, _29490_);
  and _80444_ (_29493_, _29191_, \oc8051_golden_model_1.PC [13]);
  nor _80445_ (_29494_, _29191_, \oc8051_golden_model_1.PC [13]);
  nor _80446_ (_29495_, _29494_, _29493_);
  or _80447_ (_29496_, _29495_, _12201_);
  or _80448_ (_29497_, _12211_, _12212_);
  not _80449_ (_29498_, _29497_);
  nor _80450_ (_29500_, _29498_, _12297_);
  and _80451_ (_29501_, _29498_, _12297_);
  or _80452_ (_29502_, _29501_, _29500_);
  or _80453_ (_29503_, _29502_, _10967_);
  or _80454_ (_29504_, _12210_, \oc8051_golden_model_1.PSW [7]);
  and _80455_ (_29505_, _29504_, _12310_);
  and _80456_ (_29506_, _29505_, _29503_);
  or _80457_ (_29507_, _29495_, _12320_);
  or _80458_ (_29508_, _29495_, _12333_);
  or _80459_ (_29509_, _12210_, _08626_);
  and _80460_ (_29511_, _12386_, _06037_);
  or _80461_ (_29512_, _12387_, _12388_);
  not _80462_ (_29513_, _29512_);
  nor _80463_ (_29514_, _29513_, _12483_);
  and _80464_ (_29515_, _29513_, _12483_);
  or _80465_ (_29516_, _29515_, _29514_);
  or _80466_ (_29517_, _29516_, _12648_);
  or _80467_ (_29518_, _26636_, _12386_);
  and _80468_ (_29519_, _29518_, _06490_);
  and _80469_ (_29520_, _29519_, _29517_);
  not _80470_ (_29522_, _12379_);
  or _80471_ (_29523_, _29516_, _29522_);
  or _80472_ (_29524_, _12386_, _12379_);
  and _80473_ (_29525_, _29524_, _06472_);
  and _80474_ (_29526_, _29525_, _29523_);
  or _80475_ (_29527_, _12567_, _12210_);
  and _80476_ (_29528_, _12210_, _06417_);
  and _80477_ (_29529_, _29516_, _12510_);
  and _80478_ (_29530_, _12512_, _12386_);
  or _80479_ (_29531_, _29530_, _07275_);
  or _80480_ (_29533_, _29531_, _29529_);
  and _80481_ (_29534_, _12539_, _12210_);
  and _80482_ (_29535_, _29502_, _12537_);
  or _80483_ (_29536_, _29535_, _29534_);
  and _80484_ (_29537_, _29536_, _08687_);
  or _80485_ (_29538_, _29495_, _12520_);
  and _80486_ (_29539_, _12523_, _15729_);
  nor _80487_ (_29540_, _06816_, \oc8051_golden_model_1.PC [13]);
  and _80488_ (_29541_, _29540_, _12525_);
  and _80489_ (_29542_, _29541_, _12518_);
  or _80490_ (_29544_, _29542_, _29539_);
  nand _80491_ (_29545_, _29544_, _12516_);
  and _80492_ (_29546_, _29545_, _08685_);
  and _80493_ (_29547_, _29546_, _29538_);
  or _80494_ (_29548_, _29547_, _27616_);
  or _80495_ (_29549_, _29548_, _29537_);
  and _80496_ (_29550_, _29549_, _29533_);
  or _80497_ (_29551_, _29550_, _25228_);
  or _80498_ (_29552_, _29495_, _12503_);
  and _80499_ (_29553_, _29552_, _12549_);
  and _80500_ (_29555_, _29553_, _29551_);
  nor _80501_ (_29556_, _12549_, _15729_);
  or _80502_ (_29557_, _29556_, _12552_);
  or _80503_ (_29558_, _29557_, _29555_);
  or _80504_ (_29559_, _29495_, _12551_);
  and _80505_ (_29560_, _29559_, _06426_);
  and _80506_ (_29561_, _29560_, _29558_);
  or _80507_ (_29562_, _29561_, _29528_);
  and _80508_ (_29563_, _29562_, _12561_);
  not _80509_ (_29564_, _29495_);
  or _80510_ (_29566_, _29564_, _12561_);
  nand _80511_ (_29567_, _29566_, _12567_);
  or _80512_ (_29568_, _29567_, _29563_);
  and _80513_ (_29569_, _29568_, _29527_);
  or _80514_ (_29570_, _29569_, _12611_);
  and _80515_ (_29571_, _12609_, _12386_);
  and _80516_ (_29572_, _29516_, _14270_);
  or _80517_ (_29573_, _29572_, _29571_);
  or _80518_ (_29574_, _29573_, _12574_);
  and _80519_ (_29575_, _29574_, _06473_);
  and _80520_ (_29577_, _29575_, _29570_);
  or _80521_ (_29578_, _29577_, _06431_);
  or _80522_ (_29579_, _29578_, _29526_);
  and _80523_ (_29580_, _12630_, _12386_);
  and _80524_ (_29581_, _29516_, _12632_);
  or _80525_ (_29582_, _29581_, _06500_);
  or _80526_ (_29583_, _29582_, _29580_);
  and _80527_ (_29584_, _29583_, _12349_);
  and _80528_ (_29585_, _29584_, _29579_);
  or _80529_ (_29586_, _29585_, _29520_);
  and _80530_ (_29588_, _29586_, _12348_);
  nand _80531_ (_29589_, _29495_, _12347_);
  nand _80532_ (_29590_, _29589_, _12662_);
  or _80533_ (_29591_, _29590_, _29588_);
  or _80534_ (_29592_, _12662_, _12210_);
  and _80535_ (_29593_, _29592_, _12344_);
  and _80536_ (_29594_, _29593_, _29591_);
  nor _80537_ (_29595_, _29564_, _12344_);
  or _80538_ (_29596_, _29595_, _28982_);
  or _80539_ (_29597_, _29596_, _29594_);
  or _80540_ (_29599_, _12669_, _12210_);
  and _80541_ (_29600_, _29599_, _12339_);
  and _80542_ (_29601_, _29600_, _29597_);
  nor _80543_ (_29602_, _29564_, _12339_);
  or _80544_ (_29603_, _29602_, _12337_);
  or _80545_ (_29604_, _29603_, _29601_);
  or _80546_ (_29605_, _12210_, _12336_);
  and _80547_ (_29606_, _29605_, _06043_);
  and _80548_ (_29607_, _29606_, _29604_);
  nand _80549_ (_29608_, _29495_, _06042_);
  nand _80550_ (_29610_, _29608_, _12681_);
  or _80551_ (_29611_, _29610_, _29607_);
  or _80552_ (_29612_, _12681_, _12210_);
  and _80553_ (_29613_, _29612_, _06487_);
  and _80554_ (_29614_, _29613_, _29611_);
  nand _80555_ (_29615_, _12386_, _06486_);
  nand _80556_ (_29616_, _29615_, _06334_);
  or _80557_ (_29617_, _29616_, _29614_);
  or _80558_ (_29618_, _12210_, _06334_);
  and _80559_ (_29619_, _29618_, _06313_);
  and _80560_ (_29621_, _29619_, _29617_);
  or _80561_ (_29622_, _29621_, _29511_);
  and _80562_ (_29623_, _29622_, _12694_);
  or _80563_ (_29624_, _29564_, _12694_);
  nand _80564_ (_29625_, _29624_, _12697_);
  or _80565_ (_29626_, _29625_, _29623_);
  or _80566_ (_29627_, _12697_, _12210_);
  and _80567_ (_29628_, _29627_, _12705_);
  and _80568_ (_29629_, _29628_, _29626_);
  and _80569_ (_29630_, _29502_, _12704_);
  or _80570_ (_29632_, _29630_, _08848_);
  or _80571_ (_29633_, _29632_, _29629_);
  and _80572_ (_29634_, _29633_, _29509_);
  or _80573_ (_29635_, _29634_, _06277_);
  or _80574_ (_29636_, _12386_, _06278_);
  and _80575_ (_29637_, _29636_, _11029_);
  and _80576_ (_29638_, _29637_, _29635_);
  and _80577_ (_29639_, _12210_, _11028_);
  or _80578_ (_29640_, _29639_, _29638_);
  and _80579_ (_29641_, _29640_, _12719_);
  or _80580_ (_29643_, _12754_, \oc8051_golden_model_1.DPH [5]);
  nor _80581_ (_29644_, _12755_, _12719_);
  and _80582_ (_29645_, _29644_, _29643_);
  or _80583_ (_29646_, _29645_, _12725_);
  or _80584_ (_29647_, _29646_, _29641_);
  or _80585_ (_29648_, _12724_, _12210_);
  and _80586_ (_29649_, _29648_, _12764_);
  and _80587_ (_29650_, _29649_, _29647_);
  or _80588_ (_29651_, _29502_, _11389_);
  or _80589_ (_29652_, _12210_, _12770_);
  and _80590_ (_29653_, _29652_, _12763_);
  and _80591_ (_29654_, _29653_, _29651_);
  or _80592_ (_29655_, _29654_, _12768_);
  or _80593_ (_29656_, _29655_, _29650_);
  and _80594_ (_29657_, _29656_, _29508_);
  or _80595_ (_29658_, _29657_, _12331_);
  or _80596_ (_29659_, _12210_, _12330_);
  and _80597_ (_29660_, _29659_, _07334_);
  and _80598_ (_29661_, _29660_, _29658_);
  nand _80599_ (_29662_, _12386_, _06502_);
  nand _80600_ (_29665_, _29662_, _12783_);
  or _80601_ (_29666_, _29665_, _29661_);
  or _80602_ (_29667_, _12783_, _12210_);
  and _80603_ (_29668_, _29667_, _12788_);
  and _80604_ (_29669_, _29668_, _29666_);
  or _80605_ (_29670_, _29502_, _12770_);
  or _80606_ (_29671_, _12210_, _11389_);
  and _80607_ (_29672_, _29671_, _12787_);
  and _80608_ (_29673_, _29672_, _29670_);
  or _80609_ (_29674_, _29673_, _29669_);
  and _80610_ (_29676_, _29674_, _12328_);
  nor _80611_ (_29677_, _29564_, _12328_);
  or _80612_ (_29678_, _29677_, _12323_);
  or _80613_ (_29679_, _29678_, _29676_);
  or _80614_ (_29680_, _12210_, _12322_);
  and _80615_ (_29681_, _29680_, _07339_);
  and _80616_ (_29682_, _29681_, _29679_);
  nand _80617_ (_29683_, _12386_, _06507_);
  nand _80618_ (_29684_, _29683_, _12805_);
  or _80619_ (_29685_, _29684_, _29682_);
  or _80620_ (_29687_, _12805_, _12210_);
  and _80621_ (_29688_, _29687_, _12810_);
  and _80622_ (_29689_, _29688_, _29685_);
  or _80623_ (_29690_, _29502_, \oc8051_golden_model_1.PSW [7]);
  or _80624_ (_29691_, _12210_, _10967_);
  and _80625_ (_29692_, _29691_, _12809_);
  and _80626_ (_29693_, _29692_, _29690_);
  or _80627_ (_29694_, _29693_, _12814_);
  or _80628_ (_29695_, _29694_, _29689_);
  and _80629_ (_29696_, _29695_, _29507_);
  or _80630_ (_29698_, _29696_, _12315_);
  or _80631_ (_29699_, _12210_, _12314_);
  and _80632_ (_29700_, _29699_, _09107_);
  and _80633_ (_29701_, _29700_, _29698_);
  nand _80634_ (_29702_, _12386_, _06509_);
  nand _80635_ (_29703_, _29702_, _12828_);
  or _80636_ (_29704_, _29703_, _29701_);
  or _80637_ (_29705_, _12828_, _12210_);
  and _80638_ (_29706_, _29705_, _12832_);
  and _80639_ (_29707_, _29706_, _29704_);
  or _80640_ (_29709_, _29707_, _29506_);
  and _80641_ (_29710_, _29709_, _12837_);
  nor _80642_ (_29711_, _29564_, _12837_);
  or _80643_ (_29712_, _29711_, _11188_);
  or _80644_ (_29713_, _29712_, _29710_);
  or _80645_ (_29714_, _12210_, _11187_);
  and _80646_ (_29715_, _29714_, _11217_);
  and _80647_ (_29716_, _29715_, _29713_);
  and _80648_ (_29717_, _29495_, _11216_);
  or _80649_ (_29718_, _29717_, _06621_);
  or _80650_ (_29720_, _29718_, _29716_);
  nand _80651_ (_29721_, _08305_, _06621_);
  and _80652_ (_29722_, _29721_, _29720_);
  or _80653_ (_29723_, _29722_, _07350_);
  nor _80654_ (_29724_, _12210_, _06016_);
  nor _80655_ (_29725_, _29724_, _06512_);
  and _80656_ (_29726_, _29725_, _29723_);
  or _80657_ (_29727_, _29516_, _13038_);
  or _80658_ (_29728_, _12386_, _13037_);
  and _80659_ (_29729_, _29728_, _06512_);
  and _80660_ (_29731_, _29729_, _29727_);
  or _80661_ (_29732_, _29731_, _12854_);
  or _80662_ (_29733_, _29732_, _29726_);
  and _80663_ (_29734_, _29733_, _29496_);
  or _80664_ (_29735_, _29734_, _13047_);
  or _80665_ (_29736_, _13046_, _12210_);
  and _80666_ (_29737_, _29736_, _13049_);
  and _80667_ (_29738_, _29737_, _29735_);
  and _80668_ (_29739_, _29495_, _10564_);
  or _80669_ (_29740_, _29739_, _06361_);
  or _80670_ (_29742_, _29740_, _29738_);
  nand _80671_ (_29743_, _08305_, _06361_);
  and _80672_ (_29744_, _29743_, _29742_);
  or _80673_ (_29745_, _29744_, _12187_);
  nor _80674_ (_29746_, _12210_, _06021_);
  nor _80675_ (_29747_, _29746_, _06496_);
  and _80676_ (_29748_, _29747_, _29745_);
  or _80677_ (_29749_, _29516_, _13037_);
  or _80678_ (_29750_, _12386_, _13038_);
  and _80679_ (_29751_, _29750_, _29749_);
  and _80680_ (_29753_, _29751_, _06496_);
  or _80681_ (_29754_, _29753_, _13062_);
  or _80682_ (_29755_, _29754_, _29748_);
  or _80683_ (_29756_, _29495_, _09123_);
  and _80684_ (_29757_, _29756_, _07048_);
  and _80685_ (_29758_, _29757_, _29755_);
  nand _80686_ (_29759_, _12210_, _06639_);
  nand _80687_ (_29760_, _29759_, _13072_);
  or _80688_ (_29761_, _29760_, _29758_);
  or _80689_ (_29762_, _29495_, _13072_);
  and _80690_ (_29764_, _29762_, _09534_);
  and _80691_ (_29765_, _29764_, _29761_);
  nor _80692_ (_29766_, _06685_, _09534_);
  or _80693_ (_29767_, _29766_, _05998_);
  or _80694_ (_29768_, _29767_, _29765_);
  nand _80695_ (_29769_, _15729_, _05998_);
  and _80696_ (_29770_, _29769_, _05990_);
  and _80697_ (_29771_, _29770_, _29768_);
  and _80698_ (_29772_, _29751_, _05989_);
  or _80699_ (_29773_, _29772_, _13088_);
  or _80700_ (_29775_, _29773_, _29771_);
  or _80701_ (_29776_, _29495_, _13087_);
  and _80702_ (_29777_, _29776_, _06651_);
  and _80703_ (_29778_, _29777_, _29775_);
  nand _80704_ (_29779_, _12210_, _06646_);
  nand _80705_ (_29780_, _29779_, _13095_);
  or _80706_ (_29781_, _29780_, _29778_);
  or _80707_ (_29782_, _29495_, _13095_);
  and _80708_ (_29783_, _29782_, _13098_);
  and _80709_ (_29784_, _29783_, _29781_);
  nand _80710_ (_29786_, _06685_, _13107_);
  and _80711_ (_29787_, _29786_, _25414_);
  or _80712_ (_29788_, _29787_, _29784_);
  nand _80713_ (_29789_, _15729_, _05997_);
  and _80714_ (_29790_, _29789_, _13106_);
  and _80715_ (_29791_, _29790_, _29788_);
  and _80716_ (_29792_, _29495_, _13105_);
  or _80717_ (_29793_, _29792_, _29791_);
  or _80718_ (_29794_, _29793_, _01446_);
  or _80719_ (_29795_, _01442_, \oc8051_golden_model_1.PC [13]);
  and _80720_ (_29797_, _29795_, _43634_);
  and _80721_ (_44221_, _29797_, _29794_);
  nor _80722_ (_29798_, _29493_, \oc8051_golden_model_1.PC [14]);
  nor _80723_ (_29799_, _29798_, _12197_);
  or _80724_ (_29800_, _29799_, _13106_);
  or _80725_ (_29801_, _29799_, _13049_);
  nor _80726_ (_29802_, _12828_, _15930_);
  nor _80727_ (_29803_, _12805_, _15930_);
  nor _80728_ (_29804_, _12783_, _15930_);
  nor _80729_ (_29805_, _12724_, _15930_);
  nor _80730_ (_29807_, _12486_, _12384_);
  nor _80731_ (_29808_, _29807_, _12487_);
  or _80732_ (_29809_, _29808_, _29522_);
  or _80733_ (_29810_, _12381_, _12379_);
  and _80734_ (_29811_, _29810_, _06472_);
  and _80735_ (_29812_, _29811_, _29809_);
  and _80736_ (_29813_, _29799_, _12563_);
  nor _80737_ (_29814_, _12549_, _15930_);
  or _80738_ (_29815_, _12510_, _12381_);
  or _80739_ (_29816_, _29808_, _12512_);
  and _80740_ (_29818_, _29816_, _29815_);
  or _80741_ (_29819_, _29818_, _07275_);
  and _80742_ (_29820_, _12539_, _12205_);
  nor _80743_ (_29821_, _12300_, _12208_);
  nor _80744_ (_29822_, _29821_, _12301_);
  and _80745_ (_29823_, _29822_, _12537_);
  or _80746_ (_29824_, _29823_, _29820_);
  or _80747_ (_29825_, _29824_, _08685_);
  not _80748_ (_29826_, _29799_);
  nor _80749_ (_29827_, _29826_, _12520_);
  and _80750_ (_29829_, _12523_, _12205_);
  and _80751_ (_29830_, _12525_, \oc8051_golden_model_1.PC [14]);
  and _80752_ (_29831_, _29830_, _29217_);
  or _80753_ (_29832_, _29831_, _29829_);
  and _80754_ (_29833_, _29832_, _12516_);
  or _80755_ (_29834_, _29833_, _08687_);
  or _80756_ (_29835_, _29834_, _29827_);
  and _80757_ (_29836_, _29835_, _07270_);
  and _80758_ (_29837_, _29836_, _29825_);
  and _80759_ (_29838_, _29799_, _07269_);
  or _80760_ (_29840_, _29838_, _06474_);
  or _80761_ (_29841_, _29840_, _29837_);
  and _80762_ (_29842_, _29841_, _29819_);
  or _80763_ (_29843_, _29842_, _25228_);
  or _80764_ (_29844_, _29799_, _12502_);
  and _80765_ (_29845_, _29844_, _12549_);
  and _80766_ (_29846_, _29845_, _29843_);
  or _80767_ (_29847_, _29846_, _29814_);
  and _80768_ (_29848_, _29847_, _12551_);
  and _80769_ (_29849_, _29799_, _12552_);
  or _80770_ (_29851_, _29849_, _06417_);
  or _80771_ (_29852_, _29851_, _29848_);
  nand _80772_ (_29853_, _15930_, _06417_);
  and _80773_ (_29854_, _29853_, _12561_);
  and _80774_ (_29855_, _29854_, _29852_);
  or _80775_ (_29856_, _29855_, _29813_);
  and _80776_ (_29857_, _29856_, _12567_);
  or _80777_ (_29858_, _12567_, _15930_);
  nand _80778_ (_29859_, _29858_, _12574_);
  or _80779_ (_29860_, _29859_, _29857_);
  and _80780_ (_29862_, _29808_, _14270_);
  and _80781_ (_29863_, _12609_, _12381_);
  or _80782_ (_29864_, _29863_, _12574_);
  or _80783_ (_29865_, _29864_, _29862_);
  and _80784_ (_29866_, _29865_, _06473_);
  and _80785_ (_29867_, _29866_, _29860_);
  or _80786_ (_29868_, _29867_, _06431_);
  or _80787_ (_29869_, _29868_, _29812_);
  and _80788_ (_29870_, _29808_, _12632_);
  and _80789_ (_29871_, _12630_, _12381_);
  or _80790_ (_29873_, _29871_, _06500_);
  or _80791_ (_29874_, _29873_, _29870_);
  and _80792_ (_29875_, _29874_, _12349_);
  and _80793_ (_29876_, _29875_, _29869_);
  or _80794_ (_29877_, _29808_, _12648_);
  or _80795_ (_29878_, _26636_, _12381_);
  and _80796_ (_29879_, _29878_, _06490_);
  and _80797_ (_29880_, _29879_, _29877_);
  or _80798_ (_29881_, _29880_, _12347_);
  or _80799_ (_29882_, _29881_, _29876_);
  or _80800_ (_29884_, _29799_, _12348_);
  and _80801_ (_29885_, _29884_, _12662_);
  and _80802_ (_29886_, _29885_, _29882_);
  nor _80803_ (_29887_, _12662_, _15930_);
  or _80804_ (_29888_, _29887_, _12345_);
  or _80805_ (_29889_, _29888_, _29886_);
  or _80806_ (_29890_, _29799_, _12344_);
  and _80807_ (_29891_, _29890_, _12669_);
  and _80808_ (_29892_, _29891_, _29889_);
  nor _80809_ (_29893_, _12669_, _15930_);
  or _80810_ (_29895_, _29893_, _12671_);
  or _80811_ (_29896_, _29895_, _29892_);
  or _80812_ (_29897_, _29799_, _12339_);
  and _80813_ (_29898_, _29897_, _12336_);
  and _80814_ (_29899_, _29898_, _29896_);
  nor _80815_ (_29900_, _15930_, _12336_);
  or _80816_ (_29901_, _29900_, _06042_);
  or _80817_ (_29902_, _29901_, _29899_);
  or _80818_ (_29903_, _29799_, _06043_);
  and _80819_ (_29904_, _29903_, _12681_);
  and _80820_ (_29906_, _29904_, _29902_);
  nor _80821_ (_29907_, _12681_, _15930_);
  or _80822_ (_29908_, _29907_, _06486_);
  or _80823_ (_29909_, _29908_, _29906_);
  or _80824_ (_29910_, _12381_, _06487_);
  and _80825_ (_29911_, _29910_, _06334_);
  and _80826_ (_29912_, _29911_, _29909_);
  nor _80827_ (_29913_, _15930_, _06334_);
  or _80828_ (_29914_, _29913_, _06037_);
  or _80829_ (_29915_, _29914_, _29912_);
  or _80830_ (_29917_, _12381_, _06313_);
  and _80831_ (_29918_, _29917_, _12694_);
  and _80832_ (_29919_, _29918_, _29915_);
  and _80833_ (_29920_, _29799_, _12700_);
  or _80834_ (_29921_, _29920_, _12698_);
  or _80835_ (_29922_, _29921_, _29919_);
  or _80836_ (_29923_, _12697_, _12205_);
  and _80837_ (_29924_, _29923_, _12705_);
  and _80838_ (_29925_, _29924_, _29922_);
  and _80839_ (_29926_, _29822_, _12704_);
  or _80840_ (_29928_, _29926_, _29925_);
  and _80841_ (_29929_, _29928_, _08626_);
  nor _80842_ (_29930_, _15930_, _08626_);
  or _80843_ (_29931_, _29930_, _06277_);
  or _80844_ (_29932_, _29931_, _29929_);
  or _80845_ (_29933_, _12381_, _06278_);
  and _80846_ (_29934_, _29933_, _11029_);
  and _80847_ (_29935_, _29934_, _29932_);
  and _80848_ (_29936_, _12205_, _11028_);
  or _80849_ (_29937_, _29936_, _12718_);
  or _80850_ (_29939_, _29937_, _29935_);
  nor _80851_ (_29940_, _12755_, \oc8051_golden_model_1.DPH [6]);
  nor _80852_ (_29941_, _29940_, _12756_);
  or _80853_ (_29942_, _29941_, _12719_);
  and _80854_ (_29943_, _29942_, _12724_);
  and _80855_ (_29944_, _29943_, _29939_);
  or _80856_ (_29945_, _29944_, _29805_);
  and _80857_ (_29946_, _29945_, _12764_);
  or _80858_ (_29947_, _29822_, _11389_);
  or _80859_ (_29948_, _12205_, _12770_);
  and _80860_ (_29950_, _29948_, _12763_);
  and _80861_ (_29951_, _29950_, _29947_);
  or _80862_ (_29952_, _29951_, _12768_);
  or _80863_ (_29953_, _29952_, _29946_);
  or _80864_ (_29954_, _29799_, _12333_);
  and _80865_ (_29955_, _29954_, _12330_);
  and _80866_ (_29956_, _29955_, _29953_);
  nor _80867_ (_29957_, _15930_, _12330_);
  or _80868_ (_29958_, _29957_, _06502_);
  or _80869_ (_29959_, _29958_, _29956_);
  or _80870_ (_29961_, _12381_, _07334_);
  and _80871_ (_29962_, _29961_, _12783_);
  and _80872_ (_29963_, _29962_, _29959_);
  or _80873_ (_29964_, _29963_, _29804_);
  and _80874_ (_29965_, _29964_, _12788_);
  or _80875_ (_29966_, _29822_, _12770_);
  or _80876_ (_29967_, _12205_, _11389_);
  and _80877_ (_29968_, _29967_, _12787_);
  and _80878_ (_29969_, _29968_, _29966_);
  or _80879_ (_29970_, _29969_, _12792_);
  or _80880_ (_29972_, _29970_, _29965_);
  or _80881_ (_29973_, _29799_, _12328_);
  and _80882_ (_29974_, _29973_, _12322_);
  and _80883_ (_29975_, _29974_, _29972_);
  nor _80884_ (_29976_, _15930_, _12322_);
  or _80885_ (_29977_, _29976_, _06507_);
  or _80886_ (_29978_, _29977_, _29975_);
  or _80887_ (_29979_, _12381_, _07339_);
  and _80888_ (_29980_, _29979_, _12805_);
  and _80889_ (_29981_, _29980_, _29978_);
  or _80890_ (_29983_, _29981_, _29803_);
  and _80891_ (_29984_, _29983_, _12810_);
  or _80892_ (_29985_, _29822_, \oc8051_golden_model_1.PSW [7]);
  or _80893_ (_29986_, _12205_, _10967_);
  and _80894_ (_29987_, _29986_, _12809_);
  and _80895_ (_29988_, _29987_, _29985_);
  or _80896_ (_29989_, _29988_, _12814_);
  or _80897_ (_29990_, _29989_, _29984_);
  or _80898_ (_29991_, _29799_, _12320_);
  and _80899_ (_29992_, _29991_, _12314_);
  and _80900_ (_29994_, _29992_, _29990_);
  nor _80901_ (_29995_, _15930_, _12314_);
  or _80902_ (_29996_, _29995_, _06509_);
  or _80903_ (_29997_, _29996_, _29994_);
  or _80904_ (_29998_, _12381_, _09107_);
  and _80905_ (_29999_, _29998_, _12828_);
  and _80906_ (_30000_, _29999_, _29997_);
  or _80907_ (_30001_, _30000_, _29802_);
  and _80908_ (_30002_, _30001_, _12832_);
  or _80909_ (_30003_, _29822_, _10967_);
  or _80910_ (_30005_, _12205_, \oc8051_golden_model_1.PSW [7]);
  and _80911_ (_30006_, _30005_, _12310_);
  and _80912_ (_30007_, _30006_, _30003_);
  or _80913_ (_30008_, _30007_, _12839_);
  or _80914_ (_30009_, _30008_, _30002_);
  or _80915_ (_30010_, _29799_, _12837_);
  and _80916_ (_30011_, _30010_, _11187_);
  and _80917_ (_30012_, _30011_, _30009_);
  nor _80918_ (_30013_, _15930_, _11187_);
  or _80919_ (_30014_, _30013_, _11216_);
  or _80920_ (_30016_, _30014_, _30012_);
  or _80921_ (_30017_, _29799_, _11217_);
  and _80922_ (_30018_, _30017_, _14116_);
  and _80923_ (_30019_, _30018_, _30016_);
  nor _80924_ (_30020_, _08209_, _14116_);
  or _80925_ (_30021_, _30020_, _07350_);
  or _80926_ (_30022_, _30021_, _30019_);
  nor _80927_ (_30023_, _12205_, _06016_);
  nor _80928_ (_30024_, _30023_, _06512_);
  and _80929_ (_30025_, _30024_, _30022_);
  or _80930_ (_30027_, _29808_, _13038_);
  or _80931_ (_30028_, _12381_, _13037_);
  and _80932_ (_30029_, _30028_, _06512_);
  and _80933_ (_30030_, _30029_, _30027_);
  or _80934_ (_30031_, _30030_, _12854_);
  or _80935_ (_30032_, _30031_, _30025_);
  or _80936_ (_30033_, _29799_, _12201_);
  and _80937_ (_30034_, _30033_, _13046_);
  and _80938_ (_30035_, _30034_, _30032_);
  nor _80939_ (_30036_, _13046_, _15930_);
  or _80940_ (_30038_, _30036_, _10564_);
  or _80941_ (_30039_, _30038_, _30035_);
  and _80942_ (_30040_, _30039_, _29801_);
  or _80943_ (_30041_, _30040_, _06361_);
  nand _80944_ (_30042_, _08209_, _06361_);
  and _80945_ (_30043_, _30042_, _06021_);
  and _80946_ (_30044_, _30043_, _30041_);
  nor _80947_ (_30045_, _15930_, _06021_);
  or _80948_ (_30046_, _30045_, _06496_);
  or _80949_ (_30047_, _30046_, _30044_);
  or _80950_ (_30049_, _12381_, _13038_);
  or _80951_ (_30050_, _29808_, _13037_);
  and _80952_ (_30051_, _30050_, _30049_);
  or _80953_ (_30052_, _30051_, _07035_);
  and _80954_ (_30053_, _30052_, _30047_);
  or _80955_ (_30054_, _30053_, _13062_);
  or _80956_ (_30055_, _29799_, _09123_);
  and _80957_ (_30056_, _30055_, _30054_);
  or _80958_ (_30057_, _30056_, _06639_);
  nand _80959_ (_30058_, _15930_, _06639_);
  and _80960_ (_30060_, _30058_, _13072_);
  and _80961_ (_30061_, _30060_, _30057_);
  and _80962_ (_30062_, _29799_, _26848_);
  or _80963_ (_30063_, _30062_, _06503_);
  or _80964_ (_30064_, _30063_, _30061_);
  nand _80965_ (_30065_, _06503_, _06397_);
  and _80966_ (_30066_, _30065_, _13082_);
  and _80967_ (_30067_, _30066_, _30064_);
  and _80968_ (_30068_, _12205_, _05998_);
  or _80969_ (_30069_, _30068_, _05989_);
  or _80970_ (_30071_, _30069_, _30067_);
  or _80971_ (_30072_, _30051_, _05990_);
  and _80972_ (_30073_, _30072_, _13087_);
  and _80973_ (_30074_, _30073_, _30071_);
  nor _80974_ (_30075_, _29826_, _13087_);
  or _80975_ (_30076_, _30075_, _06646_);
  or _80976_ (_30077_, _30076_, _30074_);
  nand _80977_ (_30078_, _15930_, _06646_);
  and _80978_ (_30079_, _30078_, _13095_);
  and _80979_ (_30080_, _30079_, _30077_);
  and _80980_ (_30082_, _29799_, _26866_);
  or _80981_ (_30083_, _30082_, _06488_);
  or _80982_ (_30084_, _30083_, _30080_);
  nand _80983_ (_30085_, _06488_, _06397_);
  and _80984_ (_30086_, _30085_, _13107_);
  and _80985_ (_30087_, _30086_, _30084_);
  and _80986_ (_30088_, _12205_, _05997_);
  or _80987_ (_30089_, _30088_, _13105_);
  or _80988_ (_30090_, _30089_, _30087_);
  and _80989_ (_30091_, _30090_, _29800_);
  or _80990_ (_30093_, _30091_, _01446_);
  or _80991_ (_30094_, _01442_, \oc8051_golden_model_1.PC [14]);
  and _80992_ (_30095_, _30094_, _43634_);
  and _80993_ (_44222_, _30095_, _30093_);
  nor _80994_ (_30096_, \oc8051_golden_model_1.P2 [0], rst);
  nor _80995_ (_30097_, _30096_, _00000_);
  and _80996_ (_30098_, _13248_, _08032_);
  and _80997_ (_30099_, _13139_, \oc8051_golden_model_1.P2 [0]);
  and _80998_ (_30100_, _08032_, _09008_);
  or _80999_ (_30101_, _30100_, _30099_);
  nand _81000_ (_30103_, _30101_, _06507_);
  nor _81001_ (_30104_, _30103_, _30098_);
  nand _81002_ (_30105_, _13248_, _06071_);
  or _81003_ (_30106_, _13248_, _06071_);
  and _81004_ (_30107_, _30106_, _30105_);
  and _81005_ (_30108_, _30107_, _08032_);
  or _81006_ (_30109_, _30108_, _30099_);
  and _81007_ (_30110_, _30109_, _06615_);
  or _81008_ (_30111_, _30099_, _30098_);
  or _81009_ (_30112_, _30111_, _07275_);
  and _81010_ (_30114_, _08032_, \oc8051_golden_model_1.ACC [0]);
  or _81011_ (_30115_, _30114_, _30099_);
  and _81012_ (_30116_, _30115_, _07259_);
  and _81013_ (_30117_, _07260_, \oc8051_golden_model_1.P2 [0]);
  or _81014_ (_30118_, _30117_, _06474_);
  or _81015_ (_30119_, _30118_, _30116_);
  and _81016_ (_30120_, _30119_, _06357_);
  and _81017_ (_30121_, _30120_, _30112_);
  not _81018_ (_30122_, _08655_);
  and _81019_ (_30123_, _30122_, \oc8051_golden_model_1.P2 [0]);
  and _81020_ (_30125_, _08657_, \oc8051_golden_model_1.P3 [0]);
  and _81021_ (_30126_, _08661_, \oc8051_golden_model_1.P1 [0]);
  and _81022_ (_30127_, _08655_, \oc8051_golden_model_1.P2 [0]);
  or _81023_ (_30128_, _30127_, _30126_);
  or _81024_ (_30129_, _30128_, _30125_);
  and _81025_ (_30130_, _07993_, \oc8051_golden_model_1.P0 [0]);
  nor _81026_ (_30131_, _30130_, _12947_);
  nand _81027_ (_30132_, _30131_, _12939_);
  nor _81028_ (_30133_, _30132_, _30129_);
  nand _81029_ (_30134_, _30133_, _12946_);
  or _81030_ (_30136_, _30134_, _08451_);
  or _81031_ (_30137_, _30136_, _07967_);
  and _81032_ (_30138_, _30137_, _08655_);
  or _81033_ (_30139_, _30138_, _30123_);
  and _81034_ (_30140_, _30139_, _06356_);
  or _81035_ (_30141_, _30140_, _30121_);
  and _81036_ (_30142_, _30141_, _06772_);
  and _81037_ (_30143_, _08032_, _07250_);
  or _81038_ (_30144_, _30143_, _30099_);
  and _81039_ (_30145_, _30144_, _06410_);
  or _81040_ (_30147_, _30145_, _06417_);
  or _81041_ (_30148_, _30147_, _30142_);
  or _81042_ (_30149_, _30115_, _06426_);
  and _81043_ (_30150_, _30149_, _06353_);
  and _81044_ (_30151_, _30150_, _30148_);
  and _81045_ (_30152_, _30099_, _06352_);
  or _81046_ (_30153_, _30152_, _06345_);
  or _81047_ (_30154_, _30153_, _30151_);
  or _81048_ (_30155_, _30111_, _06346_);
  and _81049_ (_30156_, _30155_, _06340_);
  and _81050_ (_30158_, _30156_, _30154_);
  or _81051_ (_30159_, _30123_, _16663_);
  and _81052_ (_30160_, _30159_, _06339_);
  and _81053_ (_30161_, _30160_, _30139_);
  or _81054_ (_30162_, _30161_, _10153_);
  or _81055_ (_30163_, _30162_, _30158_);
  or _81056_ (_30164_, _30144_, _06327_);
  and _81057_ (_30165_, _30164_, _30163_);
  or _81058_ (_30166_, _30165_, _09572_);
  and _81059_ (_30167_, _09447_, _08032_);
  or _81060_ (_30169_, _30099_, _06333_);
  or _81061_ (_30170_, _30169_, _30167_);
  and _81062_ (_30171_, _30170_, _06313_);
  and _81063_ (_30172_, _30171_, _30166_);
  and _81064_ (_30173_, _08989_, \oc8051_golden_model_1.P2 [0]);
  and _81065_ (_30174_, _08993_, \oc8051_golden_model_1.P0 [0]);
  and _81066_ (_30175_, _08998_, \oc8051_golden_model_1.P1 [0]);
  and _81067_ (_30176_, _09002_, \oc8051_golden_model_1.P3 [0]);
  or _81068_ (_30177_, _30176_, _30175_);
  or _81069_ (_30178_, _30177_, _30174_);
  or _81070_ (_30180_, _30178_, _30173_);
  or _81071_ (_30181_, _30180_, _14645_);
  or _81072_ (_30182_, _30181_, _14662_);
  or _81073_ (_30183_, _30182_, _14644_);
  or _81074_ (_30184_, _30183_, _14637_);
  or _81075_ (_30185_, _30184_, _14624_);
  and _81076_ (_30186_, _30185_, _08032_);
  or _81077_ (_30187_, _30186_, _30099_);
  and _81078_ (_30188_, _30187_, _06037_);
  or _81079_ (_30189_, _30188_, _06277_);
  or _81080_ (_30191_, _30189_, _30172_);
  or _81081_ (_30192_, _30101_, _06278_);
  and _81082_ (_30193_, _30192_, _30191_);
  or _81083_ (_30194_, _30193_, _06502_);
  nor _81084_ (_30195_, _13248_, _06950_);
  not _81085_ (_30196_, _30195_);
  nand _81086_ (_30197_, _13248_, _06950_);
  and _81087_ (_30198_, _30197_, _30196_);
  and _81088_ (_30199_, _30198_, _08032_);
  or _81089_ (_30200_, _30099_, _07334_);
  or _81090_ (_30202_, _30200_, _30199_);
  and _81091_ (_30203_, _30202_, _07337_);
  and _81092_ (_30204_, _30203_, _30194_);
  or _81093_ (_30205_, _30204_, _30110_);
  and _81094_ (_30206_, _30205_, _07339_);
  or _81095_ (_30207_, _30206_, _30104_);
  and _81096_ (_30208_, _30207_, _07331_);
  not _81097_ (_30209_, _13248_);
  or _81098_ (_30210_, _30099_, _30209_);
  and _81099_ (_30211_, _30115_, _06610_);
  and _81100_ (_30213_, _30211_, _30210_);
  or _81101_ (_30214_, _30213_, _06509_);
  or _81102_ (_30215_, _30214_, _30208_);
  and _81103_ (_30216_, _30197_, _08032_);
  or _81104_ (_30217_, _30099_, _09107_);
  or _81105_ (_30218_, _30217_, _30216_);
  and _81106_ (_30219_, _30218_, _09112_);
  and _81107_ (_30220_, _30219_, _30215_);
  and _81108_ (_30221_, _30105_, _08032_);
  or _81109_ (_30222_, _30221_, _30099_);
  and _81110_ (_30224_, _30222_, _06602_);
  or _81111_ (_30225_, _30224_, _06639_);
  or _81112_ (_30226_, _30225_, _30220_);
  or _81113_ (_30227_, _30111_, _07048_);
  and _81114_ (_30228_, _30227_, _05990_);
  and _81115_ (_30229_, _30228_, _30226_);
  and _81116_ (_30230_, _30099_, _05989_);
  or _81117_ (_30231_, _30230_, _06646_);
  or _81118_ (_30232_, _30231_, _30229_);
  or _81119_ (_30233_, _30111_, _06651_);
  and _81120_ (_30235_, _30233_, _01442_);
  and _81121_ (_30236_, _30235_, _30232_);
  or _81122_ (_44223_, _30236_, _30097_);
  nor _81123_ (_30237_, \oc8051_golden_model_1.P2 [1], rst);
  nor _81124_ (_30238_, _30237_, _00000_);
  and _81125_ (_30239_, _13139_, \oc8051_golden_model_1.P2 [1]);
  nor _81126_ (_30240_, _13139_, _07448_);
  or _81127_ (_30241_, _30240_, _30239_);
  or _81128_ (_30242_, _30241_, _06772_);
  or _81129_ (_30243_, _08032_, \oc8051_golden_model_1.P2 [1]);
  nor _81130_ (_30245_, _13363_, _13249_);
  and _81131_ (_30246_, _30245_, _08032_);
  not _81132_ (_30247_, _30246_);
  and _81133_ (_30248_, _30247_, _30243_);
  or _81134_ (_30249_, _30248_, _07275_);
  nand _81135_ (_30250_, _08032_, _06097_);
  and _81136_ (_30251_, _30250_, _30243_);
  and _81137_ (_30252_, _30251_, _07259_);
  and _81138_ (_30253_, _07260_, \oc8051_golden_model_1.P2 [1]);
  or _81139_ (_30254_, _30253_, _06474_);
  or _81140_ (_30256_, _30254_, _30252_);
  and _81141_ (_30257_, _30256_, _06357_);
  and _81142_ (_30258_, _30257_, _30249_);
  and _81143_ (_30259_, _30122_, \oc8051_golden_model_1.P2 [1]);
  and _81144_ (_30260_, _08657_, \oc8051_golden_model_1.P3 [1]);
  nor _81145_ (_30261_, _30260_, _12894_);
  and _81146_ (_30262_, _30261_, _12886_);
  and _81147_ (_30263_, _08661_, \oc8051_golden_model_1.P1 [1]);
  and _81148_ (_30264_, _07993_, \oc8051_golden_model_1.P0 [1]);
  and _81149_ (_30265_, _08655_, \oc8051_golden_model_1.P2 [1]);
  or _81150_ (_30267_, _30265_, _30264_);
  nor _81151_ (_30268_, _30267_, _30263_);
  and _81152_ (_30269_, _30268_, _12893_);
  and _81153_ (_30270_, _30269_, _30262_);
  and _81154_ (_30271_, _30270_, _08402_);
  nand _81155_ (_30272_, _30271_, _12880_);
  and _81156_ (_30273_, _30272_, _08655_);
  or _81157_ (_30274_, _30273_, _30259_);
  and _81158_ (_30275_, _30274_, _06356_);
  or _81159_ (_30276_, _30275_, _06410_);
  or _81160_ (_30277_, _30276_, _30258_);
  and _81161_ (_30278_, _30277_, _30242_);
  or _81162_ (_30279_, _30278_, _06417_);
  or _81163_ (_30280_, _30251_, _06426_);
  and _81164_ (_30281_, _30280_, _06353_);
  and _81165_ (_30282_, _30281_, _30279_);
  nor _81166_ (_30283_, _30271_, _07957_);
  and _81167_ (_30284_, _30283_, _08655_);
  or _81168_ (_30285_, _30284_, _30259_);
  and _81169_ (_30286_, _30285_, _06352_);
  or _81170_ (_30289_, _30286_, _06345_);
  or _81171_ (_30290_, _30289_, _30282_);
  or _81172_ (_30291_, _30271_, _12880_);
  and _81173_ (_30292_, _30273_, _30291_);
  or _81174_ (_30293_, _30259_, _06346_);
  or _81175_ (_30294_, _30293_, _30292_);
  and _81176_ (_30295_, _30294_, _30290_);
  and _81177_ (_30296_, _30295_, _06340_);
  or _81178_ (_30297_, _30283_, _14795_);
  and _81179_ (_30298_, _30297_, _08655_);
  or _81180_ (_30300_, _30259_, _30298_);
  and _81181_ (_30301_, _30300_, _06339_);
  or _81182_ (_30302_, _30301_, _10153_);
  or _81183_ (_30303_, _30302_, _30296_);
  or _81184_ (_30304_, _30241_, _06327_);
  and _81185_ (_30305_, _30304_, _30303_);
  or _81186_ (_30306_, _30305_, _09572_);
  and _81187_ (_30307_, _09402_, _08032_);
  or _81188_ (_30308_, _30239_, _06333_);
  or _81189_ (_30309_, _30308_, _30307_);
  and _81190_ (_30311_, _30309_, _06313_);
  and _81191_ (_30312_, _30311_, _30306_);
  and _81192_ (_30313_, _08993_, \oc8051_golden_model_1.P0 [1]);
  and _81193_ (_30314_, _08989_, \oc8051_golden_model_1.P2 [1]);
  and _81194_ (_30315_, _08998_, \oc8051_golden_model_1.P1 [1]);
  and _81195_ (_30316_, _09002_, \oc8051_golden_model_1.P3 [1]);
  or _81196_ (_30317_, _30316_, _30315_);
  or _81197_ (_30318_, _30317_, _30314_);
  or _81198_ (_30319_, _30318_, _30313_);
  or _81199_ (_30320_, _30319_, _14839_);
  or _81200_ (_30322_, _30320_, _14838_);
  or _81201_ (_30323_, _30322_, _14831_);
  or _81202_ (_30324_, _30323_, _14826_);
  or _81203_ (_30325_, _30324_, _14809_);
  and _81204_ (_30326_, _30325_, _08032_);
  or _81205_ (_30327_, _30326_, _30239_);
  and _81206_ (_30328_, _30327_, _06037_);
  or _81207_ (_30329_, _30328_, _30312_);
  and _81208_ (_30330_, _30329_, _06278_);
  nand _81209_ (_30331_, _08032_, _07160_);
  and _81210_ (_30333_, _30243_, _06277_);
  and _81211_ (_30334_, _30333_, _30331_);
  or _81212_ (_30335_, _30334_, _30330_);
  and _81213_ (_30336_, _30335_, _07334_);
  nor _81214_ (_30337_, _13237_, _07160_);
  and _81215_ (_30338_, _13237_, _07160_);
  nor _81216_ (_30339_, _30338_, _30337_);
  or _81217_ (_30340_, _30339_, _13139_);
  and _81218_ (_30341_, _30243_, _06502_);
  and _81219_ (_30342_, _30341_, _30340_);
  or _81220_ (_30344_, _30342_, _30336_);
  and _81221_ (_30345_, _30344_, _07337_);
  nand _81222_ (_30346_, _13237_, _06097_);
  or _81223_ (_30347_, _13237_, _06097_);
  and _81224_ (_30348_, _30347_, _30346_);
  or _81225_ (_30349_, _30348_, _13139_);
  and _81226_ (_30350_, _30243_, _06615_);
  and _81227_ (_30351_, _30350_, _30349_);
  or _81228_ (_30352_, _30351_, _30345_);
  and _81229_ (_30353_, _30352_, _07339_);
  or _81230_ (_30355_, _30337_, _13139_);
  and _81231_ (_30356_, _30243_, _06507_);
  and _81232_ (_30357_, _30356_, _30355_);
  or _81233_ (_30358_, _30357_, _30353_);
  and _81234_ (_30359_, _30358_, _07331_);
  not _81235_ (_30360_, _13237_);
  or _81236_ (_30361_, _30239_, _30360_);
  and _81237_ (_30362_, _30251_, _06610_);
  and _81238_ (_30363_, _30362_, _30361_);
  or _81239_ (_30364_, _30363_, _30359_);
  and _81240_ (_30366_, _30364_, _06603_);
  or _81241_ (_30367_, _30250_, _30360_);
  and _81242_ (_30368_, _30243_, _06602_);
  and _81243_ (_30369_, _30368_, _30367_);
  or _81244_ (_30370_, _30369_, _06639_);
  or _81245_ (_30371_, _30331_, _30360_);
  and _81246_ (_30372_, _30243_, _06509_);
  and _81247_ (_30373_, _30372_, _30371_);
  or _81248_ (_30374_, _30373_, _30370_);
  or _81249_ (_30375_, _30374_, _30366_);
  or _81250_ (_30377_, _30248_, _07048_);
  and _81251_ (_30378_, _30377_, _05990_);
  and _81252_ (_30379_, _30378_, _30375_);
  and _81253_ (_30380_, _30285_, _05989_);
  or _81254_ (_30381_, _30380_, _06646_);
  or _81255_ (_30382_, _30381_, _30379_);
  or _81256_ (_30383_, _30239_, _06651_);
  or _81257_ (_30384_, _30383_, _30246_);
  and _81258_ (_30385_, _30384_, _01442_);
  and _81259_ (_30386_, _30385_, _30382_);
  or _81260_ (_44225_, _30386_, _30238_);
  nor _81261_ (_30388_, \oc8051_golden_model_1.P2 [2], rst);
  nor _81262_ (_30389_, _30388_, _00000_);
  and _81263_ (_30390_, _13139_, \oc8051_golden_model_1.P2 [2]);
  nand _81264_ (_30391_, _13219_, _10280_);
  or _81265_ (_30392_, _13219_, _10280_);
  and _81266_ (_30393_, _30392_, _30391_);
  and _81267_ (_30394_, _30393_, _08032_);
  or _81268_ (_30395_, _30394_, _30390_);
  and _81269_ (_30396_, _30395_, _06615_);
  nor _81270_ (_30398_, _13139_, _07854_);
  or _81271_ (_30399_, _30398_, _30390_);
  or _81272_ (_30400_, _30399_, _06327_);
  or _81273_ (_30401_, _30399_, _06772_);
  nor _81274_ (_30402_, _13249_, _13219_);
  or _81275_ (_30403_, _30402_, _13250_);
  and _81276_ (_30404_, _30403_, _08032_);
  or _81277_ (_30405_, _30404_, _30390_);
  or _81278_ (_30406_, _30405_, _07275_);
  and _81279_ (_30407_, _08032_, \oc8051_golden_model_1.ACC [2]);
  or _81280_ (_30409_, _30407_, _30390_);
  and _81281_ (_30410_, _30409_, _07259_);
  and _81282_ (_30411_, _07260_, \oc8051_golden_model_1.P2 [2]);
  or _81283_ (_30412_, _30411_, _06474_);
  or _81284_ (_30413_, _30412_, _30410_);
  and _81285_ (_30414_, _30413_, _06357_);
  and _81286_ (_30415_, _30414_, _30406_);
  and _81287_ (_30416_, _30122_, \oc8051_golden_model_1.P2 [2]);
  and _81288_ (_30417_, _07993_, \oc8051_golden_model_1.P0 [2]);
  and _81289_ (_30418_, _08655_, \oc8051_golden_model_1.P2 [2]);
  nor _81290_ (_30420_, _30418_, _30417_);
  and _81291_ (_30421_, _08661_, \oc8051_golden_model_1.P1 [2]);
  and _81292_ (_30422_, _08657_, \oc8051_golden_model_1.P3 [2]);
  nor _81293_ (_30423_, _30422_, _30421_);
  and _81294_ (_30424_, _30423_, _30420_);
  and _81295_ (_30425_, _30424_, _12868_);
  and _81296_ (_30426_, _30425_, _12865_);
  and _81297_ (_30427_, _30426_, _08501_);
  nand _81298_ (_30428_, _30427_, _12855_);
  and _81299_ (_30429_, _30428_, _08655_);
  or _81300_ (_30431_, _30429_, _30416_);
  and _81301_ (_30432_, _30431_, _06356_);
  or _81302_ (_30433_, _30432_, _06410_);
  or _81303_ (_30434_, _30433_, _30415_);
  and _81304_ (_30435_, _30434_, _30401_);
  or _81305_ (_30436_, _30435_, _06417_);
  or _81306_ (_30437_, _30409_, _06426_);
  and _81307_ (_30438_, _30437_, _06353_);
  and _81308_ (_30439_, _30438_, _30436_);
  nor _81309_ (_30440_, _30427_, _08000_);
  and _81310_ (_30442_, _30440_, _08655_);
  or _81311_ (_30443_, _30442_, _30416_);
  and _81312_ (_30444_, _30443_, _06352_);
  or _81313_ (_30445_, _30444_, _06345_);
  or _81314_ (_30446_, _30445_, _30439_);
  or _81315_ (_30447_, _30427_, _12855_);
  and _81316_ (_30448_, _30429_, _30447_);
  or _81317_ (_30449_, _30416_, _06346_);
  or _81318_ (_30450_, _30449_, _30448_);
  and _81319_ (_30451_, _30450_, _06340_);
  and _81320_ (_30453_, _30451_, _30446_);
  or _81321_ (_30454_, _30440_, _14999_);
  and _81322_ (_30455_, _30454_, _08655_);
  or _81323_ (_30456_, _30455_, _30416_);
  and _81324_ (_30457_, _30456_, _06339_);
  or _81325_ (_30458_, _30457_, _10153_);
  or _81326_ (_30459_, _30458_, _30453_);
  and _81327_ (_30460_, _30459_, _30400_);
  or _81328_ (_30461_, _30460_, _09572_);
  and _81329_ (_30462_, _09356_, _08032_);
  or _81330_ (_30464_, _30390_, _06333_);
  or _81331_ (_30465_, _30464_, _30462_);
  and _81332_ (_30466_, _30465_, _06313_);
  and _81333_ (_30467_, _30466_, _30461_);
  and _81334_ (_30468_, _08989_, \oc8051_golden_model_1.P2 [2]);
  and _81335_ (_30469_, _08993_, \oc8051_golden_model_1.P0 [2]);
  and _81336_ (_30470_, _08998_, \oc8051_golden_model_1.P1 [2]);
  and _81337_ (_30471_, _09002_, \oc8051_golden_model_1.P3 [2]);
  or _81338_ (_30472_, _30471_, _30470_);
  or _81339_ (_30473_, _30472_, _30469_);
  or _81340_ (_30475_, _30473_, _30468_);
  or _81341_ (_30476_, _30475_, _15024_);
  or _81342_ (_30477_, _30476_, _15038_);
  or _81343_ (_30478_, _30477_, _15054_);
  or _81344_ (_30479_, _30478_, _15014_);
  and _81345_ (_30480_, _30479_, _08032_);
  or _81346_ (_30481_, _30480_, _30390_);
  and _81347_ (_30482_, _30481_, _06037_);
  or _81348_ (_30483_, _30482_, _06277_);
  or _81349_ (_30484_, _30483_, _30467_);
  and _81350_ (_30486_, _08032_, _09057_);
  or _81351_ (_30487_, _30486_, _30390_);
  or _81352_ (_30488_, _30487_, _06278_);
  and _81353_ (_30489_, _30488_, _30484_);
  or _81354_ (_30490_, _30489_, _06502_);
  nand _81355_ (_30491_, _13219_, _06769_);
  or _81356_ (_30492_, _13219_, _06769_);
  and _81357_ (_30493_, _30492_, _30491_);
  and _81358_ (_30494_, _30493_, _08032_);
  or _81359_ (_30495_, _30390_, _07334_);
  or _81360_ (_30497_, _30495_, _30494_);
  and _81361_ (_30498_, _30497_, _07337_);
  and _81362_ (_30499_, _30498_, _30490_);
  or _81363_ (_30500_, _30499_, _30396_);
  and _81364_ (_30501_, _30500_, _07339_);
  or _81365_ (_30502_, _30390_, _13362_);
  and _81366_ (_30503_, _30487_, _06507_);
  and _81367_ (_30504_, _30503_, _30502_);
  or _81368_ (_30505_, _30504_, _30501_);
  and _81369_ (_30506_, _30505_, _07331_);
  and _81370_ (_30508_, _30409_, _06610_);
  and _81371_ (_30509_, _30508_, _30502_);
  or _81372_ (_30510_, _30509_, _06509_);
  or _81373_ (_30511_, _30510_, _30506_);
  and _81374_ (_30512_, _30491_, _08032_);
  or _81375_ (_30513_, _30390_, _09107_);
  or _81376_ (_30514_, _30513_, _30512_);
  and _81377_ (_30515_, _30514_, _09112_);
  and _81378_ (_30516_, _30515_, _30511_);
  and _81379_ (_30517_, _30391_, _08032_);
  or _81380_ (_30519_, _30517_, _30390_);
  and _81381_ (_30520_, _30519_, _06602_);
  or _81382_ (_30521_, _30520_, _06639_);
  or _81383_ (_30522_, _30521_, _30516_);
  or _81384_ (_30523_, _30405_, _07048_);
  and _81385_ (_30524_, _30523_, _05990_);
  and _81386_ (_30525_, _30524_, _30522_);
  and _81387_ (_30526_, _30443_, _05989_);
  or _81388_ (_30527_, _30526_, _06646_);
  or _81389_ (_30528_, _30527_, _30525_);
  nor _81390_ (_30530_, _13363_, _13362_);
  nor _81391_ (_30531_, _30530_, _13364_);
  and _81392_ (_30532_, _30531_, _08032_);
  or _81393_ (_30533_, _30390_, _06651_);
  or _81394_ (_30534_, _30533_, _30532_);
  and _81395_ (_30535_, _30534_, _01442_);
  and _81396_ (_30536_, _30535_, _30528_);
  or _81397_ (_44226_, _30536_, _30389_);
  nor _81398_ (_30537_, \oc8051_golden_model_1.P2 [3], rst);
  nor _81399_ (_30538_, _30537_, _00000_);
  and _81400_ (_30540_, _13139_, \oc8051_golden_model_1.P2 [3]);
  nand _81401_ (_30541_, _13208_, _10334_);
  or _81402_ (_30542_, _13208_, _10334_);
  and _81403_ (_30543_, _30542_, _30541_);
  and _81404_ (_30544_, _30543_, _08032_);
  or _81405_ (_30545_, _30544_, _30540_);
  and _81406_ (_30546_, _30545_, _06615_);
  nor _81407_ (_30547_, _13139_, _07680_);
  or _81408_ (_30548_, _30547_, _30540_);
  or _81409_ (_30549_, _30548_, _06327_);
  nor _81410_ (_30551_, _13250_, _13208_);
  or _81411_ (_30552_, _30551_, _13251_);
  and _81412_ (_30553_, _30552_, _08032_);
  or _81413_ (_30554_, _30553_, _30540_);
  or _81414_ (_30555_, _30554_, _07275_);
  and _81415_ (_30556_, _08032_, \oc8051_golden_model_1.ACC [3]);
  or _81416_ (_30557_, _30556_, _30540_);
  and _81417_ (_30558_, _30557_, _07259_);
  and _81418_ (_30559_, _07260_, \oc8051_golden_model_1.P2 [3]);
  or _81419_ (_30560_, _30559_, _06474_);
  or _81420_ (_30562_, _30560_, _30558_);
  and _81421_ (_30563_, _30562_, _06357_);
  and _81422_ (_30564_, _30563_, _30555_);
  and _81423_ (_30565_, _30122_, \oc8051_golden_model_1.P2 [3]);
  and _81424_ (_30566_, _08661_, \oc8051_golden_model_1.P1 [3]);
  and _81425_ (_30567_, _08657_, \oc8051_golden_model_1.P3 [3]);
  nor _81426_ (_30568_, _30567_, _30566_);
  and _81427_ (_30569_, _07993_, \oc8051_golden_model_1.P0 [3]);
  and _81428_ (_30570_, _08655_, \oc8051_golden_model_1.P2 [3]);
  nor _81429_ (_30571_, _30570_, _30569_);
  and _81430_ (_30573_, _30571_, _30568_);
  and _81431_ (_30574_, _30573_, _12997_);
  and _81432_ (_30575_, _30574_, _12994_);
  and _81433_ (_30576_, _30575_, _08357_);
  nand _81434_ (_30577_, _30576_, _12984_);
  and _81435_ (_30578_, _30577_, _08655_);
  or _81436_ (_30579_, _30578_, _30565_);
  and _81437_ (_30580_, _30579_, _06356_);
  or _81438_ (_30581_, _30580_, _06410_);
  or _81439_ (_30582_, _30581_, _30564_);
  or _81440_ (_30584_, _30548_, _06772_);
  and _81441_ (_30585_, _30584_, _30582_);
  or _81442_ (_30586_, _30585_, _06417_);
  or _81443_ (_30587_, _30557_, _06426_);
  and _81444_ (_30588_, _30587_, _06353_);
  and _81445_ (_30589_, _30588_, _30586_);
  nor _81446_ (_30590_, _30576_, _07994_);
  and _81447_ (_30591_, _30590_, _08655_);
  or _81448_ (_30592_, _30591_, _30565_);
  and _81449_ (_30593_, _30592_, _06352_);
  or _81450_ (_30595_, _30593_, _06345_);
  or _81451_ (_30596_, _30595_, _30589_);
  or _81452_ (_30597_, _30576_, _12984_);
  or _81453_ (_30598_, _30565_, _30597_);
  and _81454_ (_30599_, _30598_, _30579_);
  or _81455_ (_30600_, _30599_, _06346_);
  and _81456_ (_30601_, _30600_, _06340_);
  and _81457_ (_30602_, _30601_, _30596_);
  or _81458_ (_30603_, _30590_, _15196_);
  and _81459_ (_30604_, _30603_, _08655_);
  or _81460_ (_30606_, _30604_, _30565_);
  and _81461_ (_30607_, _30606_, _06339_);
  or _81462_ (_30608_, _30607_, _10153_);
  or _81463_ (_30609_, _30608_, _30602_);
  and _81464_ (_30610_, _30609_, _30549_);
  or _81465_ (_30611_, _30610_, _09572_);
  and _81466_ (_30612_, _09310_, _08032_);
  or _81467_ (_30613_, _30540_, _06333_);
  or _81468_ (_30614_, _30613_, _30612_);
  and _81469_ (_30615_, _30614_, _06313_);
  and _81470_ (_30617_, _30615_, _30611_);
  and _81471_ (_30618_, _08993_, \oc8051_golden_model_1.P0 [3]);
  and _81472_ (_30619_, _08989_, \oc8051_golden_model_1.P2 [3]);
  and _81473_ (_30620_, _08998_, \oc8051_golden_model_1.P1 [3]);
  and _81474_ (_30621_, _09002_, \oc8051_golden_model_1.P3 [3]);
  or _81475_ (_30622_, _30621_, _30620_);
  or _81476_ (_30623_, _30622_, _30619_);
  or _81477_ (_30624_, _30623_, _30618_);
  or _81478_ (_30625_, _30624_, _15219_);
  or _81479_ (_30626_, _30625_, _15233_);
  or _81480_ (_30628_, _30626_, _15249_);
  or _81481_ (_30629_, _30628_, _15209_);
  and _81482_ (_30630_, _30629_, _08032_);
  or _81483_ (_30631_, _30630_, _30540_);
  and _81484_ (_30632_, _30631_, _06037_);
  or _81485_ (_30633_, _30632_, _06277_);
  or _81486_ (_30634_, _30633_, _30617_);
  and _81487_ (_30635_, _08032_, _09014_);
  or _81488_ (_30636_, _30635_, _30540_);
  or _81489_ (_30637_, _30636_, _06278_);
  and _81490_ (_30639_, _30637_, _30634_);
  or _81491_ (_30640_, _30639_, _06502_);
  nand _81492_ (_30641_, _13208_, _06595_);
  or _81493_ (_30642_, _13208_, _06595_);
  and _81494_ (_30643_, _30642_, _30641_);
  and _81495_ (_30644_, _30643_, _08032_);
  or _81496_ (_30645_, _30540_, _07334_);
  or _81497_ (_30646_, _30645_, _30644_);
  and _81498_ (_30647_, _30646_, _07337_);
  and _81499_ (_30648_, _30647_, _30640_);
  or _81500_ (_30650_, _30648_, _30546_);
  and _81501_ (_30651_, _30650_, _07339_);
  or _81502_ (_30652_, _30540_, _13361_);
  and _81503_ (_30653_, _30636_, _06507_);
  and _81504_ (_30654_, _30653_, _30652_);
  or _81505_ (_30655_, _30654_, _30651_);
  and _81506_ (_30656_, _30655_, _07331_);
  and _81507_ (_30657_, _30557_, _06610_);
  and _81508_ (_30658_, _30657_, _30652_);
  or _81509_ (_30659_, _30658_, _06509_);
  or _81510_ (_30661_, _30659_, _30656_);
  and _81511_ (_30662_, _30641_, _08032_);
  or _81512_ (_30663_, _30540_, _09107_);
  or _81513_ (_30664_, _30663_, _30662_);
  and _81514_ (_30665_, _30664_, _09112_);
  and _81515_ (_30666_, _30665_, _30661_);
  and _81516_ (_30667_, _30541_, _08032_);
  or _81517_ (_30668_, _30667_, _30540_);
  and _81518_ (_30669_, _30668_, _06602_);
  or _81519_ (_30670_, _30669_, _06639_);
  or _81520_ (_30672_, _30670_, _30666_);
  or _81521_ (_30673_, _30554_, _07048_);
  and _81522_ (_30674_, _30673_, _05990_);
  and _81523_ (_30675_, _30674_, _30672_);
  and _81524_ (_30676_, _30592_, _05989_);
  or _81525_ (_30677_, _30676_, _06646_);
  or _81526_ (_30678_, _30677_, _30675_);
  nor _81527_ (_30679_, _13364_, _13361_);
  nor _81528_ (_30680_, _30679_, _13365_);
  and _81529_ (_30681_, _30680_, _08032_);
  or _81530_ (_30683_, _30540_, _06651_);
  or _81531_ (_30684_, _30683_, _30681_);
  and _81532_ (_30685_, _30684_, _01442_);
  and _81533_ (_30686_, _30685_, _30678_);
  or _81534_ (_44227_, _30686_, _30538_);
  nor _81535_ (_30687_, \oc8051_golden_model_1.P2 [4], rst);
  nor _81536_ (_30688_, _30687_, _00000_);
  and _81537_ (_30689_, _13139_, \oc8051_golden_model_1.P2 [4]);
  nand _81538_ (_30690_, _13197_, _10204_);
  or _81539_ (_30691_, _13197_, _10204_);
  and _81540_ (_30693_, _30691_, _30690_);
  and _81541_ (_30694_, _30693_, _08032_);
  or _81542_ (_30695_, _30694_, _30689_);
  and _81543_ (_30696_, _30695_, _06615_);
  nor _81544_ (_30697_, _08596_, _13139_);
  or _81545_ (_30698_, _30697_, _30689_);
  or _81546_ (_30699_, _30698_, _06327_);
  and _81547_ (_30700_, _30122_, \oc8051_golden_model_1.P2 [4]);
  and _81548_ (_30701_, _07993_, \oc8051_golden_model_1.P0 [4]);
  and _81549_ (_30702_, _08655_, \oc8051_golden_model_1.P2 [4]);
  nor _81550_ (_30704_, _30702_, _30701_);
  and _81551_ (_30705_, _08661_, \oc8051_golden_model_1.P1 [4]);
  and _81552_ (_30706_, _08657_, \oc8051_golden_model_1.P3 [4]);
  nor _81553_ (_30707_, _30706_, _30705_);
  and _81554_ (_30708_, _30707_, _30704_);
  and _81555_ (_30709_, _30708_, _12917_);
  and _81556_ (_30710_, _30709_, _12914_);
  and _81557_ (_30711_, _30710_, _08597_);
  nor _81558_ (_30712_, _30711_, _12928_);
  and _81559_ (_30713_, _30712_, _08655_);
  or _81560_ (_30715_, _30713_, _30700_);
  and _81561_ (_30716_, _30715_, _06352_);
  nor _81562_ (_30717_, _13251_, _13197_);
  or _81563_ (_30718_, _30717_, _13252_);
  and _81564_ (_30719_, _30718_, _08032_);
  or _81565_ (_30720_, _30719_, _30689_);
  or _81566_ (_30721_, _30720_, _07275_);
  and _81567_ (_30722_, _08032_, \oc8051_golden_model_1.ACC [4]);
  or _81568_ (_30723_, _30722_, _30689_);
  and _81569_ (_30724_, _30723_, _07259_);
  and _81570_ (_30726_, _07260_, \oc8051_golden_model_1.P2 [4]);
  or _81571_ (_30727_, _30726_, _06474_);
  or _81572_ (_30728_, _30727_, _30724_);
  and _81573_ (_30729_, _30728_, _06357_);
  and _81574_ (_30730_, _30729_, _30721_);
  nand _81575_ (_30731_, _30711_, _12929_);
  and _81576_ (_30732_, _30731_, _08655_);
  or _81577_ (_30733_, _30732_, _30700_);
  and _81578_ (_30734_, _30733_, _06356_);
  or _81579_ (_30735_, _30734_, _06410_);
  or _81580_ (_30737_, _30735_, _30730_);
  or _81581_ (_30738_, _30698_, _06772_);
  and _81582_ (_30739_, _30738_, _30737_);
  or _81583_ (_30740_, _30739_, _06417_);
  or _81584_ (_30741_, _30723_, _06426_);
  and _81585_ (_30742_, _30741_, _06353_);
  and _81586_ (_30743_, _30742_, _30740_);
  or _81587_ (_30744_, _30743_, _30716_);
  and _81588_ (_30745_, _30744_, _06346_);
  or _81589_ (_30746_, _30711_, _12929_);
  or _81590_ (_30748_, _30700_, _30746_);
  and _81591_ (_30749_, _30733_, _06345_);
  and _81592_ (_30750_, _30749_, _30748_);
  or _81593_ (_30751_, _30750_, _30745_);
  and _81594_ (_30752_, _30751_, _06340_);
  or _81595_ (_30753_, _30712_, _15349_);
  and _81596_ (_30754_, _30753_, _08655_);
  or _81597_ (_30755_, _30754_, _30700_);
  and _81598_ (_30756_, _30755_, _06339_);
  or _81599_ (_30757_, _30756_, _10153_);
  or _81600_ (_30759_, _30757_, _30752_);
  and _81601_ (_30760_, _30759_, _30699_);
  or _81602_ (_30761_, _30760_, _09572_);
  and _81603_ (_30762_, _09264_, _08032_);
  or _81604_ (_30763_, _30689_, _06333_);
  or _81605_ (_30764_, _30763_, _30762_);
  and _81606_ (_30765_, _30764_, _06313_);
  and _81607_ (_30766_, _30765_, _30761_);
  and _81608_ (_30767_, _08993_, \oc8051_golden_model_1.P0 [4]);
  and _81609_ (_30768_, _08989_, \oc8051_golden_model_1.P2 [4]);
  and _81610_ (_30770_, _08998_, \oc8051_golden_model_1.P1 [4]);
  and _81611_ (_30771_, _09002_, \oc8051_golden_model_1.P3 [4]);
  or _81612_ (_30772_, _30771_, _30770_);
  or _81613_ (_30773_, _30772_, _30768_);
  or _81614_ (_30774_, _30773_, _30767_);
  or _81615_ (_30775_, _30774_, _15420_);
  or _81616_ (_30776_, _30775_, _15434_);
  or _81617_ (_30777_, _30776_, _15450_);
  or _81618_ (_30778_, _30777_, _15410_);
  and _81619_ (_30779_, _30778_, _08032_);
  or _81620_ (_30781_, _30779_, _30689_);
  and _81621_ (_30782_, _30781_, _06037_);
  or _81622_ (_30783_, _30782_, _06277_);
  or _81623_ (_30784_, _30783_, _30766_);
  and _81624_ (_30785_, _08995_, _08032_);
  or _81625_ (_30786_, _30785_, _30689_);
  or _81626_ (_30787_, _30786_, _06278_);
  and _81627_ (_30788_, _30787_, _30784_);
  or _81628_ (_30789_, _30788_, _06502_);
  nand _81629_ (_30790_, _13197_, _08986_);
  or _81630_ (_30792_, _13197_, _08986_);
  and _81631_ (_30793_, _30792_, _30790_);
  and _81632_ (_30794_, _30793_, _08032_);
  or _81633_ (_30795_, _30689_, _07334_);
  or _81634_ (_30796_, _30795_, _30794_);
  and _81635_ (_30797_, _30796_, _07337_);
  and _81636_ (_30798_, _30797_, _30789_);
  or _81637_ (_30799_, _30798_, _30696_);
  and _81638_ (_30800_, _30799_, _07339_);
  or _81639_ (_30801_, _30689_, _13360_);
  and _81640_ (_30803_, _30786_, _06507_);
  and _81641_ (_30804_, _30803_, _30801_);
  or _81642_ (_30805_, _30804_, _30800_);
  and _81643_ (_30806_, _30805_, _07331_);
  and _81644_ (_30807_, _30723_, _06610_);
  and _81645_ (_30808_, _30807_, _30801_);
  or _81646_ (_30809_, _30808_, _06509_);
  or _81647_ (_30810_, _30809_, _30806_);
  and _81648_ (_30811_, _30790_, _08032_);
  or _81649_ (_30812_, _30689_, _09107_);
  or _81650_ (_30814_, _30812_, _30811_);
  and _81651_ (_30815_, _30814_, _09112_);
  and _81652_ (_30816_, _30815_, _30810_);
  and _81653_ (_30817_, _30690_, _08032_);
  or _81654_ (_30818_, _30817_, _30689_);
  and _81655_ (_30819_, _30818_, _06602_);
  or _81656_ (_30820_, _30819_, _06639_);
  or _81657_ (_30821_, _30820_, _30816_);
  or _81658_ (_30822_, _30720_, _07048_);
  and _81659_ (_30823_, _30822_, _05990_);
  and _81660_ (_30825_, _30823_, _30821_);
  and _81661_ (_30826_, _30715_, _05989_);
  or _81662_ (_30827_, _30826_, _06646_);
  or _81663_ (_30828_, _30827_, _30825_);
  nor _81664_ (_30829_, _13365_, _13360_);
  nor _81665_ (_30830_, _30829_, _13366_);
  and _81666_ (_30831_, _30830_, _08032_);
  or _81667_ (_30832_, _30689_, _06651_);
  or _81668_ (_30833_, _30832_, _30831_);
  and _81669_ (_30834_, _30833_, _01442_);
  and _81670_ (_30836_, _30834_, _30828_);
  or _81671_ (_44228_, _30836_, _30688_);
  nor _81672_ (_30837_, \oc8051_golden_model_1.P2 [5], rst);
  nor _81673_ (_30838_, _30837_, _00000_);
  and _81674_ (_30839_, _13139_, \oc8051_golden_model_1.P2 [5]);
  nand _81675_ (_30840_, _13186_, _10237_);
  or _81676_ (_30841_, _13186_, _10237_);
  and _81677_ (_30842_, _30841_, _30840_);
  and _81678_ (_30843_, _30842_, _08032_);
  or _81679_ (_30844_, _30843_, _30839_);
  and _81680_ (_30846_, _30844_, _06615_);
  nor _81681_ (_30847_, _13252_, _13186_);
  or _81682_ (_30848_, _30847_, _13253_);
  and _81683_ (_30849_, _30848_, _08032_);
  or _81684_ (_30850_, _30849_, _30839_);
  or _81685_ (_30851_, _30850_, _07275_);
  and _81686_ (_30852_, _08032_, \oc8051_golden_model_1.ACC [5]);
  or _81687_ (_30853_, _30852_, _30839_);
  and _81688_ (_30854_, _30853_, _07259_);
  and _81689_ (_30855_, _07260_, \oc8051_golden_model_1.P2 [5]);
  or _81690_ (_30857_, _30855_, _06474_);
  or _81691_ (_30858_, _30857_, _30854_);
  and _81692_ (_30859_, _30858_, _06357_);
  and _81693_ (_30860_, _30859_, _30851_);
  and _81694_ (_30861_, _30122_, \oc8051_golden_model_1.P2 [5]);
  and _81695_ (_30862_, _07993_, \oc8051_golden_model_1.P0 [5]);
  and _81696_ (_30863_, _08655_, \oc8051_golden_model_1.P2 [5]);
  nor _81697_ (_30864_, _30863_, _30862_);
  and _81698_ (_30865_, _08661_, \oc8051_golden_model_1.P1 [5]);
  and _81699_ (_30866_, _08657_, \oc8051_golden_model_1.P3 [5]);
  nor _81700_ (_30868_, _30866_, _30865_);
  and _81701_ (_30869_, _30868_, _30864_);
  and _81702_ (_30870_, _30869_, _13021_);
  and _81703_ (_30871_, _30870_, _13018_);
  and _81704_ (_30872_, _30871_, _08306_);
  nand _81705_ (_30873_, _30872_, _13033_);
  and _81706_ (_30874_, _30873_, _08655_);
  or _81707_ (_30875_, _30874_, _30861_);
  and _81708_ (_30876_, _30875_, _06356_);
  or _81709_ (_30877_, _30876_, _06410_);
  or _81710_ (_30879_, _30877_, _30860_);
  nor _81711_ (_30880_, _08305_, _13139_);
  or _81712_ (_30881_, _30880_, _30839_);
  or _81713_ (_30882_, _30881_, _06772_);
  and _81714_ (_30883_, _30882_, _30879_);
  or _81715_ (_30884_, _30883_, _06417_);
  or _81716_ (_30885_, _30853_, _06426_);
  and _81717_ (_30886_, _30885_, _06353_);
  and _81718_ (_30887_, _30886_, _30884_);
  nor _81719_ (_30888_, _30872_, _13032_);
  and _81720_ (_30890_, _30888_, _08655_);
  or _81721_ (_30891_, _30890_, _30861_);
  and _81722_ (_30892_, _30891_, _06352_);
  or _81723_ (_30893_, _30892_, _06345_);
  or _81724_ (_30894_, _30893_, _30887_);
  or _81725_ (_30895_, _30872_, _13033_);
  or _81726_ (_30896_, _30861_, _30895_);
  and _81727_ (_30897_, _30896_, _30875_);
  or _81728_ (_30898_, _30897_, _06346_);
  and _81729_ (_30899_, _30898_, _06340_);
  and _81730_ (_30901_, _30899_, _30894_);
  or _81731_ (_30902_, _30888_, _15545_);
  and _81732_ (_30903_, _30902_, _08655_);
  or _81733_ (_30904_, _30903_, _30861_);
  and _81734_ (_30905_, _30904_, _06339_);
  or _81735_ (_30906_, _30905_, _10153_);
  or _81736_ (_30907_, _30906_, _30901_);
  or _81737_ (_30908_, _30881_, _06327_);
  and _81738_ (_30909_, _30908_, _30907_);
  or _81739_ (_30910_, _30909_, _09572_);
  and _81740_ (_30912_, _09218_, _08032_);
  or _81741_ (_30913_, _30839_, _06333_);
  or _81742_ (_30914_, _30913_, _30912_);
  and _81743_ (_30915_, _30914_, _06313_);
  and _81744_ (_30916_, _30915_, _30910_);
  and _81745_ (_30917_, _08989_, \oc8051_golden_model_1.P2 [5]);
  and _81746_ (_30918_, _08993_, \oc8051_golden_model_1.P0 [5]);
  and _81747_ (_30919_, _08998_, \oc8051_golden_model_1.P1 [5]);
  and _81748_ (_30920_, _09002_, \oc8051_golden_model_1.P3 [5]);
  or _81749_ (_30921_, _30920_, _30919_);
  or _81750_ (_30923_, _30921_, _30918_);
  or _81751_ (_30924_, _30923_, _30917_);
  or _81752_ (_30925_, _30924_, _15617_);
  or _81753_ (_30926_, _30925_, _15631_);
  or _81754_ (_30927_, _30926_, _15647_);
  or _81755_ (_30928_, _30927_, _15607_);
  and _81756_ (_30929_, _30928_, _08032_);
  or _81757_ (_30930_, _30929_, _30839_);
  and _81758_ (_30931_, _30930_, _06037_);
  or _81759_ (_30932_, _30931_, _06277_);
  or _81760_ (_30934_, _30932_, _30916_);
  and _81761_ (_30935_, _08954_, _08032_);
  or _81762_ (_30936_, _30935_, _30839_);
  or _81763_ (_30937_, _30936_, _06278_);
  and _81764_ (_30938_, _30937_, _30934_);
  or _81765_ (_30939_, _30938_, _06502_);
  nand _81766_ (_30940_, _13186_, _08953_);
  or _81767_ (_30941_, _13186_, _08953_);
  and _81768_ (_30942_, _30941_, _30940_);
  and _81769_ (_30943_, _30942_, _08032_);
  or _81770_ (_30945_, _30839_, _07334_);
  or _81771_ (_30946_, _30945_, _30943_);
  and _81772_ (_30947_, _30946_, _07337_);
  and _81773_ (_30948_, _30947_, _30939_);
  or _81774_ (_30949_, _30948_, _30846_);
  and _81775_ (_30950_, _30949_, _07339_);
  or _81776_ (_30951_, _30839_, _13359_);
  and _81777_ (_30952_, _30936_, _06507_);
  and _81778_ (_30953_, _30952_, _30951_);
  or _81779_ (_30954_, _30953_, _30950_);
  and _81780_ (_30956_, _30954_, _07331_);
  and _81781_ (_30957_, _30853_, _06610_);
  and _81782_ (_30958_, _30957_, _30951_);
  or _81783_ (_30959_, _30958_, _06509_);
  or _81784_ (_30960_, _30959_, _30956_);
  and _81785_ (_30961_, _30940_, _08032_);
  or _81786_ (_30962_, _30839_, _09107_);
  or _81787_ (_30963_, _30962_, _30961_);
  and _81788_ (_30964_, _30963_, _09112_);
  and _81789_ (_30965_, _30964_, _30960_);
  and _81790_ (_30967_, _30840_, _08032_);
  or _81791_ (_30968_, _30967_, _30839_);
  and _81792_ (_30969_, _30968_, _06602_);
  or _81793_ (_30970_, _30969_, _06639_);
  or _81794_ (_30971_, _30970_, _30965_);
  or _81795_ (_30972_, _30850_, _07048_);
  and _81796_ (_30973_, _30972_, _05990_);
  and _81797_ (_30974_, _30973_, _30971_);
  and _81798_ (_30975_, _30891_, _05989_);
  or _81799_ (_30976_, _30975_, _06646_);
  or _81800_ (_30978_, _30976_, _30974_);
  nor _81801_ (_30979_, _13366_, _13359_);
  nor _81802_ (_30980_, _30979_, _13367_);
  and _81803_ (_30981_, _30980_, _08032_);
  or _81804_ (_30982_, _30839_, _06651_);
  or _81805_ (_30983_, _30982_, _30981_);
  and _81806_ (_30984_, _30983_, _01442_);
  and _81807_ (_30985_, _30984_, _30978_);
  or _81808_ (_44229_, _30985_, _30838_);
  nor _81809_ (_30986_, \oc8051_golden_model_1.P2 [6], rst);
  nor _81810_ (_30988_, _30986_, _00000_);
  and _81811_ (_30989_, _13139_, \oc8051_golden_model_1.P2 [6]);
  nand _81812_ (_30990_, _13175_, _10193_);
  or _81813_ (_30991_, _13175_, _10193_);
  and _81814_ (_30992_, _30991_, _30990_);
  and _81815_ (_30993_, _30992_, _08032_);
  or _81816_ (_30994_, _30993_, _30989_);
  and _81817_ (_30995_, _30994_, _06615_);
  nor _81818_ (_30996_, _08209_, _13139_);
  or _81819_ (_30997_, _30996_, _30989_);
  or _81820_ (_31000_, _30997_, _06327_);
  and _81821_ (_31001_, _30122_, \oc8051_golden_model_1.P2 [6]);
  and _81822_ (_31002_, _07993_, \oc8051_golden_model_1.P0 [6]);
  and _81823_ (_31003_, _08655_, \oc8051_golden_model_1.P2 [6]);
  nor _81824_ (_31004_, _31003_, _31002_);
  and _81825_ (_31005_, _08661_, \oc8051_golden_model_1.P1 [6]);
  and _81826_ (_31006_, _08657_, \oc8051_golden_model_1.P3 [6]);
  nor _81827_ (_31007_, _31006_, _31005_);
  and _81828_ (_31008_, _31007_, _31004_);
  and _81829_ (_31009_, _31008_, _12969_);
  and _81830_ (_31011_, _31009_, _12966_);
  and _81831_ (_31012_, _31011_, _08210_);
  nor _81832_ (_31013_, _31012_, _12980_);
  and _81833_ (_31014_, _31013_, _08655_);
  or _81834_ (_31015_, _31014_, _31001_);
  and _81835_ (_31016_, _31015_, _06352_);
  nor _81836_ (_31017_, _13253_, _13175_);
  or _81837_ (_31018_, _31017_, _13254_);
  and _81838_ (_31019_, _31018_, _08032_);
  or _81839_ (_31020_, _31019_, _30989_);
  or _81840_ (_31023_, _31020_, _07275_);
  and _81841_ (_31024_, _08032_, \oc8051_golden_model_1.ACC [6]);
  or _81842_ (_31025_, _31024_, _30989_);
  and _81843_ (_31026_, _31025_, _07259_);
  and _81844_ (_31027_, _07260_, \oc8051_golden_model_1.P2 [6]);
  or _81845_ (_31028_, _31027_, _06474_);
  or _81846_ (_31029_, _31028_, _31026_);
  and _81847_ (_31030_, _31029_, _06357_);
  and _81848_ (_31031_, _31030_, _31023_);
  nand _81849_ (_31032_, _31012_, _12981_);
  and _81850_ (_31034_, _31032_, _08655_);
  or _81851_ (_31035_, _31034_, _31001_);
  and _81852_ (_31036_, _31035_, _06356_);
  or _81853_ (_31037_, _31036_, _06410_);
  or _81854_ (_31038_, _31037_, _31031_);
  or _81855_ (_31039_, _30997_, _06772_);
  and _81856_ (_31040_, _31039_, _31038_);
  or _81857_ (_31041_, _31040_, _06417_);
  or _81858_ (_31042_, _31025_, _06426_);
  and _81859_ (_31043_, _31042_, _06353_);
  and _81860_ (_31046_, _31043_, _31041_);
  or _81861_ (_31047_, _31046_, _31016_);
  and _81862_ (_31048_, _31047_, _06346_);
  or _81863_ (_31049_, _31012_, _12981_);
  or _81864_ (_31050_, _31001_, _31049_);
  and _81865_ (_31051_, _31035_, _06345_);
  and _81866_ (_31052_, _31051_, _31050_);
  or _81867_ (_31053_, _31052_, _31048_);
  and _81868_ (_31054_, _31053_, _06340_);
  or _81869_ (_31055_, _31013_, _15744_);
  and _81870_ (_31057_, _31055_, _08655_);
  or _81871_ (_31058_, _31057_, _31001_);
  and _81872_ (_31059_, _31058_, _06339_);
  or _81873_ (_31060_, _31059_, _10153_);
  or _81874_ (_31061_, _31060_, _31054_);
  and _81875_ (_31062_, _31061_, _31000_);
  or _81876_ (_31063_, _31062_, _09572_);
  and _81877_ (_31064_, _09172_, _08032_);
  or _81878_ (_31065_, _30989_, _06333_);
  or _81879_ (_31066_, _31065_, _31064_);
  and _81880_ (_31069_, _31066_, _06313_);
  and _81881_ (_31070_, _31069_, _31063_);
  and _81882_ (_31071_, _08993_, \oc8051_golden_model_1.P0 [6]);
  and _81883_ (_31072_, _08989_, \oc8051_golden_model_1.P2 [6]);
  and _81884_ (_31073_, _08998_, \oc8051_golden_model_1.P1 [6]);
  and _81885_ (_31074_, _09002_, \oc8051_golden_model_1.P3 [6]);
  or _81886_ (_31075_, _31074_, _31073_);
  or _81887_ (_31076_, _31075_, _31072_);
  or _81888_ (_31077_, _31076_, _31071_);
  or _81889_ (_31078_, _31077_, _15814_);
  or _81890_ (_31080_, _31078_, _15828_);
  or _81891_ (_31081_, _31080_, _15844_);
  or _81892_ (_31082_, _31081_, _15804_);
  and _81893_ (_31083_, _31082_, _08032_);
  or _81894_ (_31084_, _31083_, _30989_);
  and _81895_ (_31085_, _31084_, _06037_);
  or _81896_ (_31086_, _31085_, _06277_);
  or _81897_ (_31087_, _31086_, _31070_);
  and _81898_ (_31088_, _15853_, _08032_);
  or _81899_ (_31089_, _31088_, _30989_);
  or _81900_ (_31091_, _31089_, _06278_);
  and _81901_ (_31092_, _31091_, _31087_);
  or _81902_ (_31093_, _31092_, _06502_);
  nand _81903_ (_31094_, _13175_, _08918_);
  or _81904_ (_31095_, _13175_, _08918_);
  and _81905_ (_31096_, _31095_, _31094_);
  and _81906_ (_31097_, _31096_, _08032_);
  or _81907_ (_31098_, _30989_, _07334_);
  or _81908_ (_31099_, _31098_, _31097_);
  and _81909_ (_31100_, _31099_, _07337_);
  and _81910_ (_31102_, _31100_, _31093_);
  or _81911_ (_31103_, _31102_, _30995_);
  and _81912_ (_31104_, _31103_, _07339_);
  or _81913_ (_31105_, _30989_, _13358_);
  and _81914_ (_31106_, _31089_, _06507_);
  and _81915_ (_31107_, _31106_, _31105_);
  or _81916_ (_31108_, _31107_, _31104_);
  and _81917_ (_31109_, _31108_, _07331_);
  and _81918_ (_31110_, _31025_, _06610_);
  and _81919_ (_31111_, _31110_, _31105_);
  or _81920_ (_31113_, _31111_, _06509_);
  or _81921_ (_31114_, _31113_, _31109_);
  and _81922_ (_31115_, _31094_, _08032_);
  or _81923_ (_31116_, _30989_, _09107_);
  or _81924_ (_31117_, _31116_, _31115_);
  and _81925_ (_31118_, _31117_, _09112_);
  and _81926_ (_31119_, _31118_, _31114_);
  and _81927_ (_31120_, _30990_, _08032_);
  or _81928_ (_31121_, _31120_, _30989_);
  and _81929_ (_31122_, _31121_, _06602_);
  or _81930_ (_31124_, _31122_, _06639_);
  or _81931_ (_31125_, _31124_, _31119_);
  or _81932_ (_31126_, _31020_, _07048_);
  and _81933_ (_31127_, _31126_, _05990_);
  and _81934_ (_31128_, _31127_, _31125_);
  and _81935_ (_31129_, _31015_, _05989_);
  or _81936_ (_31130_, _31129_, _06646_);
  or _81937_ (_31131_, _31130_, _31128_);
  nor _81938_ (_31132_, _13367_, _13358_);
  nor _81939_ (_31133_, _31132_, _13368_);
  and _81940_ (_31135_, _31133_, _08032_);
  or _81941_ (_31136_, _30989_, _06651_);
  or _81942_ (_31137_, _31136_, _31135_);
  and _81943_ (_31138_, _31137_, _01442_);
  and _81944_ (_31139_, _31138_, _31131_);
  or _81945_ (_44230_, _31139_, _30988_);
  nor _81946_ (_31140_, \oc8051_golden_model_1.P3 [0], rst);
  nor _81947_ (_31141_, _31140_, _00000_);
  and _81948_ (_31142_, _13248_, _08034_);
  and _81949_ (_31143_, _13379_, \oc8051_golden_model_1.P3 [0]);
  and _81950_ (_31145_, _08034_, _09008_);
  or _81951_ (_31146_, _31145_, _31143_);
  nand _81952_ (_31147_, _31146_, _06507_);
  nor _81953_ (_31148_, _31147_, _31142_);
  and _81954_ (_31149_, _30107_, _08034_);
  or _81955_ (_31150_, _31149_, _31143_);
  and _81956_ (_31151_, _31150_, _06615_);
  or _81957_ (_31152_, _31143_, _31142_);
  or _81958_ (_31153_, _31152_, _07275_);
  and _81959_ (_31154_, _08034_, \oc8051_golden_model_1.ACC [0]);
  or _81960_ (_31156_, _31154_, _31143_);
  and _81961_ (_31157_, _31156_, _07259_);
  and _81962_ (_31158_, _07260_, \oc8051_golden_model_1.P3 [0]);
  or _81963_ (_31159_, _31158_, _06474_);
  or _81964_ (_31160_, _31159_, _31157_);
  and _81965_ (_31161_, _31160_, _06357_);
  and _81966_ (_31162_, _31161_, _31153_);
  and _81967_ (_31163_, _13387_, \oc8051_golden_model_1.P3 [0]);
  and _81968_ (_31164_, _30137_, _08657_);
  or _81969_ (_31165_, _31164_, _31163_);
  and _81970_ (_31167_, _31165_, _06356_);
  or _81971_ (_31168_, _31167_, _31162_);
  and _81972_ (_31169_, _31168_, _06772_);
  and _81973_ (_31170_, _08034_, _07250_);
  or _81974_ (_31171_, _31170_, _31143_);
  and _81975_ (_31172_, _31171_, _06410_);
  or _81976_ (_31173_, _31172_, _06417_);
  or _81977_ (_31174_, _31173_, _31169_);
  or _81978_ (_31175_, _31156_, _06426_);
  and _81979_ (_31176_, _31175_, _06353_);
  and _81980_ (_31178_, _31176_, _31174_);
  and _81981_ (_31179_, _31143_, _06352_);
  or _81982_ (_31180_, _31179_, _06345_);
  or _81983_ (_31181_, _31180_, _31178_);
  or _81984_ (_31182_, _31152_, _06346_);
  and _81985_ (_31183_, _31182_, _06340_);
  and _81986_ (_31184_, _31183_, _31181_);
  or _81987_ (_31185_, _31163_, _16663_);
  and _81988_ (_31186_, _31185_, _06339_);
  and _81989_ (_31187_, _31186_, _31165_);
  or _81990_ (_31189_, _31187_, _10153_);
  or _81991_ (_31190_, _31189_, _31184_);
  or _81992_ (_31191_, _31171_, _06327_);
  and _81993_ (_31192_, _31191_, _31190_);
  or _81994_ (_31193_, _31192_, _09572_);
  and _81995_ (_31194_, _09447_, _08034_);
  or _81996_ (_31195_, _31143_, _06333_);
  or _81997_ (_31196_, _31195_, _31194_);
  and _81998_ (_31197_, _31196_, _06313_);
  and _81999_ (_31198_, _31197_, _31193_);
  and _82000_ (_31200_, _30185_, _08034_);
  or _82001_ (_31201_, _31200_, _31143_);
  and _82002_ (_31202_, _31201_, _06037_);
  or _82003_ (_31203_, _31202_, _06277_);
  or _82004_ (_31204_, _31203_, _31198_);
  or _82005_ (_31205_, _31146_, _06278_);
  and _82006_ (_31206_, _31205_, _31204_);
  or _82007_ (_31207_, _31206_, _06502_);
  and _82008_ (_31208_, _30198_, _08034_);
  or _82009_ (_31209_, _31143_, _07334_);
  or _82010_ (_31211_, _31209_, _31208_);
  and _82011_ (_31212_, _31211_, _07337_);
  and _82012_ (_31213_, _31212_, _31207_);
  or _82013_ (_31214_, _31213_, _31151_);
  and _82014_ (_31215_, _31214_, _07339_);
  or _82015_ (_31216_, _31215_, _31148_);
  and _82016_ (_31217_, _31216_, _07331_);
  or _82017_ (_31218_, _31143_, _30209_);
  and _82018_ (_31219_, _31156_, _06610_);
  and _82019_ (_31220_, _31219_, _31218_);
  or _82020_ (_31222_, _31220_, _06509_);
  or _82021_ (_31223_, _31222_, _31217_);
  and _82022_ (_31224_, _30197_, _08034_);
  or _82023_ (_31225_, _31143_, _09107_);
  or _82024_ (_31226_, _31225_, _31224_);
  and _82025_ (_31227_, _31226_, _09112_);
  and _82026_ (_31228_, _31227_, _31223_);
  and _82027_ (_31229_, _30105_, _08034_);
  or _82028_ (_31230_, _31229_, _31143_);
  and _82029_ (_31231_, _31230_, _06602_);
  or _82030_ (_31233_, _31231_, _06639_);
  or _82031_ (_31234_, _31233_, _31228_);
  or _82032_ (_31235_, _31152_, _07048_);
  and _82033_ (_31236_, _31235_, _05990_);
  and _82034_ (_31237_, _31236_, _31234_);
  and _82035_ (_31238_, _31143_, _05989_);
  or _82036_ (_31239_, _31238_, _06646_);
  or _82037_ (_31240_, _31239_, _31237_);
  or _82038_ (_31241_, _31152_, _06651_);
  and _82039_ (_31242_, _31241_, _01442_);
  and _82040_ (_31244_, _31242_, _31240_);
  or _82041_ (_44232_, _31244_, _31141_);
  nor _82042_ (_31245_, \oc8051_golden_model_1.P3 [1], rst);
  nor _82043_ (_31246_, _31245_, _00000_);
  nand _82044_ (_31247_, _08034_, _07160_);
  or _82045_ (_31248_, _08034_, \oc8051_golden_model_1.P3 [1]);
  and _82046_ (_31249_, _31248_, _06277_);
  and _82047_ (_31250_, _31249_, _31247_);
  and _82048_ (_31251_, _13379_, \oc8051_golden_model_1.P3 [1]);
  nor _82049_ (_31252_, _13379_, _07448_);
  or _82050_ (_31254_, _31252_, _31251_);
  or _82051_ (_31255_, _31254_, _06772_);
  and _82052_ (_31256_, _30245_, _08034_);
  not _82053_ (_31257_, _31256_);
  and _82054_ (_31258_, _31257_, _31248_);
  or _82055_ (_31259_, _31258_, _07275_);
  nand _82056_ (_31260_, _08034_, _06097_);
  and _82057_ (_31261_, _31260_, _31248_);
  and _82058_ (_31262_, _31261_, _07259_);
  and _82059_ (_31263_, _07260_, \oc8051_golden_model_1.P3 [1]);
  or _82060_ (_31265_, _31263_, _06474_);
  or _82061_ (_31266_, _31265_, _31262_);
  and _82062_ (_31267_, _31266_, _06357_);
  and _82063_ (_31268_, _31267_, _31259_);
  and _82064_ (_31269_, _13387_, \oc8051_golden_model_1.P3 [1]);
  and _82065_ (_31270_, _30272_, _08657_);
  or _82066_ (_31271_, _31270_, _31269_);
  and _82067_ (_31272_, _31271_, _06356_);
  or _82068_ (_31273_, _31272_, _06410_);
  or _82069_ (_31274_, _31273_, _31268_);
  and _82070_ (_31276_, _31274_, _31255_);
  or _82071_ (_31277_, _31276_, _06417_);
  or _82072_ (_31278_, _31261_, _06426_);
  and _82073_ (_31279_, _31278_, _06353_);
  and _82074_ (_31280_, _31279_, _31277_);
  and _82075_ (_31281_, _30283_, _08657_);
  or _82076_ (_31282_, _31281_, _31269_);
  and _82077_ (_31283_, _31282_, _06352_);
  or _82078_ (_31284_, _31283_, _06345_);
  or _82079_ (_31285_, _31284_, _31280_);
  and _82080_ (_31287_, _31270_, _30291_);
  or _82081_ (_31288_, _31269_, _06346_);
  or _82082_ (_31289_, _31288_, _31287_);
  and _82083_ (_31290_, _31289_, _31285_);
  and _82084_ (_31291_, _31290_, _06340_);
  and _82085_ (_31292_, _30297_, _08657_);
  or _82086_ (_31293_, _31269_, _31292_);
  and _82087_ (_31294_, _31293_, _06339_);
  or _82088_ (_31295_, _31294_, _10153_);
  or _82089_ (_31296_, _31295_, _31291_);
  or _82090_ (_31298_, _31254_, _06327_);
  and _82091_ (_31299_, _31298_, _31296_);
  or _82092_ (_31300_, _31299_, _09572_);
  and _82093_ (_31301_, _09402_, _08034_);
  or _82094_ (_31302_, _31251_, _06333_);
  or _82095_ (_31303_, _31302_, _31301_);
  and _82096_ (_31304_, _31303_, _06313_);
  and _82097_ (_31305_, _31304_, _31300_);
  and _82098_ (_31306_, _30325_, _08034_);
  or _82099_ (_31307_, _31306_, _31251_);
  and _82100_ (_31309_, _31307_, _06037_);
  or _82101_ (_31310_, _31309_, _31305_);
  and _82102_ (_31311_, _31310_, _06278_);
  or _82103_ (_31312_, _31311_, _31250_);
  and _82104_ (_31313_, _31312_, _07334_);
  or _82105_ (_31314_, _30339_, _13379_);
  and _82106_ (_31315_, _31248_, _06502_);
  and _82107_ (_31316_, _31315_, _31314_);
  or _82108_ (_31317_, _31316_, _31313_);
  and _82109_ (_31318_, _31317_, _07337_);
  or _82110_ (_31320_, _30348_, _13379_);
  and _82111_ (_31321_, _31248_, _06615_);
  and _82112_ (_31322_, _31321_, _31320_);
  or _82113_ (_31323_, _31322_, _31318_);
  and _82114_ (_31324_, _31323_, _07339_);
  or _82115_ (_31325_, _30337_, _13379_);
  and _82116_ (_31326_, _31248_, _06507_);
  and _82117_ (_31327_, _31326_, _31325_);
  or _82118_ (_31328_, _31327_, _31324_);
  and _82119_ (_31329_, _31328_, _07331_);
  or _82120_ (_31331_, _31251_, _30360_);
  and _82121_ (_31332_, _31261_, _06610_);
  and _82122_ (_31333_, _31332_, _31331_);
  or _82123_ (_31334_, _31333_, _31329_);
  and _82124_ (_31335_, _31334_, _06603_);
  or _82125_ (_31336_, _31260_, _30360_);
  and _82126_ (_31337_, _31248_, _06602_);
  and _82127_ (_31338_, _31337_, _31336_);
  or _82128_ (_31339_, _31338_, _06639_);
  or _82129_ (_31340_, _31247_, _30360_);
  and _82130_ (_31342_, _31248_, _06509_);
  and _82131_ (_31343_, _31342_, _31340_);
  or _82132_ (_31344_, _31343_, _31339_);
  or _82133_ (_31345_, _31344_, _31335_);
  or _82134_ (_31346_, _31258_, _07048_);
  and _82135_ (_31347_, _31346_, _05990_);
  and _82136_ (_31348_, _31347_, _31345_);
  and _82137_ (_31349_, _31282_, _05989_);
  or _82138_ (_31350_, _31349_, _06646_);
  or _82139_ (_31351_, _31350_, _31348_);
  or _82140_ (_31353_, _31251_, _06651_);
  or _82141_ (_31354_, _31353_, _31256_);
  and _82142_ (_31355_, _31354_, _01442_);
  and _82143_ (_31356_, _31355_, _31351_);
  or _82144_ (_44233_, _31356_, _31246_);
  nor _82145_ (_31357_, \oc8051_golden_model_1.P3 [2], rst);
  nor _82146_ (_31358_, _31357_, _00000_);
  and _82147_ (_31359_, _13379_, \oc8051_golden_model_1.P3 [2]);
  and _82148_ (_31360_, _30393_, _08034_);
  or _82149_ (_31361_, _31360_, _31359_);
  and _82150_ (_31363_, _31361_, _06615_);
  nor _82151_ (_31364_, _13379_, _07854_);
  or _82152_ (_31365_, _31364_, _31359_);
  or _82153_ (_31366_, _31365_, _06327_);
  or _82154_ (_31367_, _31365_, _06772_);
  and _82155_ (_31368_, _30403_, _08034_);
  or _82156_ (_31369_, _31368_, _31359_);
  or _82157_ (_31370_, _31369_, _07275_);
  and _82158_ (_31371_, _08034_, \oc8051_golden_model_1.ACC [2]);
  or _82159_ (_31372_, _31371_, _31359_);
  and _82160_ (_31374_, _31372_, _07259_);
  and _82161_ (_31375_, _07260_, \oc8051_golden_model_1.P3 [2]);
  or _82162_ (_31376_, _31375_, _06474_);
  or _82163_ (_31377_, _31376_, _31374_);
  and _82164_ (_31378_, _31377_, _06357_);
  and _82165_ (_31379_, _31378_, _31370_);
  and _82166_ (_31380_, _13387_, \oc8051_golden_model_1.P3 [2]);
  and _82167_ (_31381_, _30428_, _08657_);
  or _82168_ (_31382_, _31381_, _31380_);
  and _82169_ (_31383_, _31382_, _06356_);
  or _82170_ (_31385_, _31383_, _06410_);
  or _82171_ (_31386_, _31385_, _31379_);
  and _82172_ (_31387_, _31386_, _31367_);
  or _82173_ (_31388_, _31387_, _06417_);
  or _82174_ (_31389_, _31372_, _06426_);
  and _82175_ (_31390_, _31389_, _06353_);
  and _82176_ (_31391_, _31390_, _31388_);
  and _82177_ (_31392_, _30440_, _08657_);
  or _82178_ (_31393_, _31392_, _31380_);
  and _82179_ (_31394_, _31393_, _06352_);
  or _82180_ (_31396_, _31394_, _06345_);
  or _82181_ (_31397_, _31396_, _31391_);
  and _82182_ (_31398_, _31381_, _30447_);
  or _82183_ (_31399_, _31380_, _06346_);
  or _82184_ (_31400_, _31399_, _31398_);
  and _82185_ (_31401_, _31400_, _06340_);
  and _82186_ (_31402_, _31401_, _31397_);
  and _82187_ (_31403_, _30454_, _08657_);
  or _82188_ (_31404_, _31403_, _31380_);
  and _82189_ (_31405_, _31404_, _06339_);
  or _82190_ (_31407_, _31405_, _10153_);
  or _82191_ (_31408_, _31407_, _31402_);
  and _82192_ (_31409_, _31408_, _31366_);
  or _82193_ (_31410_, _31409_, _09572_);
  and _82194_ (_31411_, _09356_, _08034_);
  or _82195_ (_31412_, _31359_, _06333_);
  or _82196_ (_31413_, _31412_, _31411_);
  and _82197_ (_31414_, _31413_, _06313_);
  and _82198_ (_31415_, _31414_, _31410_);
  and _82199_ (_31416_, _30479_, _08034_);
  or _82200_ (_31418_, _31416_, _31359_);
  and _82201_ (_31419_, _31418_, _06037_);
  or _82202_ (_31420_, _31419_, _06277_);
  or _82203_ (_31421_, _31420_, _31415_);
  and _82204_ (_31422_, _08034_, _09057_);
  or _82205_ (_31423_, _31422_, _31359_);
  or _82206_ (_31424_, _31423_, _06278_);
  and _82207_ (_31425_, _31424_, _31421_);
  or _82208_ (_31426_, _31425_, _06502_);
  and _82209_ (_31427_, _30493_, _08034_);
  or _82210_ (_31429_, _31359_, _07334_);
  or _82211_ (_31430_, _31429_, _31427_);
  and _82212_ (_31431_, _31430_, _07337_);
  and _82213_ (_31432_, _31431_, _31426_);
  or _82214_ (_31433_, _31432_, _31363_);
  and _82215_ (_31434_, _31433_, _07339_);
  or _82216_ (_31435_, _31359_, _13362_);
  and _82217_ (_31436_, _31423_, _06507_);
  and _82218_ (_31437_, _31436_, _31435_);
  or _82219_ (_31438_, _31437_, _31434_);
  and _82220_ (_31440_, _31438_, _07331_);
  and _82221_ (_31441_, _31372_, _06610_);
  and _82222_ (_31442_, _31441_, _31435_);
  or _82223_ (_31443_, _31442_, _06509_);
  or _82224_ (_31444_, _31443_, _31440_);
  and _82225_ (_31445_, _30491_, _08034_);
  or _82226_ (_31446_, _31359_, _09107_);
  or _82227_ (_31447_, _31446_, _31445_);
  and _82228_ (_31448_, _31447_, _09112_);
  and _82229_ (_31449_, _31448_, _31444_);
  and _82230_ (_31451_, _30391_, _08034_);
  or _82231_ (_31452_, _31451_, _31359_);
  and _82232_ (_31453_, _31452_, _06602_);
  or _82233_ (_31454_, _31453_, _06639_);
  or _82234_ (_31455_, _31454_, _31449_);
  or _82235_ (_31456_, _31369_, _07048_);
  and _82236_ (_31457_, _31456_, _05990_);
  and _82237_ (_31458_, _31457_, _31455_);
  and _82238_ (_31459_, _31393_, _05989_);
  or _82239_ (_31460_, _31459_, _06646_);
  or _82240_ (_31462_, _31460_, _31458_);
  and _82241_ (_31463_, _30531_, _08034_);
  or _82242_ (_31464_, _31359_, _06651_);
  or _82243_ (_31465_, _31464_, _31463_);
  and _82244_ (_31466_, _31465_, _01442_);
  and _82245_ (_31467_, _31466_, _31462_);
  or _82246_ (_44234_, _31467_, _31358_);
  nor _82247_ (_31468_, \oc8051_golden_model_1.P3 [3], rst);
  nor _82248_ (_31469_, _31468_, _00000_);
  and _82249_ (_31470_, _13379_, \oc8051_golden_model_1.P3 [3]);
  and _82250_ (_31472_, _30543_, _08034_);
  or _82251_ (_31473_, _31472_, _31470_);
  and _82252_ (_31474_, _31473_, _06615_);
  nor _82253_ (_31475_, _13379_, _07680_);
  or _82254_ (_31476_, _31475_, _31470_);
  or _82255_ (_31477_, _31476_, _06327_);
  and _82256_ (_31478_, _30552_, _08034_);
  or _82257_ (_31479_, _31478_, _31470_);
  or _82258_ (_31480_, _31479_, _07275_);
  and _82259_ (_31481_, _08034_, \oc8051_golden_model_1.ACC [3]);
  or _82260_ (_31483_, _31481_, _31470_);
  and _82261_ (_31484_, _31483_, _07259_);
  and _82262_ (_31485_, _07260_, \oc8051_golden_model_1.P3 [3]);
  or _82263_ (_31486_, _31485_, _06474_);
  or _82264_ (_31487_, _31486_, _31484_);
  and _82265_ (_31488_, _31487_, _06357_);
  and _82266_ (_31489_, _31488_, _31480_);
  and _82267_ (_31490_, _13387_, \oc8051_golden_model_1.P3 [3]);
  and _82268_ (_31491_, _30577_, _08657_);
  or _82269_ (_31492_, _31491_, _31490_);
  and _82270_ (_31494_, _31492_, _06356_);
  or _82271_ (_31495_, _31494_, _06410_);
  or _82272_ (_31496_, _31495_, _31489_);
  or _82273_ (_31497_, _31476_, _06772_);
  and _82274_ (_31498_, _31497_, _31496_);
  or _82275_ (_31499_, _31498_, _06417_);
  or _82276_ (_31500_, _31483_, _06426_);
  and _82277_ (_31501_, _31500_, _06353_);
  and _82278_ (_31502_, _31501_, _31499_);
  and _82279_ (_31503_, _30590_, _08657_);
  or _82280_ (_31505_, _31503_, _31490_);
  and _82281_ (_31506_, _31505_, _06352_);
  or _82282_ (_31507_, _31506_, _06345_);
  or _82283_ (_31508_, _31507_, _31502_);
  or _82284_ (_31509_, _31490_, _30597_);
  and _82285_ (_31510_, _31509_, _31492_);
  or _82286_ (_31511_, _31510_, _06346_);
  and _82287_ (_31512_, _31511_, _06340_);
  and _82288_ (_31513_, _31512_, _31508_);
  and _82289_ (_31514_, _30603_, _08657_);
  or _82290_ (_31516_, _31514_, _31490_);
  and _82291_ (_31517_, _31516_, _06339_);
  or _82292_ (_31518_, _31517_, _10153_);
  or _82293_ (_31519_, _31518_, _31513_);
  and _82294_ (_31520_, _31519_, _31477_);
  or _82295_ (_31521_, _31520_, _09572_);
  and _82296_ (_31522_, _09310_, _08034_);
  or _82297_ (_31523_, _31470_, _06333_);
  or _82298_ (_31524_, _31523_, _31522_);
  and _82299_ (_31525_, _31524_, _06313_);
  and _82300_ (_31527_, _31525_, _31521_);
  and _82301_ (_31528_, _30629_, _08034_);
  or _82302_ (_31529_, _31528_, _31470_);
  and _82303_ (_31530_, _31529_, _06037_);
  or _82304_ (_31531_, _31530_, _06277_);
  or _82305_ (_31532_, _31531_, _31527_);
  and _82306_ (_31533_, _08034_, _09014_);
  or _82307_ (_31534_, _31533_, _31470_);
  or _82308_ (_31535_, _31534_, _06278_);
  and _82309_ (_31536_, _31535_, _31532_);
  or _82310_ (_31538_, _31536_, _06502_);
  and _82311_ (_31539_, _30643_, _08034_);
  or _82312_ (_31540_, _31470_, _07334_);
  or _82313_ (_31541_, _31540_, _31539_);
  and _82314_ (_31542_, _31541_, _07337_);
  and _82315_ (_31543_, _31542_, _31538_);
  or _82316_ (_31544_, _31543_, _31474_);
  and _82317_ (_31545_, _31544_, _07339_);
  or _82318_ (_31546_, _31470_, _13361_);
  and _82319_ (_31547_, _31534_, _06507_);
  and _82320_ (_31549_, _31547_, _31546_);
  or _82321_ (_31550_, _31549_, _31545_);
  and _82322_ (_31551_, _31550_, _07331_);
  and _82323_ (_31552_, _31483_, _06610_);
  and _82324_ (_31553_, _31552_, _31546_);
  or _82325_ (_31554_, _31553_, _06509_);
  or _82326_ (_31555_, _31554_, _31551_);
  and _82327_ (_31556_, _30641_, _08034_);
  or _82328_ (_31557_, _31470_, _09107_);
  or _82329_ (_31558_, _31557_, _31556_);
  and _82330_ (_31560_, _31558_, _09112_);
  and _82331_ (_31561_, _31560_, _31555_);
  and _82332_ (_31562_, _30541_, _08034_);
  or _82333_ (_31563_, _31562_, _31470_);
  and _82334_ (_31564_, _31563_, _06602_);
  or _82335_ (_31565_, _31564_, _06639_);
  or _82336_ (_31566_, _31565_, _31561_);
  or _82337_ (_31567_, _31479_, _07048_);
  and _82338_ (_31568_, _31567_, _05990_);
  and _82339_ (_31569_, _31568_, _31566_);
  and _82340_ (_31571_, _31505_, _05989_);
  or _82341_ (_31572_, _31571_, _06646_);
  or _82342_ (_31573_, _31572_, _31569_);
  and _82343_ (_31574_, _30680_, _08034_);
  or _82344_ (_31575_, _31470_, _06651_);
  or _82345_ (_31576_, _31575_, _31574_);
  and _82346_ (_31577_, _31576_, _01442_);
  and _82347_ (_31578_, _31577_, _31573_);
  or _82348_ (_44235_, _31578_, _31469_);
  nor _82349_ (_31579_, \oc8051_golden_model_1.P3 [4], rst);
  nor _82350_ (_31581_, _31579_, _00000_);
  and _82351_ (_31582_, _13379_, \oc8051_golden_model_1.P3 [4]);
  and _82352_ (_31583_, _30693_, _08034_);
  or _82353_ (_31584_, _31583_, _31582_);
  and _82354_ (_31585_, _31584_, _06615_);
  nor _82355_ (_31586_, _08596_, _13379_);
  or _82356_ (_31587_, _31586_, _31582_);
  or _82357_ (_31588_, _31587_, _06327_);
  and _82358_ (_31589_, _13387_, \oc8051_golden_model_1.P3 [4]);
  and _82359_ (_31590_, _30712_, _08657_);
  or _82360_ (_31592_, _31590_, _31589_);
  and _82361_ (_31593_, _31592_, _06352_);
  and _82362_ (_31594_, _30718_, _08034_);
  or _82363_ (_31595_, _31594_, _31582_);
  or _82364_ (_31596_, _31595_, _07275_);
  and _82365_ (_31597_, _08034_, \oc8051_golden_model_1.ACC [4]);
  or _82366_ (_31598_, _31597_, _31582_);
  and _82367_ (_31599_, _31598_, _07259_);
  and _82368_ (_31600_, _07260_, \oc8051_golden_model_1.P3 [4]);
  or _82369_ (_31601_, _31600_, _06474_);
  or _82370_ (_31603_, _31601_, _31599_);
  and _82371_ (_31604_, _31603_, _06357_);
  and _82372_ (_31605_, _31604_, _31596_);
  and _82373_ (_31606_, _30731_, _08657_);
  or _82374_ (_31607_, _31606_, _31589_);
  and _82375_ (_31608_, _31607_, _06356_);
  or _82376_ (_31609_, _31608_, _06410_);
  or _82377_ (_31610_, _31609_, _31605_);
  or _82378_ (_31611_, _31587_, _06772_);
  and _82379_ (_31612_, _31611_, _31610_);
  or _82380_ (_31614_, _31612_, _06417_);
  or _82381_ (_31615_, _31598_, _06426_);
  and _82382_ (_31616_, _31615_, _06353_);
  and _82383_ (_31617_, _31616_, _31614_);
  or _82384_ (_31618_, _31617_, _31593_);
  and _82385_ (_31619_, _31618_, _06346_);
  or _82386_ (_31620_, _31589_, _30746_);
  and _82387_ (_31621_, _31607_, _06345_);
  and _82388_ (_31622_, _31621_, _31620_);
  or _82389_ (_31623_, _31622_, _31619_);
  and _82390_ (_31625_, _31623_, _06340_);
  and _82391_ (_31626_, _30753_, _08657_);
  or _82392_ (_31627_, _31626_, _31589_);
  and _82393_ (_31628_, _31627_, _06339_);
  or _82394_ (_31629_, _31628_, _10153_);
  or _82395_ (_31630_, _31629_, _31625_);
  and _82396_ (_31631_, _31630_, _31588_);
  or _82397_ (_31632_, _31631_, _09572_);
  and _82398_ (_31633_, _09264_, _08034_);
  or _82399_ (_31634_, _31582_, _06333_);
  or _82400_ (_31636_, _31634_, _31633_);
  and _82401_ (_31637_, _31636_, _06313_);
  and _82402_ (_31638_, _31637_, _31632_);
  and _82403_ (_31639_, _30778_, _08034_);
  or _82404_ (_31640_, _31639_, _31582_);
  and _82405_ (_31641_, _31640_, _06037_);
  or _82406_ (_31642_, _31641_, _06277_);
  or _82407_ (_31643_, _31642_, _31638_);
  and _82408_ (_31644_, _08995_, _08034_);
  or _82409_ (_31645_, _31644_, _31582_);
  or _82410_ (_31647_, _31645_, _06278_);
  and _82411_ (_31648_, _31647_, _31643_);
  or _82412_ (_31649_, _31648_, _06502_);
  and _82413_ (_31650_, _30793_, _08034_);
  or _82414_ (_31651_, _31582_, _07334_);
  or _82415_ (_31652_, _31651_, _31650_);
  and _82416_ (_31653_, _31652_, _07337_);
  and _82417_ (_31654_, _31653_, _31649_);
  or _82418_ (_31655_, _31654_, _31585_);
  and _82419_ (_31656_, _31655_, _07339_);
  or _82420_ (_31658_, _31582_, _13360_);
  and _82421_ (_31659_, _31645_, _06507_);
  and _82422_ (_31660_, _31659_, _31658_);
  or _82423_ (_31661_, _31660_, _31656_);
  and _82424_ (_31662_, _31661_, _07331_);
  and _82425_ (_31663_, _31598_, _06610_);
  and _82426_ (_31664_, _31663_, _31658_);
  or _82427_ (_31665_, _31664_, _06509_);
  or _82428_ (_31666_, _31665_, _31662_);
  and _82429_ (_31667_, _30790_, _08034_);
  or _82430_ (_31669_, _31582_, _09107_);
  or _82431_ (_31670_, _31669_, _31667_);
  and _82432_ (_31671_, _31670_, _09112_);
  and _82433_ (_31672_, _31671_, _31666_);
  and _82434_ (_31673_, _30690_, _08034_);
  or _82435_ (_31674_, _31673_, _31582_);
  and _82436_ (_31675_, _31674_, _06602_);
  or _82437_ (_31676_, _31675_, _06639_);
  or _82438_ (_31677_, _31676_, _31672_);
  or _82439_ (_31678_, _31595_, _07048_);
  and _82440_ (_31680_, _31678_, _05990_);
  and _82441_ (_31681_, _31680_, _31677_);
  and _82442_ (_31682_, _31592_, _05989_);
  or _82443_ (_31683_, _31682_, _06646_);
  or _82444_ (_31684_, _31683_, _31681_);
  and _82445_ (_31685_, _30830_, _08034_);
  or _82446_ (_31686_, _31582_, _06651_);
  or _82447_ (_31687_, _31686_, _31685_);
  and _82448_ (_31688_, _31687_, _01442_);
  and _82449_ (_31689_, _31688_, _31684_);
  or _82450_ (_44236_, _31689_, _31581_);
  nor _82451_ (_31691_, \oc8051_golden_model_1.P3 [5], rst);
  nor _82452_ (_31692_, _31691_, _00000_);
  and _82453_ (_31693_, _13379_, \oc8051_golden_model_1.P3 [5]);
  and _82454_ (_31694_, _30842_, _08034_);
  or _82455_ (_31695_, _31694_, _31693_);
  and _82456_ (_31696_, _31695_, _06615_);
  and _82457_ (_31697_, _30848_, _08034_);
  or _82458_ (_31698_, _31697_, _31693_);
  or _82459_ (_31699_, _31698_, _07275_);
  and _82460_ (_31701_, _08034_, \oc8051_golden_model_1.ACC [5]);
  or _82461_ (_31702_, _31701_, _31693_);
  and _82462_ (_31703_, _31702_, _07259_);
  and _82463_ (_31704_, _07260_, \oc8051_golden_model_1.P3 [5]);
  or _82464_ (_31705_, _31704_, _06474_);
  or _82465_ (_31706_, _31705_, _31703_);
  and _82466_ (_31707_, _31706_, _06357_);
  and _82467_ (_31708_, _31707_, _31699_);
  and _82468_ (_31709_, _13387_, \oc8051_golden_model_1.P3 [5]);
  and _82469_ (_31710_, _30873_, _08657_);
  or _82470_ (_31712_, _31710_, _31709_);
  and _82471_ (_31713_, _31712_, _06356_);
  or _82472_ (_31714_, _31713_, _06410_);
  or _82473_ (_31715_, _31714_, _31708_);
  nor _82474_ (_31716_, _08305_, _13379_);
  or _82475_ (_31717_, _31716_, _31693_);
  or _82476_ (_31718_, _31717_, _06772_);
  and _82477_ (_31719_, _31718_, _31715_);
  or _82478_ (_31720_, _31719_, _06417_);
  or _82479_ (_31721_, _31702_, _06426_);
  and _82480_ (_31723_, _31721_, _06353_);
  and _82481_ (_31724_, _31723_, _31720_);
  and _82482_ (_31725_, _30888_, _08657_);
  or _82483_ (_31726_, _31725_, _31709_);
  and _82484_ (_31727_, _31726_, _06352_);
  or _82485_ (_31728_, _31727_, _06345_);
  or _82486_ (_31729_, _31728_, _31724_);
  or _82487_ (_31730_, _31709_, _30895_);
  and _82488_ (_31731_, _31730_, _31712_);
  or _82489_ (_31732_, _31731_, _06346_);
  and _82490_ (_31734_, _31732_, _06340_);
  and _82491_ (_31735_, _31734_, _31729_);
  and _82492_ (_31736_, _30902_, _08657_);
  or _82493_ (_31737_, _31736_, _31709_);
  and _82494_ (_31738_, _31737_, _06339_);
  or _82495_ (_31739_, _31738_, _10153_);
  or _82496_ (_31740_, _31739_, _31735_);
  or _82497_ (_31741_, _31717_, _06327_);
  and _82498_ (_31742_, _31741_, _31740_);
  or _82499_ (_31743_, _31742_, _09572_);
  and _82500_ (_31745_, _09218_, _08034_);
  or _82501_ (_31746_, _31693_, _06333_);
  or _82502_ (_31747_, _31746_, _31745_);
  and _82503_ (_31748_, _31747_, _06313_);
  and _82504_ (_31749_, _31748_, _31743_);
  and _82505_ (_31750_, _30928_, _08034_);
  or _82506_ (_31751_, _31750_, _31693_);
  and _82507_ (_31752_, _31751_, _06037_);
  or _82508_ (_31753_, _31752_, _06277_);
  or _82509_ (_31754_, _31753_, _31749_);
  and _82510_ (_31756_, _08954_, _08034_);
  or _82511_ (_31757_, _31756_, _31693_);
  or _82512_ (_31758_, _31757_, _06278_);
  and _82513_ (_31759_, _31758_, _31754_);
  or _82514_ (_31760_, _31759_, _06502_);
  and _82515_ (_31761_, _30942_, _08034_);
  or _82516_ (_31762_, _31693_, _07334_);
  or _82517_ (_31763_, _31762_, _31761_);
  and _82518_ (_31764_, _31763_, _07337_);
  and _82519_ (_31765_, _31764_, _31760_);
  or _82520_ (_31767_, _31765_, _31696_);
  and _82521_ (_31768_, _31767_, _07339_);
  or _82522_ (_31769_, _31693_, _13359_);
  and _82523_ (_31770_, _31757_, _06507_);
  and _82524_ (_31771_, _31770_, _31769_);
  or _82525_ (_31772_, _31771_, _31768_);
  and _82526_ (_31773_, _31772_, _07331_);
  and _82527_ (_31774_, _31702_, _06610_);
  and _82528_ (_31775_, _31774_, _31769_);
  or _82529_ (_31776_, _31775_, _06509_);
  or _82530_ (_31778_, _31776_, _31773_);
  and _82531_ (_31779_, _30940_, _08034_);
  or _82532_ (_31780_, _31693_, _09107_);
  or _82533_ (_31781_, _31780_, _31779_);
  and _82534_ (_31782_, _31781_, _09112_);
  and _82535_ (_31783_, _31782_, _31778_);
  and _82536_ (_31784_, _30840_, _08034_);
  or _82537_ (_31785_, _31784_, _31693_);
  and _82538_ (_31786_, _31785_, _06602_);
  or _82539_ (_31787_, _31786_, _06639_);
  or _82540_ (_31789_, _31787_, _31783_);
  or _82541_ (_31790_, _31698_, _07048_);
  and _82542_ (_31791_, _31790_, _05990_);
  and _82543_ (_31792_, _31791_, _31789_);
  and _82544_ (_31793_, _31726_, _05989_);
  or _82545_ (_31794_, _31793_, _06646_);
  or _82546_ (_31795_, _31794_, _31792_);
  and _82547_ (_31796_, _30980_, _08034_);
  or _82548_ (_31797_, _31693_, _06651_);
  or _82549_ (_31798_, _31797_, _31796_);
  and _82550_ (_31800_, _31798_, _01442_);
  and _82551_ (_31801_, _31800_, _31795_);
  or _82552_ (_44237_, _31801_, _31692_);
  nor _82553_ (_31802_, \oc8051_golden_model_1.P3 [6], rst);
  nor _82554_ (_31803_, _31802_, _00000_);
  and _82555_ (_31804_, _13379_, \oc8051_golden_model_1.P3 [6]);
  and _82556_ (_31805_, _30992_, _08034_);
  or _82557_ (_31806_, _31805_, _31804_);
  and _82558_ (_31807_, _31806_, _06615_);
  nor _82559_ (_31808_, _08209_, _13379_);
  or _82560_ (_31810_, _31808_, _31804_);
  or _82561_ (_31811_, _31810_, _06327_);
  and _82562_ (_31812_, _13387_, \oc8051_golden_model_1.P3 [6]);
  and _82563_ (_31813_, _31013_, _08657_);
  or _82564_ (_31814_, _31813_, _31812_);
  and _82565_ (_31815_, _31814_, _06352_);
  and _82566_ (_31816_, _31018_, _08034_);
  or _82567_ (_31817_, _31816_, _31804_);
  or _82568_ (_31818_, _31817_, _07275_);
  and _82569_ (_31819_, _08034_, \oc8051_golden_model_1.ACC [6]);
  or _82570_ (_31821_, _31819_, _31804_);
  and _82571_ (_31822_, _31821_, _07259_);
  and _82572_ (_31823_, _07260_, \oc8051_golden_model_1.P3 [6]);
  or _82573_ (_31824_, _31823_, _06474_);
  or _82574_ (_31825_, _31824_, _31822_);
  and _82575_ (_31826_, _31825_, _06357_);
  and _82576_ (_31827_, _31826_, _31818_);
  and _82577_ (_31828_, _31032_, _08657_);
  or _82578_ (_31829_, _31828_, _31812_);
  and _82579_ (_31830_, _31829_, _06356_);
  or _82580_ (_31832_, _31830_, _06410_);
  or _82581_ (_31833_, _31832_, _31827_);
  or _82582_ (_31834_, _31810_, _06772_);
  and _82583_ (_31835_, _31834_, _31833_);
  or _82584_ (_31836_, _31835_, _06417_);
  or _82585_ (_31837_, _31821_, _06426_);
  and _82586_ (_31838_, _31837_, _06353_);
  and _82587_ (_31839_, _31838_, _31836_);
  or _82588_ (_31840_, _31839_, _31815_);
  and _82589_ (_31841_, _31840_, _06346_);
  or _82590_ (_31843_, _31812_, _31049_);
  and _82591_ (_31844_, _31829_, _06345_);
  and _82592_ (_31845_, _31844_, _31843_);
  or _82593_ (_31846_, _31845_, _31841_);
  and _82594_ (_31847_, _31846_, _06340_);
  and _82595_ (_31848_, _31055_, _08657_);
  or _82596_ (_31849_, _31848_, _31812_);
  and _82597_ (_31850_, _31849_, _06339_);
  or _82598_ (_31851_, _31850_, _10153_);
  or _82599_ (_31852_, _31851_, _31847_);
  and _82600_ (_31854_, _31852_, _31811_);
  or _82601_ (_31855_, _31854_, _09572_);
  and _82602_ (_31856_, _09172_, _08034_);
  or _82603_ (_31857_, _31804_, _06333_);
  or _82604_ (_31858_, _31857_, _31856_);
  and _82605_ (_31859_, _31858_, _06313_);
  and _82606_ (_31860_, _31859_, _31855_);
  and _82607_ (_31861_, _31082_, _08034_);
  or _82608_ (_31862_, _31861_, _31804_);
  and _82609_ (_31863_, _31862_, _06037_);
  or _82610_ (_31865_, _31863_, _06277_);
  or _82611_ (_31866_, _31865_, _31860_);
  and _82612_ (_31867_, _15853_, _08034_);
  or _82613_ (_31868_, _31867_, _31804_);
  or _82614_ (_31869_, _31868_, _06278_);
  and _82615_ (_31870_, _31869_, _31866_);
  or _82616_ (_31871_, _31870_, _06502_);
  and _82617_ (_31872_, _31096_, _08034_);
  or _82618_ (_31873_, _31804_, _07334_);
  or _82619_ (_31874_, _31873_, _31872_);
  and _82620_ (_31876_, _31874_, _07337_);
  and _82621_ (_31877_, _31876_, _31871_);
  or _82622_ (_31878_, _31877_, _31807_);
  and _82623_ (_31879_, _31878_, _07339_);
  or _82624_ (_31880_, _31804_, _13358_);
  and _82625_ (_31881_, _31868_, _06507_);
  and _82626_ (_31882_, _31881_, _31880_);
  or _82627_ (_31883_, _31882_, _31879_);
  and _82628_ (_31884_, _31883_, _07331_);
  and _82629_ (_31885_, _31821_, _06610_);
  and _82630_ (_31887_, _31885_, _31880_);
  or _82631_ (_31888_, _31887_, _06509_);
  or _82632_ (_31889_, _31888_, _31884_);
  and _82633_ (_31890_, _31094_, _08034_);
  or _82634_ (_31891_, _31804_, _09107_);
  or _82635_ (_31892_, _31891_, _31890_);
  and _82636_ (_31893_, _31892_, _09112_);
  and _82637_ (_31894_, _31893_, _31889_);
  and _82638_ (_31895_, _30990_, _08034_);
  or _82639_ (_31896_, _31895_, _31804_);
  and _82640_ (_31898_, _31896_, _06602_);
  or _82641_ (_31899_, _31898_, _06639_);
  or _82642_ (_31900_, _31899_, _31894_);
  or _82643_ (_31901_, _31817_, _07048_);
  and _82644_ (_31902_, _31901_, _05990_);
  and _82645_ (_31903_, _31902_, _31900_);
  and _82646_ (_31904_, _31814_, _05989_);
  or _82647_ (_31905_, _31904_, _06646_);
  or _82648_ (_31906_, _31905_, _31903_);
  and _82649_ (_31907_, _31133_, _08034_);
  or _82650_ (_31909_, _31804_, _06651_);
  or _82651_ (_31910_, _31909_, _31907_);
  and _82652_ (_31911_, _31910_, _01442_);
  and _82653_ (_31912_, _31911_, _31906_);
  or _82654_ (_44238_, _31912_, _31803_);
  nor _82655_ (_31913_, \oc8051_golden_model_1.P0 [0], rst);
  nor _82656_ (_31914_, _31913_, _00000_);
  and _82657_ (_31915_, _13248_, _08039_);
  and _82658_ (_31916_, _13482_, \oc8051_golden_model_1.P0 [0]);
  and _82659_ (_31917_, _08039_, _09008_);
  or _82660_ (_31919_, _31917_, _31916_);
  nand _82661_ (_31920_, _31919_, _06507_);
  nor _82662_ (_31921_, _31920_, _31915_);
  and _82663_ (_31922_, _30107_, _08039_);
  or _82664_ (_31923_, _31922_, _31916_);
  and _82665_ (_31924_, _31923_, _06615_);
  or _82666_ (_31925_, _31916_, _31915_);
  or _82667_ (_31926_, _31925_, _07275_);
  and _82668_ (_31927_, _08039_, \oc8051_golden_model_1.ACC [0]);
  or _82669_ (_31928_, _31927_, _31916_);
  and _82670_ (_31930_, _31928_, _07259_);
  and _82671_ (_31931_, _07260_, \oc8051_golden_model_1.P0 [0]);
  or _82672_ (_31932_, _31931_, _06474_);
  or _82673_ (_31933_, _31932_, _31930_);
  and _82674_ (_31934_, _31933_, _06357_);
  and _82675_ (_31935_, _31934_, _31926_);
  and _82676_ (_31936_, _13490_, \oc8051_golden_model_1.P0 [0]);
  and _82677_ (_31937_, _30137_, _07993_);
  or _82678_ (_31938_, _31937_, _31936_);
  and _82679_ (_31939_, _31938_, _06356_);
  or _82680_ (_31941_, _31939_, _31935_);
  and _82681_ (_31942_, _31941_, _06772_);
  and _82682_ (_31943_, _08039_, _07250_);
  or _82683_ (_31944_, _31943_, _31916_);
  and _82684_ (_31945_, _31944_, _06410_);
  or _82685_ (_31946_, _31945_, _06417_);
  or _82686_ (_31947_, _31946_, _31942_);
  or _82687_ (_31948_, _31928_, _06426_);
  and _82688_ (_31949_, _31948_, _06353_);
  and _82689_ (_31950_, _31949_, _31947_);
  and _82690_ (_31952_, _31916_, _06352_);
  or _82691_ (_31953_, _31952_, _06345_);
  or _82692_ (_31954_, _31953_, _31950_);
  or _82693_ (_31955_, _31925_, _06346_);
  and _82694_ (_31956_, _31955_, _06340_);
  and _82695_ (_31957_, _31956_, _31954_);
  or _82696_ (_31958_, _31936_, _16663_);
  and _82697_ (_31959_, _31958_, _06339_);
  and _82698_ (_31960_, _31959_, _31938_);
  or _82699_ (_31961_, _31960_, _10153_);
  or _82700_ (_31963_, _31961_, _31957_);
  or _82701_ (_31964_, _31944_, _06327_);
  and _82702_ (_31965_, _31964_, _31963_);
  or _82703_ (_31966_, _31965_, _09572_);
  and _82704_ (_31967_, _09447_, _08039_);
  or _82705_ (_31968_, _31916_, _06333_);
  or _82706_ (_31969_, _31968_, _31967_);
  and _82707_ (_31970_, _31969_, _06313_);
  and _82708_ (_31971_, _31970_, _31966_);
  and _82709_ (_31972_, _30185_, _08039_);
  or _82710_ (_31974_, _31972_, _31916_);
  and _82711_ (_31975_, _31974_, _06037_);
  or _82712_ (_31976_, _31975_, _06277_);
  or _82713_ (_31977_, _31976_, _31971_);
  or _82714_ (_31978_, _31919_, _06278_);
  and _82715_ (_31979_, _31978_, _31977_);
  or _82716_ (_31980_, _31979_, _06502_);
  and _82717_ (_31981_, _30198_, _08039_);
  or _82718_ (_31982_, _31916_, _07334_);
  or _82719_ (_31983_, _31982_, _31981_);
  and _82720_ (_31985_, _31983_, _07337_);
  and _82721_ (_31986_, _31985_, _31980_);
  or _82722_ (_31987_, _31986_, _31924_);
  and _82723_ (_31988_, _31987_, _07339_);
  or _82724_ (_31989_, _31988_, _31921_);
  and _82725_ (_31990_, _31989_, _07331_);
  or _82726_ (_31991_, _31916_, _30209_);
  and _82727_ (_31992_, _31928_, _06610_);
  and _82728_ (_31993_, _31992_, _31991_);
  or _82729_ (_31994_, _31993_, _06509_);
  or _82730_ (_31996_, _31994_, _31990_);
  and _82731_ (_31997_, _30197_, _08039_);
  or _82732_ (_31998_, _31916_, _09107_);
  or _82733_ (_31999_, _31998_, _31997_);
  and _82734_ (_32000_, _31999_, _09112_);
  and _82735_ (_32001_, _32000_, _31996_);
  and _82736_ (_32002_, _30105_, _08039_);
  or _82737_ (_32003_, _32002_, _31916_);
  and _82738_ (_32004_, _32003_, _06602_);
  or _82739_ (_32005_, _32004_, _06639_);
  or _82740_ (_32007_, _32005_, _32001_);
  or _82741_ (_32008_, _31925_, _07048_);
  and _82742_ (_32009_, _32008_, _05990_);
  and _82743_ (_32010_, _32009_, _32007_);
  and _82744_ (_32011_, _31916_, _05989_);
  or _82745_ (_32012_, _32011_, _06646_);
  or _82746_ (_32013_, _32012_, _32010_);
  or _82747_ (_32014_, _31925_, _06651_);
  and _82748_ (_32015_, _32014_, _01442_);
  and _82749_ (_32016_, _32015_, _32013_);
  or _82750_ (_44240_, _32016_, _31914_);
  nor _82751_ (_32018_, \oc8051_golden_model_1.P0 [1], rst);
  nor _82752_ (_32019_, _32018_, _00000_);
  nand _82753_ (_32020_, _08039_, _07160_);
  or _82754_ (_32021_, _08039_, \oc8051_golden_model_1.P0 [1]);
  and _82755_ (_32022_, _32021_, _06277_);
  and _82756_ (_32023_, _32022_, _32020_);
  and _82757_ (_32024_, _13482_, \oc8051_golden_model_1.P0 [1]);
  nor _82758_ (_32025_, _13482_, _07448_);
  or _82759_ (_32026_, _32025_, _32024_);
  or _82760_ (_32028_, _32026_, _06772_);
  and _82761_ (_32029_, _30245_, _08039_);
  not _82762_ (_32030_, _32029_);
  and _82763_ (_32031_, _32030_, _32021_);
  or _82764_ (_32032_, _32031_, _07275_);
  nand _82765_ (_32033_, _08039_, _06097_);
  and _82766_ (_32034_, _32033_, _32021_);
  and _82767_ (_32035_, _32034_, _07259_);
  and _82768_ (_32036_, _07260_, \oc8051_golden_model_1.P0 [1]);
  or _82769_ (_32037_, _32036_, _06474_);
  or _82770_ (_32039_, _32037_, _32035_);
  and _82771_ (_32040_, _32039_, _06357_);
  and _82772_ (_32041_, _32040_, _32032_);
  and _82773_ (_32042_, _13490_, \oc8051_golden_model_1.P0 [1]);
  and _82774_ (_32043_, _30272_, _07993_);
  or _82775_ (_32044_, _32043_, _32042_);
  and _82776_ (_32045_, _32044_, _06356_);
  or _82777_ (_32046_, _32045_, _06410_);
  or _82778_ (_32047_, _32046_, _32041_);
  and _82779_ (_32048_, _32047_, _32028_);
  or _82780_ (_32050_, _32048_, _06417_);
  or _82781_ (_32051_, _32034_, _06426_);
  and _82782_ (_32052_, _32051_, _06353_);
  and _82783_ (_32053_, _32052_, _32050_);
  and _82784_ (_32054_, _30283_, _07993_);
  or _82785_ (_32055_, _32054_, _32042_);
  and _82786_ (_32056_, _32055_, _06352_);
  or _82787_ (_32057_, _32056_, _06345_);
  or _82788_ (_32058_, _32057_, _32053_);
  and _82789_ (_32059_, _32043_, _30291_);
  or _82790_ (_32061_, _32042_, _06346_);
  or _82791_ (_32062_, _32061_, _32059_);
  and _82792_ (_32063_, _32062_, _32058_);
  and _82793_ (_32064_, _32063_, _06340_);
  and _82794_ (_32065_, _30297_, _07993_);
  or _82795_ (_32066_, _32042_, _32065_);
  and _82796_ (_32067_, _32066_, _06339_);
  or _82797_ (_32068_, _32067_, _10153_);
  or _82798_ (_32069_, _32068_, _32064_);
  or _82799_ (_32070_, _32026_, _06327_);
  and _82800_ (_32072_, _32070_, _32069_);
  or _82801_ (_32073_, _32072_, _09572_);
  and _82802_ (_32074_, _09402_, _08039_);
  or _82803_ (_32075_, _32024_, _06333_);
  or _82804_ (_32076_, _32075_, _32074_);
  and _82805_ (_32077_, _32076_, _06313_);
  and _82806_ (_32078_, _32077_, _32073_);
  and _82807_ (_32079_, _30325_, _08039_);
  or _82808_ (_32080_, _32079_, _32024_);
  and _82809_ (_32081_, _32080_, _06037_);
  or _82810_ (_32083_, _32081_, _32078_);
  and _82811_ (_32084_, _32083_, _06278_);
  or _82812_ (_32085_, _32084_, _32023_);
  and _82813_ (_32086_, _32085_, _07334_);
  or _82814_ (_32087_, _30339_, _13482_);
  and _82815_ (_32088_, _32021_, _06502_);
  and _82816_ (_32089_, _32088_, _32087_);
  or _82817_ (_32090_, _32089_, _32086_);
  and _82818_ (_32091_, _32090_, _07337_);
  or _82819_ (_32092_, _30348_, _13482_);
  and _82820_ (_32094_, _32021_, _06615_);
  and _82821_ (_32095_, _32094_, _32092_);
  or _82822_ (_32096_, _32095_, _32091_);
  and _82823_ (_32097_, _32096_, _07339_);
  or _82824_ (_32098_, _30337_, _13482_);
  and _82825_ (_32099_, _32021_, _06507_);
  and _82826_ (_32100_, _32099_, _32098_);
  or _82827_ (_32101_, _32100_, _32097_);
  and _82828_ (_32102_, _32101_, _07331_);
  or _82829_ (_32103_, _32024_, _30360_);
  and _82830_ (_32105_, _32034_, _06610_);
  and _82831_ (_32106_, _32105_, _32103_);
  or _82832_ (_32107_, _32106_, _32102_);
  and _82833_ (_32108_, _32107_, _06603_);
  or _82834_ (_32109_, _32020_, _30360_);
  and _82835_ (_32110_, _32021_, _06509_);
  and _82836_ (_32111_, _32110_, _32109_);
  or _82837_ (_32112_, _30346_, _13482_);
  and _82838_ (_32113_, _32021_, _06602_);
  and _82839_ (_32114_, _32113_, _32112_);
  or _82840_ (_32116_, _32114_, _06639_);
  or _82841_ (_32117_, _32116_, _32111_);
  or _82842_ (_32118_, _32117_, _32108_);
  or _82843_ (_32119_, _32031_, _07048_);
  and _82844_ (_32120_, _32119_, _05990_);
  and _82845_ (_32121_, _32120_, _32118_);
  and _82846_ (_32122_, _32055_, _05989_);
  or _82847_ (_32123_, _32122_, _06646_);
  or _82848_ (_32124_, _32123_, _32121_);
  or _82849_ (_32125_, _32024_, _06651_);
  or _82850_ (_32127_, _32125_, _32029_);
  and _82851_ (_32128_, _32127_, _01442_);
  and _82852_ (_32129_, _32128_, _32124_);
  or _82853_ (_44241_, _32129_, _32019_);
  nor _82854_ (_32130_, \oc8051_golden_model_1.P0 [2], rst);
  nor _82855_ (_32131_, _32130_, _00000_);
  and _82856_ (_32132_, _13482_, \oc8051_golden_model_1.P0 [2]);
  and _82857_ (_32133_, _30393_, _08039_);
  or _82858_ (_32134_, _32133_, _32132_);
  and _82859_ (_32135_, _32134_, _06615_);
  nor _82860_ (_32137_, _13482_, _07854_);
  or _82861_ (_32138_, _32137_, _32132_);
  or _82862_ (_32139_, _32138_, _06327_);
  or _82863_ (_32140_, _32138_, _06772_);
  and _82864_ (_32141_, _30403_, _08039_);
  or _82865_ (_32142_, _32141_, _32132_);
  or _82866_ (_32143_, _32142_, _07275_);
  and _82867_ (_32144_, _08039_, \oc8051_golden_model_1.ACC [2]);
  or _82868_ (_32145_, _32144_, _32132_);
  and _82869_ (_32146_, _32145_, _07259_);
  and _82870_ (_32148_, _07260_, \oc8051_golden_model_1.P0 [2]);
  or _82871_ (_32149_, _32148_, _06474_);
  or _82872_ (_32150_, _32149_, _32146_);
  and _82873_ (_32151_, _32150_, _06357_);
  and _82874_ (_32152_, _32151_, _32143_);
  and _82875_ (_32153_, _13490_, \oc8051_golden_model_1.P0 [2]);
  and _82876_ (_32154_, _30428_, _07993_);
  or _82877_ (_32155_, _32154_, _32153_);
  and _82878_ (_32156_, _32155_, _06356_);
  or _82879_ (_32157_, _32156_, _06410_);
  or _82880_ (_32159_, _32157_, _32152_);
  and _82881_ (_32160_, _32159_, _32140_);
  or _82882_ (_32161_, _32160_, _06417_);
  or _82883_ (_32162_, _32145_, _06426_);
  and _82884_ (_32163_, _32162_, _06353_);
  and _82885_ (_32164_, _32163_, _32161_);
  and _82886_ (_32165_, _30440_, _07993_);
  or _82887_ (_32166_, _32165_, _32153_);
  and _82888_ (_32167_, _32166_, _06352_);
  or _82889_ (_32168_, _32167_, _06345_);
  or _82890_ (_32170_, _32168_, _32164_);
  and _82891_ (_32171_, _32154_, _30447_);
  or _82892_ (_32172_, _32153_, _06346_);
  or _82893_ (_32173_, _32172_, _32171_);
  and _82894_ (_32174_, _32173_, _06340_);
  and _82895_ (_32175_, _32174_, _32170_);
  and _82896_ (_32176_, _30454_, _07993_);
  or _82897_ (_32177_, _32176_, _32153_);
  and _82898_ (_32178_, _32177_, _06339_);
  or _82899_ (_32179_, _32178_, _10153_);
  or _82900_ (_32181_, _32179_, _32175_);
  and _82901_ (_32182_, _32181_, _32139_);
  or _82902_ (_32183_, _32182_, _09572_);
  and _82903_ (_32184_, _09356_, _08039_);
  or _82904_ (_32185_, _32132_, _06333_);
  or _82905_ (_32186_, _32185_, _32184_);
  and _82906_ (_32187_, _32186_, _06313_);
  and _82907_ (_32188_, _32187_, _32183_);
  and _82908_ (_32189_, _30479_, _08039_);
  or _82909_ (_32190_, _32189_, _32132_);
  and _82910_ (_32192_, _32190_, _06037_);
  or _82911_ (_32193_, _32192_, _06277_);
  or _82912_ (_32194_, _32193_, _32188_);
  and _82913_ (_32195_, _08039_, _09057_);
  or _82914_ (_32196_, _32195_, _32132_);
  or _82915_ (_32197_, _32196_, _06278_);
  and _82916_ (_32198_, _32197_, _32194_);
  or _82917_ (_32199_, _32198_, _06502_);
  and _82918_ (_32200_, _30493_, _08039_);
  or _82919_ (_32201_, _32132_, _07334_);
  or _82920_ (_32203_, _32201_, _32200_);
  and _82921_ (_32204_, _32203_, _07337_);
  and _82922_ (_32205_, _32204_, _32199_);
  or _82923_ (_32206_, _32205_, _32135_);
  and _82924_ (_32207_, _32206_, _07339_);
  or _82925_ (_32208_, _32132_, _13362_);
  and _82926_ (_32209_, _32196_, _06507_);
  and _82927_ (_32210_, _32209_, _32208_);
  or _82928_ (_32211_, _32210_, _32207_);
  and _82929_ (_32212_, _32211_, _07331_);
  and _82930_ (_32214_, _32145_, _06610_);
  and _82931_ (_32215_, _32214_, _32208_);
  or _82932_ (_32216_, _32215_, _06509_);
  or _82933_ (_32217_, _32216_, _32212_);
  and _82934_ (_32218_, _30491_, _08039_);
  or _82935_ (_32219_, _32132_, _09107_);
  or _82936_ (_32220_, _32219_, _32218_);
  and _82937_ (_32221_, _32220_, _09112_);
  and _82938_ (_32222_, _32221_, _32217_);
  and _82939_ (_32223_, _30391_, _08039_);
  or _82940_ (_32225_, _32223_, _32132_);
  and _82941_ (_32226_, _32225_, _06602_);
  or _82942_ (_32227_, _32226_, _06639_);
  or _82943_ (_32228_, _32227_, _32222_);
  or _82944_ (_32229_, _32142_, _07048_);
  and _82945_ (_32230_, _32229_, _05990_);
  and _82946_ (_32231_, _32230_, _32228_);
  and _82947_ (_32232_, _32166_, _05989_);
  or _82948_ (_32233_, _32232_, _06646_);
  or _82949_ (_32234_, _32233_, _32231_);
  and _82950_ (_32236_, _30531_, _08039_);
  or _82951_ (_32237_, _32132_, _06651_);
  or _82952_ (_32238_, _32237_, _32236_);
  and _82953_ (_32239_, _32238_, _01442_);
  and _82954_ (_32240_, _32239_, _32234_);
  or _82955_ (_44242_, _32240_, _32131_);
  nor _82956_ (_32241_, \oc8051_golden_model_1.P0 [3], rst);
  nor _82957_ (_32242_, _32241_, _00000_);
  and _82958_ (_32243_, _13482_, \oc8051_golden_model_1.P0 [3]);
  and _82959_ (_32244_, _30543_, _08039_);
  or _82960_ (_32246_, _32244_, _32243_);
  and _82961_ (_32247_, _32246_, _06615_);
  nor _82962_ (_32248_, _13482_, _07680_);
  or _82963_ (_32249_, _32248_, _32243_);
  or _82964_ (_32250_, _32249_, _06327_);
  and _82965_ (_32251_, _30552_, _08039_);
  or _82966_ (_32252_, _32251_, _32243_);
  or _82967_ (_32253_, _32252_, _07275_);
  and _82968_ (_32254_, _08039_, \oc8051_golden_model_1.ACC [3]);
  or _82969_ (_32255_, _32254_, _32243_);
  and _82970_ (_32257_, _32255_, _07259_);
  and _82971_ (_32258_, _07260_, \oc8051_golden_model_1.P0 [3]);
  or _82972_ (_32259_, _32258_, _06474_);
  or _82973_ (_32260_, _32259_, _32257_);
  and _82974_ (_32261_, _32260_, _06357_);
  and _82975_ (_32262_, _32261_, _32253_);
  and _82976_ (_32263_, _13490_, \oc8051_golden_model_1.P0 [3]);
  and _82977_ (_32264_, _30577_, _07993_);
  or _82978_ (_32265_, _32264_, _32263_);
  and _82979_ (_32266_, _32265_, _06356_);
  or _82980_ (_32268_, _32266_, _06410_);
  or _82981_ (_32269_, _32268_, _32262_);
  or _82982_ (_32270_, _32249_, _06772_);
  and _82983_ (_32271_, _32270_, _32269_);
  or _82984_ (_32272_, _32271_, _06417_);
  or _82985_ (_32273_, _32255_, _06426_);
  and _82986_ (_32274_, _32273_, _06353_);
  and _82987_ (_32275_, _32274_, _32272_);
  and _82988_ (_32276_, _30590_, _07993_);
  or _82989_ (_32277_, _32276_, _32263_);
  and _82990_ (_32279_, _32277_, _06352_);
  or _82991_ (_32280_, _32279_, _06345_);
  or _82992_ (_32281_, _32280_, _32275_);
  or _82993_ (_32282_, _32263_, _30597_);
  and _82994_ (_32283_, _32282_, _32265_);
  or _82995_ (_32284_, _32283_, _06346_);
  and _82996_ (_32285_, _32284_, _06340_);
  and _82997_ (_32286_, _32285_, _32281_);
  and _82998_ (_32287_, _30603_, _07993_);
  or _82999_ (_32288_, _32287_, _32263_);
  and _83000_ (_32290_, _32288_, _06339_);
  or _83001_ (_32291_, _32290_, _10153_);
  or _83002_ (_32292_, _32291_, _32286_);
  and _83003_ (_32293_, _32292_, _32250_);
  or _83004_ (_32294_, _32293_, _09572_);
  and _83005_ (_32295_, _09310_, _08039_);
  or _83006_ (_32296_, _32243_, _06333_);
  or _83007_ (_32297_, _32296_, _32295_);
  and _83008_ (_32298_, _32297_, _06313_);
  and _83009_ (_32299_, _32298_, _32294_);
  and _83010_ (_32301_, _30629_, _08039_);
  or _83011_ (_32302_, _32301_, _32243_);
  and _83012_ (_32303_, _32302_, _06037_);
  or _83013_ (_32304_, _32303_, _06277_);
  or _83014_ (_32305_, _32304_, _32299_);
  and _83015_ (_32306_, _08039_, _09014_);
  or _83016_ (_32307_, _32306_, _32243_);
  or _83017_ (_32308_, _32307_, _06278_);
  and _83018_ (_32309_, _32308_, _32305_);
  or _83019_ (_32310_, _32309_, _06502_);
  and _83020_ (_32312_, _30643_, _08039_);
  or _83021_ (_32313_, _32243_, _07334_);
  or _83022_ (_32314_, _32313_, _32312_);
  and _83023_ (_32315_, _32314_, _07337_);
  and _83024_ (_32316_, _32315_, _32310_);
  or _83025_ (_32317_, _32316_, _32247_);
  and _83026_ (_32318_, _32317_, _07339_);
  or _83027_ (_32319_, _32243_, _13361_);
  and _83028_ (_32320_, _32307_, _06507_);
  and _83029_ (_32321_, _32320_, _32319_);
  or _83030_ (_32323_, _32321_, _32318_);
  and _83031_ (_32324_, _32323_, _07331_);
  and _83032_ (_32325_, _32255_, _06610_);
  and _83033_ (_32326_, _32325_, _32319_);
  or _83034_ (_32327_, _32326_, _06509_);
  or _83035_ (_32328_, _32327_, _32324_);
  and _83036_ (_32329_, _30641_, _08039_);
  or _83037_ (_32330_, _32243_, _09107_);
  or _83038_ (_32331_, _32330_, _32329_);
  and _83039_ (_32332_, _32331_, _09112_);
  and _83040_ (_32334_, _32332_, _32328_);
  and _83041_ (_32335_, _30541_, _08039_);
  or _83042_ (_32336_, _32335_, _32243_);
  and _83043_ (_32337_, _32336_, _06602_);
  or _83044_ (_32338_, _32337_, _06639_);
  or _83045_ (_32339_, _32338_, _32334_);
  or _83046_ (_32340_, _32252_, _07048_);
  and _83047_ (_32341_, _32340_, _05990_);
  and _83048_ (_32342_, _32341_, _32339_);
  and _83049_ (_32343_, _32277_, _05989_);
  or _83050_ (_32345_, _32343_, _06646_);
  or _83051_ (_32346_, _32345_, _32342_);
  and _83052_ (_32347_, _30680_, _08039_);
  or _83053_ (_32348_, _32243_, _06651_);
  or _83054_ (_32349_, _32348_, _32347_);
  and _83055_ (_32350_, _32349_, _01442_);
  and _83056_ (_32351_, _32350_, _32346_);
  or _83057_ (_44244_, _32351_, _32242_);
  nor _83058_ (_32352_, \oc8051_golden_model_1.P0 [4], rst);
  nor _83059_ (_32353_, _32352_, _00000_);
  and _83060_ (_32355_, _13482_, \oc8051_golden_model_1.P0 [4]);
  and _83061_ (_32356_, _30693_, _08039_);
  or _83062_ (_32357_, _32356_, _32355_);
  and _83063_ (_32358_, _32357_, _06615_);
  nor _83064_ (_32359_, _08596_, _13482_);
  or _83065_ (_32360_, _32359_, _32355_);
  or _83066_ (_32361_, _32360_, _06327_);
  and _83067_ (_32362_, _13490_, \oc8051_golden_model_1.P0 [4]);
  and _83068_ (_32363_, _30712_, _07993_);
  or _83069_ (_32364_, _32363_, _32362_);
  and _83070_ (_32366_, _32364_, _06352_);
  and _83071_ (_32367_, _30718_, _08039_);
  or _83072_ (_32368_, _32367_, _32355_);
  or _83073_ (_32369_, _32368_, _07275_);
  and _83074_ (_32370_, _08039_, \oc8051_golden_model_1.ACC [4]);
  or _83075_ (_32371_, _32370_, _32355_);
  and _83076_ (_32372_, _32371_, _07259_);
  and _83077_ (_32373_, _07260_, \oc8051_golden_model_1.P0 [4]);
  or _83078_ (_32374_, _32373_, _06474_);
  or _83079_ (_32375_, _32374_, _32372_);
  and _83080_ (_32377_, _32375_, _06357_);
  and _83081_ (_32378_, _32377_, _32369_);
  and _83082_ (_32379_, _30731_, _07993_);
  or _83083_ (_32380_, _32379_, _32362_);
  and _83084_ (_32381_, _32380_, _06356_);
  or _83085_ (_32382_, _32381_, _06410_);
  or _83086_ (_32383_, _32382_, _32378_);
  or _83087_ (_32384_, _32360_, _06772_);
  and _83088_ (_32385_, _32384_, _32383_);
  or _83089_ (_32386_, _32385_, _06417_);
  or _83090_ (_32388_, _32371_, _06426_);
  and _83091_ (_32389_, _32388_, _06353_);
  and _83092_ (_32390_, _32389_, _32386_);
  or _83093_ (_32391_, _32390_, _32366_);
  and _83094_ (_32392_, _32391_, _06346_);
  or _83095_ (_32393_, _32362_, _30746_);
  and _83096_ (_32394_, _32380_, _06345_);
  and _83097_ (_32395_, _32394_, _32393_);
  or _83098_ (_32396_, _32395_, _32392_);
  and _83099_ (_32397_, _32396_, _06340_);
  and _83100_ (_32399_, _30753_, _07993_);
  or _83101_ (_32400_, _32399_, _32362_);
  and _83102_ (_32401_, _32400_, _06339_);
  or _83103_ (_32402_, _32401_, _10153_);
  or _83104_ (_32403_, _32402_, _32397_);
  and _83105_ (_32404_, _32403_, _32361_);
  or _83106_ (_32405_, _32404_, _09572_);
  and _83107_ (_32406_, _09264_, _08039_);
  or _83108_ (_32407_, _32355_, _06333_);
  or _83109_ (_32408_, _32407_, _32406_);
  and _83110_ (_32410_, _32408_, _06313_);
  and _83111_ (_32411_, _32410_, _32405_);
  and _83112_ (_32412_, _30778_, _08039_);
  or _83113_ (_32413_, _32412_, _32355_);
  and _83114_ (_32414_, _32413_, _06037_);
  or _83115_ (_32415_, _32414_, _06277_);
  or _83116_ (_32416_, _32415_, _32411_);
  and _83117_ (_32417_, _08995_, _08039_);
  or _83118_ (_32418_, _32417_, _32355_);
  or _83119_ (_32419_, _32418_, _06278_);
  and _83120_ (_32421_, _32419_, _32416_);
  or _83121_ (_32422_, _32421_, _06502_);
  and _83122_ (_32423_, _30793_, _08039_);
  or _83123_ (_32424_, _32355_, _07334_);
  or _83124_ (_32425_, _32424_, _32423_);
  and _83125_ (_32426_, _32425_, _07337_);
  and _83126_ (_32427_, _32426_, _32422_);
  or _83127_ (_32428_, _32427_, _32358_);
  and _83128_ (_32429_, _32428_, _07339_);
  or _83129_ (_32430_, _32355_, _13360_);
  and _83130_ (_32432_, _32418_, _06507_);
  and _83131_ (_32433_, _32432_, _32430_);
  or _83132_ (_32434_, _32433_, _32429_);
  and _83133_ (_32435_, _32434_, _07331_);
  and _83134_ (_32436_, _32371_, _06610_);
  and _83135_ (_32437_, _32436_, _32430_);
  or _83136_ (_32438_, _32437_, _06509_);
  or _83137_ (_32439_, _32438_, _32435_);
  and _83138_ (_32440_, _30790_, _08039_);
  or _83139_ (_32441_, _32355_, _09107_);
  or _83140_ (_32443_, _32441_, _32440_);
  and _83141_ (_32444_, _32443_, _09112_);
  and _83142_ (_32445_, _32444_, _32439_);
  and _83143_ (_32446_, _30690_, _08039_);
  or _83144_ (_32447_, _32446_, _32355_);
  and _83145_ (_32448_, _32447_, _06602_);
  or _83146_ (_32449_, _32448_, _06639_);
  or _83147_ (_32450_, _32449_, _32445_);
  or _83148_ (_32451_, _32368_, _07048_);
  and _83149_ (_32452_, _32451_, _05990_);
  and _83150_ (_32454_, _32452_, _32450_);
  and _83151_ (_32455_, _32364_, _05989_);
  or _83152_ (_32456_, _32455_, _06646_);
  or _83153_ (_32457_, _32456_, _32454_);
  and _83154_ (_32458_, _30830_, _08039_);
  or _83155_ (_32459_, _32355_, _06651_);
  or _83156_ (_32460_, _32459_, _32458_);
  and _83157_ (_32461_, _32460_, _01442_);
  and _83158_ (_32462_, _32461_, _32457_);
  or _83159_ (_44245_, _32462_, _32353_);
  nor _83160_ (_32464_, \oc8051_golden_model_1.P0 [5], rst);
  nor _83161_ (_32465_, _32464_, _00000_);
  and _83162_ (_32466_, _13482_, \oc8051_golden_model_1.P0 [5]);
  and _83163_ (_32467_, _30842_, _08039_);
  or _83164_ (_32468_, _32467_, _32466_);
  and _83165_ (_32469_, _32468_, _06615_);
  and _83166_ (_32470_, _30848_, _08039_);
  or _83167_ (_32471_, _32470_, _32466_);
  or _83168_ (_32472_, _32471_, _07275_);
  and _83169_ (_32473_, _08039_, \oc8051_golden_model_1.ACC [5]);
  or _83170_ (_32475_, _32473_, _32466_);
  and _83171_ (_32476_, _32475_, _07259_);
  and _83172_ (_32477_, _07260_, \oc8051_golden_model_1.P0 [5]);
  or _83173_ (_32478_, _32477_, _06474_);
  or _83174_ (_32479_, _32478_, _32476_);
  and _83175_ (_32480_, _32479_, _06357_);
  and _83176_ (_32481_, _32480_, _32472_);
  and _83177_ (_32482_, _13490_, \oc8051_golden_model_1.P0 [5]);
  and _83178_ (_32483_, _30873_, _07993_);
  or _83179_ (_32484_, _32483_, _32482_);
  and _83180_ (_32486_, _32484_, _06356_);
  or _83181_ (_32487_, _32486_, _06410_);
  or _83182_ (_32488_, _32487_, _32481_);
  nor _83183_ (_32489_, _08305_, _13482_);
  or _83184_ (_32490_, _32489_, _32466_);
  or _83185_ (_32491_, _32490_, _06772_);
  and _83186_ (_32492_, _32491_, _32488_);
  or _83187_ (_32493_, _32492_, _06417_);
  or _83188_ (_32494_, _32475_, _06426_);
  and _83189_ (_32495_, _32494_, _06353_);
  and _83190_ (_32497_, _32495_, _32493_);
  and _83191_ (_32498_, _30888_, _07993_);
  or _83192_ (_32499_, _32498_, _32482_);
  and _83193_ (_32500_, _32499_, _06352_);
  or _83194_ (_32501_, _32500_, _06345_);
  or _83195_ (_32502_, _32501_, _32497_);
  or _83196_ (_32503_, _32482_, _30895_);
  and _83197_ (_32504_, _32503_, _32484_);
  or _83198_ (_32505_, _32504_, _06346_);
  and _83199_ (_32506_, _32505_, _06340_);
  and _83200_ (_32508_, _32506_, _32502_);
  and _83201_ (_32509_, _30902_, _07993_);
  or _83202_ (_32510_, _32509_, _32482_);
  and _83203_ (_32511_, _32510_, _06339_);
  or _83204_ (_32512_, _32511_, _10153_);
  or _83205_ (_32513_, _32512_, _32508_);
  or _83206_ (_32514_, _32490_, _06327_);
  and _83207_ (_32515_, _32514_, _32513_);
  or _83208_ (_32516_, _32515_, _09572_);
  and _83209_ (_32517_, _09218_, _08039_);
  or _83210_ (_32519_, _32466_, _06333_);
  or _83211_ (_32520_, _32519_, _32517_);
  and _83212_ (_32521_, _32520_, _06313_);
  and _83213_ (_32522_, _32521_, _32516_);
  and _83214_ (_32523_, _30928_, _08039_);
  or _83215_ (_32524_, _32523_, _32466_);
  and _83216_ (_32525_, _32524_, _06037_);
  or _83217_ (_32526_, _32525_, _06277_);
  or _83218_ (_32527_, _32526_, _32522_);
  and _83219_ (_32528_, _08954_, _08039_);
  or _83220_ (_32530_, _32528_, _32466_);
  or _83221_ (_32531_, _32530_, _06278_);
  and _83222_ (_32532_, _32531_, _32527_);
  or _83223_ (_32533_, _32532_, _06502_);
  and _83224_ (_32534_, _30942_, _08039_);
  or _83225_ (_32535_, _32466_, _07334_);
  or _83226_ (_32536_, _32535_, _32534_);
  and _83227_ (_32537_, _32536_, _07337_);
  and _83228_ (_32538_, _32537_, _32533_);
  or _83229_ (_32539_, _32538_, _32469_);
  and _83230_ (_32541_, _32539_, _07339_);
  or _83231_ (_32542_, _32466_, _13359_);
  and _83232_ (_32543_, _32530_, _06507_);
  and _83233_ (_32544_, _32543_, _32542_);
  or _83234_ (_32545_, _32544_, _32541_);
  and _83235_ (_32546_, _32545_, _07331_);
  and _83236_ (_32547_, _32475_, _06610_);
  and _83237_ (_32548_, _32547_, _32542_);
  or _83238_ (_32549_, _32548_, _06509_);
  or _83239_ (_32550_, _32549_, _32546_);
  and _83240_ (_32552_, _30940_, _08039_);
  or _83241_ (_32553_, _32466_, _09107_);
  or _83242_ (_32554_, _32553_, _32552_);
  and _83243_ (_32555_, _32554_, _09112_);
  and _83244_ (_32556_, _32555_, _32550_);
  and _83245_ (_32557_, _30840_, _08039_);
  or _83246_ (_32558_, _32557_, _32466_);
  and _83247_ (_32559_, _32558_, _06602_);
  or _83248_ (_32560_, _32559_, _06639_);
  or _83249_ (_32561_, _32560_, _32556_);
  or _83250_ (_32562_, _32471_, _07048_);
  and _83251_ (_32563_, _32562_, _05990_);
  and _83252_ (_32564_, _32563_, _32561_);
  and _83253_ (_32565_, _32499_, _05989_);
  or _83254_ (_32566_, _32565_, _06646_);
  or _83255_ (_32567_, _32566_, _32564_);
  and _83256_ (_32568_, _30980_, _08039_);
  or _83257_ (_32569_, _32466_, _06651_);
  or _83258_ (_32570_, _32569_, _32568_);
  and _83259_ (_32571_, _32570_, _01442_);
  and _83260_ (_32573_, _32571_, _32567_);
  or _83261_ (_44246_, _32573_, _32465_);
  nor _83262_ (_32574_, \oc8051_golden_model_1.P0 [6], rst);
  nor _83263_ (_32575_, _32574_, _00000_);
  and _83264_ (_32576_, _13482_, \oc8051_golden_model_1.P0 [6]);
  and _83265_ (_32577_, _30992_, _08039_);
  or _83266_ (_32578_, _32577_, _32576_);
  and _83267_ (_32579_, _32578_, _06615_);
  nor _83268_ (_32580_, _08209_, _13482_);
  or _83269_ (_32581_, _32580_, _32576_);
  or _83270_ (_32583_, _32581_, _06327_);
  and _83271_ (_32584_, _13490_, \oc8051_golden_model_1.P0 [6]);
  and _83272_ (_32585_, _31013_, _07993_);
  or _83273_ (_32586_, _32585_, _32584_);
  and _83274_ (_32587_, _32586_, _06352_);
  and _83275_ (_32588_, _31018_, _08039_);
  or _83276_ (_32589_, _32588_, _32576_);
  or _83277_ (_32590_, _32589_, _07275_);
  and _83278_ (_32591_, _08039_, \oc8051_golden_model_1.ACC [6]);
  or _83279_ (_32592_, _32591_, _32576_);
  and _83280_ (_32594_, _32592_, _07259_);
  and _83281_ (_32595_, _07260_, \oc8051_golden_model_1.P0 [6]);
  or _83282_ (_32596_, _32595_, _06474_);
  or _83283_ (_32597_, _32596_, _32594_);
  and _83284_ (_32598_, _32597_, _06357_);
  and _83285_ (_32599_, _32598_, _32590_);
  and _83286_ (_32600_, _31032_, _07993_);
  or _83287_ (_32601_, _32600_, _32584_);
  and _83288_ (_32602_, _32601_, _06356_);
  or _83289_ (_32603_, _32602_, _06410_);
  or _83290_ (_32605_, _32603_, _32599_);
  or _83291_ (_32606_, _32581_, _06772_);
  and _83292_ (_32607_, _32606_, _32605_);
  or _83293_ (_32608_, _32607_, _06417_);
  or _83294_ (_32609_, _32592_, _06426_);
  and _83295_ (_32610_, _32609_, _06353_);
  and _83296_ (_32611_, _32610_, _32608_);
  or _83297_ (_32612_, _32611_, _32587_);
  and _83298_ (_32613_, _32612_, _06346_);
  or _83299_ (_32614_, _32584_, _31049_);
  and _83300_ (_32616_, _32601_, _06345_);
  and _83301_ (_32617_, _32616_, _32614_);
  or _83302_ (_32618_, _32617_, _32613_);
  and _83303_ (_32619_, _32618_, _06340_);
  and _83304_ (_32620_, _31055_, _07993_);
  or _83305_ (_32621_, _32620_, _32584_);
  and _83306_ (_32622_, _32621_, _06339_);
  or _83307_ (_32623_, _32622_, _10153_);
  or _83308_ (_32624_, _32623_, _32619_);
  and _83309_ (_32625_, _32624_, _32583_);
  or _83310_ (_32627_, _32625_, _09572_);
  and _83311_ (_32628_, _09172_, _08039_);
  or _83312_ (_32629_, _32576_, _06333_);
  or _83313_ (_32630_, _32629_, _32628_);
  and _83314_ (_32631_, _32630_, _06313_);
  and _83315_ (_32632_, _32631_, _32627_);
  and _83316_ (_32633_, _31082_, _08039_);
  or _83317_ (_32634_, _32633_, _32576_);
  and _83318_ (_32635_, _32634_, _06037_);
  or _83319_ (_32636_, _32635_, _06277_);
  or _83320_ (_32638_, _32636_, _32632_);
  and _83321_ (_32639_, _15853_, _08039_);
  or _83322_ (_32640_, _32639_, _32576_);
  or _83323_ (_32641_, _32640_, _06278_);
  and _83324_ (_32642_, _32641_, _32638_);
  or _83325_ (_32643_, _32642_, _06502_);
  and _83326_ (_32644_, _31096_, _08039_);
  or _83327_ (_32645_, _32576_, _07334_);
  or _83328_ (_32646_, _32645_, _32644_);
  and _83329_ (_32647_, _32646_, _07337_);
  and _83330_ (_32649_, _32647_, _32643_);
  or _83331_ (_32650_, _32649_, _32579_);
  and _83332_ (_32651_, _32650_, _07339_);
  or _83333_ (_32652_, _32576_, _13358_);
  and _83334_ (_32653_, _32640_, _06507_);
  and _83335_ (_32654_, _32653_, _32652_);
  or _83336_ (_32655_, _32654_, _32651_);
  and _83337_ (_32656_, _32655_, _07331_);
  and _83338_ (_32657_, _32592_, _06610_);
  and _83339_ (_32658_, _32657_, _32652_);
  or _83340_ (_32660_, _32658_, _06509_);
  or _83341_ (_32661_, _32660_, _32656_);
  and _83342_ (_32662_, _31094_, _08039_);
  or _83343_ (_32663_, _32576_, _09107_);
  or _83344_ (_32664_, _32663_, _32662_);
  and _83345_ (_32665_, _32664_, _09112_);
  and _83346_ (_32666_, _32665_, _32661_);
  and _83347_ (_32667_, _30990_, _08039_);
  or _83348_ (_32668_, _32667_, _32576_);
  and _83349_ (_32669_, _32668_, _06602_);
  or _83350_ (_32671_, _32669_, _06639_);
  or _83351_ (_32672_, _32671_, _32666_);
  or _83352_ (_32673_, _32589_, _07048_);
  and _83353_ (_32674_, _32673_, _05990_);
  and _83354_ (_32675_, _32674_, _32672_);
  and _83355_ (_32676_, _32586_, _05989_);
  or _83356_ (_32677_, _32676_, _06646_);
  or _83357_ (_32678_, _32677_, _32675_);
  and _83358_ (_32679_, _31133_, _08039_);
  or _83359_ (_32680_, _32576_, _06651_);
  or _83360_ (_32682_, _32680_, _32679_);
  and _83361_ (_32683_, _32682_, _01442_);
  and _83362_ (_32684_, _32683_, _32678_);
  or _83363_ (_44247_, _32684_, _32575_);
  nor _83364_ (_32685_, \oc8051_golden_model_1.P1 [0], rst);
  nor _83365_ (_32686_, _32685_, _00000_);
  and _83366_ (_32687_, _13585_, \oc8051_golden_model_1.P1 [0]);
  and _83367_ (_32688_, _30107_, _08029_);
  or _83368_ (_32689_, _32688_, _32687_);
  and _83369_ (_32690_, _32689_, _06615_);
  and _83370_ (_32692_, _13248_, _08029_);
  or _83371_ (_32693_, _32692_, _32687_);
  or _83372_ (_32694_, _32693_, _07275_);
  and _83373_ (_32695_, _08029_, \oc8051_golden_model_1.ACC [0]);
  or _83374_ (_32696_, _32695_, _32687_);
  and _83375_ (_32697_, _32696_, _07259_);
  and _83376_ (_32698_, _07260_, \oc8051_golden_model_1.P1 [0]);
  or _83377_ (_32699_, _32698_, _06474_);
  or _83378_ (_32700_, _32699_, _32697_);
  and _83379_ (_32701_, _32700_, _06357_);
  and _83380_ (_32703_, _32701_, _32694_);
  and _83381_ (_32704_, _13593_, \oc8051_golden_model_1.P1 [0]);
  and _83382_ (_32705_, _30137_, _08661_);
  or _83383_ (_32706_, _32705_, _32704_);
  and _83384_ (_32707_, _32706_, _06356_);
  or _83385_ (_32708_, _32707_, _32703_);
  and _83386_ (_32709_, _32708_, _06772_);
  and _83387_ (_32710_, _08029_, _07250_);
  or _83388_ (_32711_, _32710_, _32687_);
  and _83389_ (_32712_, _32711_, _06410_);
  or _83390_ (_32714_, _32712_, _06417_);
  or _83391_ (_32715_, _32714_, _32709_);
  or _83392_ (_32716_, _32696_, _06426_);
  and _83393_ (_32717_, _32716_, _06353_);
  and _83394_ (_32718_, _32717_, _32715_);
  and _83395_ (_32719_, _32687_, _06352_);
  or _83396_ (_32720_, _32719_, _06345_);
  or _83397_ (_32721_, _32720_, _32718_);
  or _83398_ (_32722_, _32693_, _06346_);
  and _83399_ (_32723_, _32722_, _06340_);
  and _83400_ (_32725_, _32723_, _32721_);
  or _83401_ (_32726_, _32704_, _16663_);
  and _83402_ (_32727_, _32726_, _06339_);
  and _83403_ (_32728_, _32727_, _32706_);
  or _83404_ (_32729_, _32728_, _10153_);
  or _83405_ (_32730_, _32729_, _32725_);
  or _83406_ (_32731_, _32711_, _06327_);
  and _83407_ (_32732_, _32731_, _32730_);
  or _83408_ (_32733_, _32732_, _09572_);
  and _83409_ (_32734_, _09447_, _08029_);
  or _83410_ (_32736_, _32687_, _06333_);
  or _83411_ (_32737_, _32736_, _32734_);
  and _83412_ (_32738_, _32737_, _06313_);
  and _83413_ (_32739_, _32738_, _32733_);
  and _83414_ (_32740_, _30185_, _08029_);
  or _83415_ (_32741_, _32740_, _32687_);
  and _83416_ (_32742_, _32741_, _06037_);
  or _83417_ (_32743_, _32742_, _06277_);
  or _83418_ (_32744_, _32743_, _32739_);
  and _83419_ (_32745_, _08029_, _09008_);
  or _83420_ (_32747_, _32745_, _32687_);
  or _83421_ (_32748_, _32747_, _06278_);
  and _83422_ (_32749_, _32748_, _32744_);
  or _83423_ (_32750_, _32749_, _06502_);
  and _83424_ (_32751_, _30198_, _08029_);
  or _83425_ (_32752_, _32687_, _07334_);
  or _83426_ (_32753_, _32752_, _32751_);
  and _83427_ (_32754_, _32753_, _07337_);
  and _83428_ (_32755_, _32754_, _32750_);
  or _83429_ (_32756_, _32755_, _32690_);
  and _83430_ (_32758_, _32756_, _07339_);
  nand _83431_ (_32759_, _32747_, _06507_);
  nor _83432_ (_32760_, _32759_, _32692_);
  or _83433_ (_32761_, _32760_, _32758_);
  and _83434_ (_32762_, _32761_, _07331_);
  or _83435_ (_32763_, _32687_, _30209_);
  and _83436_ (_32764_, _32696_, _06610_);
  and _83437_ (_32765_, _32764_, _32763_);
  or _83438_ (_32766_, _32765_, _06509_);
  or _83439_ (_32767_, _32766_, _32762_);
  and _83440_ (_32769_, _30197_, _08029_);
  or _83441_ (_32770_, _32687_, _09107_);
  or _83442_ (_32771_, _32770_, _32769_);
  and _83443_ (_32772_, _32771_, _09112_);
  and _83444_ (_32773_, _32772_, _32767_);
  and _83445_ (_32774_, _30105_, _08029_);
  or _83446_ (_32775_, _32774_, _32687_);
  and _83447_ (_32776_, _32775_, _06602_);
  or _83448_ (_32777_, _32776_, _06639_);
  or _83449_ (_32778_, _32777_, _32773_);
  or _83450_ (_32780_, _32693_, _07048_);
  and _83451_ (_32781_, _32780_, _05990_);
  and _83452_ (_32782_, _32781_, _32778_);
  and _83453_ (_32783_, _32687_, _05989_);
  or _83454_ (_32784_, _32783_, _06646_);
  or _83455_ (_32785_, _32784_, _32782_);
  or _83456_ (_32786_, _32693_, _06651_);
  and _83457_ (_32787_, _32786_, _01442_);
  and _83458_ (_32788_, _32787_, _32785_);
  or _83459_ (_44249_, _32788_, _32686_);
  nor _83460_ (_32790_, \oc8051_golden_model_1.P1 [1], rst);
  nor _83461_ (_32791_, _32790_, _00000_);
  nand _83462_ (_32792_, _08029_, _07160_);
  or _83463_ (_32793_, _08029_, \oc8051_golden_model_1.P1 [1]);
  and _83464_ (_32794_, _32793_, _06277_);
  and _83465_ (_32795_, _32794_, _32792_);
  and _83466_ (_32796_, _13585_, \oc8051_golden_model_1.P1 [1]);
  nor _83467_ (_32797_, _13585_, _07448_);
  or _83468_ (_32798_, _32797_, _32796_);
  or _83469_ (_32799_, _32798_, _06772_);
  and _83470_ (_32801_, _30245_, _08029_);
  not _83471_ (_32802_, _32801_);
  and _83472_ (_32803_, _32802_, _32793_);
  or _83473_ (_32804_, _32803_, _07275_);
  nand _83474_ (_32805_, _08029_, _06097_);
  and _83475_ (_32806_, _32805_, _32793_);
  and _83476_ (_32807_, _32806_, _07259_);
  and _83477_ (_32808_, _07260_, \oc8051_golden_model_1.P1 [1]);
  or _83478_ (_32809_, _32808_, _06474_);
  or _83479_ (_32810_, _32809_, _32807_);
  and _83480_ (_32812_, _32810_, _06357_);
  and _83481_ (_32813_, _32812_, _32804_);
  and _83482_ (_32814_, _13593_, \oc8051_golden_model_1.P1 [1]);
  and _83483_ (_32815_, _30272_, _08661_);
  or _83484_ (_32816_, _32815_, _32814_);
  and _83485_ (_32817_, _32816_, _06356_);
  or _83486_ (_32818_, _32817_, _06410_);
  or _83487_ (_32819_, _32818_, _32813_);
  and _83488_ (_32820_, _32819_, _32799_);
  or _83489_ (_32821_, _32820_, _06417_);
  or _83490_ (_32823_, _32806_, _06426_);
  and _83491_ (_32824_, _32823_, _06353_);
  and _83492_ (_32825_, _32824_, _32821_);
  and _83493_ (_32826_, _30283_, _08661_);
  or _83494_ (_32827_, _32826_, _32814_);
  and _83495_ (_32828_, _32827_, _06352_);
  or _83496_ (_32829_, _32828_, _06345_);
  or _83497_ (_32830_, _32829_, _32825_);
  and _83498_ (_32831_, _32815_, _30291_);
  or _83499_ (_32832_, _32814_, _06346_);
  or _83500_ (_32834_, _32832_, _32831_);
  and _83501_ (_32835_, _32834_, _32830_);
  and _83502_ (_32836_, _32835_, _06340_);
  and _83503_ (_32837_, _30297_, _08661_);
  or _83504_ (_32838_, _32814_, _32837_);
  and _83505_ (_32839_, _32838_, _06339_);
  or _83506_ (_32840_, _32839_, _10153_);
  or _83507_ (_32841_, _32840_, _32836_);
  or _83508_ (_32842_, _32798_, _06327_);
  and _83509_ (_32843_, _32842_, _32841_);
  or _83510_ (_32845_, _32843_, _09572_);
  and _83511_ (_32846_, _09402_, _08029_);
  or _83512_ (_32847_, _32796_, _06333_);
  or _83513_ (_32848_, _32847_, _32846_);
  and _83514_ (_32849_, _32848_, _06313_);
  and _83515_ (_32850_, _32849_, _32845_);
  and _83516_ (_32851_, _30325_, _08029_);
  or _83517_ (_32852_, _32851_, _32796_);
  and _83518_ (_32853_, _32852_, _06037_);
  or _83519_ (_32854_, _32853_, _32850_);
  and _83520_ (_32856_, _32854_, _06278_);
  or _83521_ (_32857_, _32856_, _32795_);
  and _83522_ (_32858_, _32857_, _07334_);
  or _83523_ (_32859_, _30339_, _13585_);
  and _83524_ (_32860_, _32793_, _06502_);
  and _83525_ (_32861_, _32860_, _32859_);
  or _83526_ (_32862_, _32861_, _32858_);
  and _83527_ (_32863_, _32862_, _07337_);
  or _83528_ (_32864_, _30348_, _13585_);
  and _83529_ (_32865_, _32793_, _06615_);
  and _83530_ (_32867_, _32865_, _32864_);
  or _83531_ (_32868_, _32867_, _32863_);
  and _83532_ (_32869_, _32868_, _07339_);
  or _83533_ (_32870_, _30337_, _13585_);
  and _83534_ (_32871_, _32793_, _06507_);
  and _83535_ (_32872_, _32871_, _32870_);
  or _83536_ (_32873_, _32872_, _32869_);
  and _83537_ (_32874_, _32873_, _07331_);
  or _83538_ (_32875_, _32796_, _30360_);
  and _83539_ (_32876_, _32806_, _06610_);
  and _83540_ (_32878_, _32876_, _32875_);
  or _83541_ (_32879_, _32878_, _32874_);
  and _83542_ (_32880_, _32879_, _06603_);
  or _83543_ (_32881_, _32805_, _30360_);
  and _83544_ (_32882_, _32793_, _06602_);
  and _83545_ (_32883_, _32882_, _32881_);
  or _83546_ (_32884_, _32883_, _06639_);
  or _83547_ (_32885_, _32792_, _30360_);
  and _83548_ (_32886_, _32793_, _06509_);
  and _83549_ (_32887_, _32886_, _32885_);
  or _83550_ (_32889_, _32887_, _32884_);
  or _83551_ (_32890_, _32889_, _32880_);
  or _83552_ (_32891_, _32803_, _07048_);
  and _83553_ (_32892_, _32891_, _05990_);
  and _83554_ (_32893_, _32892_, _32890_);
  and _83555_ (_32894_, _32827_, _05989_);
  or _83556_ (_32895_, _32894_, _06646_);
  or _83557_ (_32896_, _32895_, _32893_);
  or _83558_ (_32897_, _32796_, _06651_);
  or _83559_ (_32898_, _32897_, _32801_);
  and _83560_ (_32900_, _32898_, _01442_);
  and _83561_ (_32901_, _32900_, _32896_);
  or _83562_ (_44250_, _32901_, _32791_);
  nor _83563_ (_32902_, \oc8051_golden_model_1.P1 [2], rst);
  nor _83564_ (_32903_, _32902_, _00000_);
  and _83565_ (_32904_, _13585_, \oc8051_golden_model_1.P1 [2]);
  and _83566_ (_32905_, _30393_, _08029_);
  or _83567_ (_32906_, _32905_, _32904_);
  and _83568_ (_32907_, _32906_, _06615_);
  nor _83569_ (_32908_, _13585_, _07854_);
  or _83570_ (_32910_, _32908_, _32904_);
  or _83571_ (_32911_, _32910_, _06327_);
  or _83572_ (_32912_, _32910_, _06772_);
  and _83573_ (_32913_, _30403_, _08029_);
  or _83574_ (_32914_, _32913_, _32904_);
  or _83575_ (_32915_, _32914_, _07275_);
  and _83576_ (_32916_, _08029_, \oc8051_golden_model_1.ACC [2]);
  or _83577_ (_32917_, _32916_, _32904_);
  and _83578_ (_32918_, _32917_, _07259_);
  and _83579_ (_32919_, _07260_, \oc8051_golden_model_1.P1 [2]);
  or _83580_ (_32921_, _32919_, _06474_);
  or _83581_ (_32922_, _32921_, _32918_);
  and _83582_ (_32923_, _32922_, _06357_);
  and _83583_ (_32924_, _32923_, _32915_);
  and _83584_ (_32925_, _13593_, \oc8051_golden_model_1.P1 [2]);
  and _83585_ (_32926_, _30428_, _08661_);
  or _83586_ (_32927_, _32926_, _32925_);
  and _83587_ (_32928_, _32927_, _06356_);
  or _83588_ (_32929_, _32928_, _06410_);
  or _83589_ (_32930_, _32929_, _32924_);
  and _83590_ (_32932_, _32930_, _32912_);
  or _83591_ (_32933_, _32932_, _06417_);
  or _83592_ (_32934_, _32917_, _06426_);
  and _83593_ (_32935_, _32934_, _06353_);
  and _83594_ (_32936_, _32935_, _32933_);
  and _83595_ (_32937_, _30440_, _08661_);
  or _83596_ (_32938_, _32937_, _32925_);
  and _83597_ (_32939_, _32938_, _06352_);
  or _83598_ (_32940_, _32939_, _06345_);
  or _83599_ (_32941_, _32940_, _32936_);
  and _83600_ (_32943_, _32926_, _30447_);
  or _83601_ (_32944_, _32925_, _06346_);
  or _83602_ (_32945_, _32944_, _32943_);
  and _83603_ (_32946_, _32945_, _06340_);
  and _83604_ (_32947_, _32946_, _32941_);
  and _83605_ (_32948_, _30454_, _08661_);
  or _83606_ (_32949_, _32948_, _32925_);
  and _83607_ (_32950_, _32949_, _06339_);
  or _83608_ (_32951_, _32950_, _10153_);
  or _83609_ (_32952_, _32951_, _32947_);
  and _83610_ (_32954_, _32952_, _32911_);
  or _83611_ (_32955_, _32954_, _09572_);
  and _83612_ (_32956_, _09356_, _08029_);
  or _83613_ (_32957_, _32904_, _06333_);
  or _83614_ (_32958_, _32957_, _32956_);
  and _83615_ (_32959_, _32958_, _06313_);
  and _83616_ (_32960_, _32959_, _32955_);
  and _83617_ (_32961_, _30479_, _08029_);
  or _83618_ (_32962_, _32961_, _32904_);
  and _83619_ (_32963_, _32962_, _06037_);
  or _83620_ (_32965_, _32963_, _06277_);
  or _83621_ (_32966_, _32965_, _32960_);
  and _83622_ (_32967_, _08029_, _09057_);
  or _83623_ (_32968_, _32967_, _32904_);
  or _83624_ (_32969_, _32968_, _06278_);
  and _83625_ (_32970_, _32969_, _32966_);
  or _83626_ (_32971_, _32970_, _06502_);
  and _83627_ (_32972_, _30493_, _08029_);
  or _83628_ (_32973_, _32904_, _07334_);
  or _83629_ (_32974_, _32973_, _32972_);
  and _83630_ (_32976_, _32974_, _07337_);
  and _83631_ (_32977_, _32976_, _32971_);
  or _83632_ (_32978_, _32977_, _32907_);
  and _83633_ (_32979_, _32978_, _07339_);
  or _83634_ (_32980_, _32904_, _13362_);
  and _83635_ (_32981_, _32968_, _06507_);
  and _83636_ (_32982_, _32981_, _32980_);
  or _83637_ (_32983_, _32982_, _32979_);
  and _83638_ (_32984_, _32983_, _07331_);
  and _83639_ (_32985_, _32917_, _06610_);
  and _83640_ (_32987_, _32985_, _32980_);
  or _83641_ (_32988_, _32987_, _06509_);
  or _83642_ (_32989_, _32988_, _32984_);
  and _83643_ (_32990_, _30491_, _08029_);
  or _83644_ (_32991_, _32904_, _09107_);
  or _83645_ (_32992_, _32991_, _32990_);
  and _83646_ (_32993_, _32992_, _09112_);
  and _83647_ (_32994_, _32993_, _32989_);
  and _83648_ (_32995_, _30391_, _08029_);
  or _83649_ (_32996_, _32995_, _32904_);
  and _83650_ (_32998_, _32996_, _06602_);
  or _83651_ (_32999_, _32998_, _06639_);
  or _83652_ (_33000_, _32999_, _32994_);
  or _83653_ (_33001_, _32914_, _07048_);
  and _83654_ (_33002_, _33001_, _05990_);
  and _83655_ (_33003_, _33002_, _33000_);
  and _83656_ (_33004_, _32938_, _05989_);
  or _83657_ (_33005_, _33004_, _06646_);
  or _83658_ (_33006_, _33005_, _33003_);
  and _83659_ (_33007_, _30531_, _08029_);
  or _83660_ (_33009_, _32904_, _06651_);
  or _83661_ (_33010_, _33009_, _33007_);
  and _83662_ (_33011_, _33010_, _01442_);
  and _83663_ (_33012_, _33011_, _33006_);
  or _83664_ (_44251_, _33012_, _32903_);
  nor _83665_ (_33013_, \oc8051_golden_model_1.P1 [3], rst);
  nor _83666_ (_33014_, _33013_, _00000_);
  and _83667_ (_33015_, _13585_, \oc8051_golden_model_1.P1 [3]);
  and _83668_ (_33016_, _30543_, _08029_);
  or _83669_ (_33017_, _33016_, _33015_);
  and _83670_ (_33019_, _33017_, _06615_);
  nor _83671_ (_33020_, _13585_, _07680_);
  or _83672_ (_33021_, _33020_, _33015_);
  or _83673_ (_33022_, _33021_, _06327_);
  and _83674_ (_33023_, _30552_, _08029_);
  or _83675_ (_33024_, _33023_, _33015_);
  or _83676_ (_33025_, _33024_, _07275_);
  and _83677_ (_33026_, _08029_, \oc8051_golden_model_1.ACC [3]);
  or _83678_ (_33027_, _33026_, _33015_);
  and _83679_ (_33028_, _33027_, _07259_);
  and _83680_ (_33030_, _07260_, \oc8051_golden_model_1.P1 [3]);
  or _83681_ (_33031_, _33030_, _06474_);
  or _83682_ (_33032_, _33031_, _33028_);
  and _83683_ (_33033_, _33032_, _06357_);
  and _83684_ (_33034_, _33033_, _33025_);
  and _83685_ (_33035_, _13593_, \oc8051_golden_model_1.P1 [3]);
  and _83686_ (_33036_, _30577_, _08661_);
  or _83687_ (_33037_, _33036_, _33035_);
  and _83688_ (_33038_, _33037_, _06356_);
  or _83689_ (_33039_, _33038_, _06410_);
  or _83690_ (_33041_, _33039_, _33034_);
  or _83691_ (_33042_, _33021_, _06772_);
  and _83692_ (_33043_, _33042_, _33041_);
  or _83693_ (_33044_, _33043_, _06417_);
  or _83694_ (_33045_, _33027_, _06426_);
  and _83695_ (_33046_, _33045_, _06353_);
  and _83696_ (_33047_, _33046_, _33044_);
  and _83697_ (_33048_, _30590_, _08661_);
  or _83698_ (_33049_, _33048_, _33035_);
  and _83699_ (_33050_, _33049_, _06352_);
  or _83700_ (_33052_, _33050_, _06345_);
  or _83701_ (_33053_, _33052_, _33047_);
  or _83702_ (_33054_, _33035_, _30597_);
  and _83703_ (_33055_, _33054_, _33037_);
  or _83704_ (_33056_, _33055_, _06346_);
  and _83705_ (_33057_, _33056_, _06340_);
  and _83706_ (_33058_, _33057_, _33053_);
  and _83707_ (_33059_, _30603_, _08661_);
  or _83708_ (_33060_, _33059_, _33035_);
  and _83709_ (_33061_, _33060_, _06339_);
  or _83710_ (_33063_, _33061_, _10153_);
  or _83711_ (_33064_, _33063_, _33058_);
  and _83712_ (_33065_, _33064_, _33022_);
  or _83713_ (_33066_, _33065_, _09572_);
  and _83714_ (_33067_, _09310_, _08029_);
  or _83715_ (_33068_, _33015_, _06333_);
  or _83716_ (_33069_, _33068_, _33067_);
  and _83717_ (_33070_, _33069_, _06313_);
  and _83718_ (_33071_, _33070_, _33066_);
  and _83719_ (_33072_, _30629_, _08029_);
  or _83720_ (_33074_, _33072_, _33015_);
  and _83721_ (_33075_, _33074_, _06037_);
  or _83722_ (_33076_, _33075_, _06277_);
  or _83723_ (_33077_, _33076_, _33071_);
  and _83724_ (_33078_, _08029_, _09014_);
  or _83725_ (_33079_, _33078_, _33015_);
  or _83726_ (_33080_, _33079_, _06278_);
  and _83727_ (_33081_, _33080_, _33077_);
  or _83728_ (_33082_, _33081_, _06502_);
  and _83729_ (_33083_, _30643_, _08029_);
  or _83730_ (_33085_, _33015_, _07334_);
  or _83731_ (_33086_, _33085_, _33083_);
  and _83732_ (_33087_, _33086_, _07337_);
  and _83733_ (_33088_, _33087_, _33082_);
  or _83734_ (_33089_, _33088_, _33019_);
  and _83735_ (_33090_, _33089_, _07339_);
  or _83736_ (_33091_, _33015_, _13361_);
  and _83737_ (_33092_, _33079_, _06507_);
  and _83738_ (_33093_, _33092_, _33091_);
  or _83739_ (_33094_, _33093_, _33090_);
  and _83740_ (_33096_, _33094_, _07331_);
  and _83741_ (_33097_, _33027_, _06610_);
  and _83742_ (_33098_, _33097_, _33091_);
  or _83743_ (_33099_, _33098_, _06509_);
  or _83744_ (_33100_, _33099_, _33096_);
  and _83745_ (_33101_, _30641_, _08029_);
  or _83746_ (_33102_, _33015_, _09107_);
  or _83747_ (_33103_, _33102_, _33101_);
  and _83748_ (_33104_, _33103_, _09112_);
  and _83749_ (_33105_, _33104_, _33100_);
  and _83750_ (_33106_, _30541_, _08029_);
  or _83751_ (_33107_, _33106_, _33015_);
  and _83752_ (_33108_, _33107_, _06602_);
  or _83753_ (_33109_, _33108_, _06639_);
  or _83754_ (_33110_, _33109_, _33105_);
  or _83755_ (_33111_, _33024_, _07048_);
  and _83756_ (_33112_, _33111_, _05990_);
  and _83757_ (_33113_, _33112_, _33110_);
  and _83758_ (_33114_, _33049_, _05989_);
  or _83759_ (_33115_, _33114_, _06646_);
  or _83760_ (_33117_, _33115_, _33113_);
  and _83761_ (_33118_, _30680_, _08029_);
  or _83762_ (_33119_, _33015_, _06651_);
  or _83763_ (_33120_, _33119_, _33118_);
  and _83764_ (_33121_, _33120_, _01442_);
  and _83765_ (_33122_, _33121_, _33117_);
  or _83766_ (_44252_, _33122_, _33014_);
  nor _83767_ (_33123_, \oc8051_golden_model_1.P1 [4], rst);
  nor _83768_ (_33124_, _33123_, _00000_);
  and _83769_ (_33125_, _13585_, \oc8051_golden_model_1.P1 [4]);
  and _83770_ (_33127_, _30693_, _08029_);
  or _83771_ (_33128_, _33127_, _33125_);
  and _83772_ (_33129_, _33128_, _06615_);
  nor _83773_ (_33130_, _08596_, _13585_);
  or _83774_ (_33131_, _33130_, _33125_);
  or _83775_ (_33132_, _33131_, _06327_);
  and _83776_ (_33133_, _13593_, \oc8051_golden_model_1.P1 [4]);
  and _83777_ (_33134_, _30712_, _08661_);
  or _83778_ (_33135_, _33134_, _33133_);
  and _83779_ (_33136_, _33135_, _06352_);
  and _83780_ (_33138_, _30718_, _08029_);
  or _83781_ (_33139_, _33138_, _33125_);
  or _83782_ (_33140_, _33139_, _07275_);
  and _83783_ (_33141_, _08029_, \oc8051_golden_model_1.ACC [4]);
  or _83784_ (_33142_, _33141_, _33125_);
  and _83785_ (_33143_, _33142_, _07259_);
  and _83786_ (_33144_, _07260_, \oc8051_golden_model_1.P1 [4]);
  or _83787_ (_33145_, _33144_, _06474_);
  or _83788_ (_33146_, _33145_, _33143_);
  and _83789_ (_33147_, _33146_, _06357_);
  and _83790_ (_33149_, _33147_, _33140_);
  and _83791_ (_33150_, _30731_, _08661_);
  or _83792_ (_33151_, _33150_, _33133_);
  and _83793_ (_33152_, _33151_, _06356_);
  or _83794_ (_33153_, _33152_, _06410_);
  or _83795_ (_33154_, _33153_, _33149_);
  or _83796_ (_33155_, _33131_, _06772_);
  and _83797_ (_33156_, _33155_, _33154_);
  or _83798_ (_33157_, _33156_, _06417_);
  or _83799_ (_33158_, _33142_, _06426_);
  and _83800_ (_33160_, _33158_, _06353_);
  and _83801_ (_33161_, _33160_, _33157_);
  or _83802_ (_33162_, _33161_, _33136_);
  and _83803_ (_33163_, _33162_, _06346_);
  or _83804_ (_33164_, _33133_, _30746_);
  and _83805_ (_33165_, _33151_, _06345_);
  and _83806_ (_33166_, _33165_, _33164_);
  or _83807_ (_33167_, _33166_, _33163_);
  and _83808_ (_33168_, _33167_, _06340_);
  and _83809_ (_33169_, _30753_, _08661_);
  or _83810_ (_33171_, _33169_, _33133_);
  and _83811_ (_33172_, _33171_, _06339_);
  or _83812_ (_33173_, _33172_, _10153_);
  or _83813_ (_33174_, _33173_, _33168_);
  and _83814_ (_33175_, _33174_, _33132_);
  or _83815_ (_33176_, _33175_, _09572_);
  and _83816_ (_33177_, _09264_, _08029_);
  or _83817_ (_33178_, _33125_, _06333_);
  or _83818_ (_33179_, _33178_, _33177_);
  and _83819_ (_33180_, _33179_, _06313_);
  and _83820_ (_33182_, _33180_, _33176_);
  and _83821_ (_33183_, _30778_, _08029_);
  or _83822_ (_33184_, _33183_, _33125_);
  and _83823_ (_33185_, _33184_, _06037_);
  or _83824_ (_33186_, _33185_, _06277_);
  or _83825_ (_33187_, _33186_, _33182_);
  and _83826_ (_33188_, _08995_, _08029_);
  or _83827_ (_33189_, _33188_, _33125_);
  or _83828_ (_33190_, _33189_, _06278_);
  and _83829_ (_33191_, _33190_, _33187_);
  or _83830_ (_33193_, _33191_, _06502_);
  and _83831_ (_33194_, _30793_, _08029_);
  or _83832_ (_33195_, _33125_, _07334_);
  or _83833_ (_33196_, _33195_, _33194_);
  and _83834_ (_33197_, _33196_, _07337_);
  and _83835_ (_33198_, _33197_, _33193_);
  or _83836_ (_33199_, _33198_, _33129_);
  and _83837_ (_33200_, _33199_, _07339_);
  or _83838_ (_33201_, _33125_, _13360_);
  and _83839_ (_33202_, _33189_, _06507_);
  and _83840_ (_33204_, _33202_, _33201_);
  or _83841_ (_33205_, _33204_, _33200_);
  and _83842_ (_33206_, _33205_, _07331_);
  and _83843_ (_33207_, _33142_, _06610_);
  and _83844_ (_33208_, _33207_, _33201_);
  or _83845_ (_33209_, _33208_, _06509_);
  or _83846_ (_33210_, _33209_, _33206_);
  and _83847_ (_33211_, _30790_, _08029_);
  or _83848_ (_33212_, _33125_, _09107_);
  or _83849_ (_33213_, _33212_, _33211_);
  and _83850_ (_33215_, _33213_, _09112_);
  and _83851_ (_33216_, _33215_, _33210_);
  and _83852_ (_33217_, _30690_, _08029_);
  or _83853_ (_33218_, _33217_, _33125_);
  and _83854_ (_33219_, _33218_, _06602_);
  or _83855_ (_33220_, _33219_, _06639_);
  or _83856_ (_33221_, _33220_, _33216_);
  or _83857_ (_33222_, _33139_, _07048_);
  and _83858_ (_33223_, _33222_, _05990_);
  and _83859_ (_33224_, _33223_, _33221_);
  and _83860_ (_33226_, _33135_, _05989_);
  or _83861_ (_33227_, _33226_, _06646_);
  or _83862_ (_33228_, _33227_, _33224_);
  and _83863_ (_33229_, _30830_, _08029_);
  or _83864_ (_33230_, _33125_, _06651_);
  or _83865_ (_33231_, _33230_, _33229_);
  and _83866_ (_33232_, _33231_, _01442_);
  and _83867_ (_33233_, _33232_, _33228_);
  or _83868_ (_44253_, _33233_, _33124_);
  nor _83869_ (_33234_, \oc8051_golden_model_1.P1 [5], rst);
  nor _83870_ (_33236_, _33234_, _00000_);
  and _83871_ (_33237_, _13585_, \oc8051_golden_model_1.P1 [5]);
  and _83872_ (_33238_, _30842_, _08029_);
  or _83873_ (_33239_, _33238_, _33237_);
  and _83874_ (_33240_, _33239_, _06615_);
  and _83875_ (_33241_, _30848_, _08029_);
  or _83876_ (_33242_, _33241_, _33237_);
  or _83877_ (_33243_, _33242_, _07275_);
  and _83878_ (_33244_, _08029_, \oc8051_golden_model_1.ACC [5]);
  or _83879_ (_33245_, _33244_, _33237_);
  and _83880_ (_33247_, _33245_, _07259_);
  and _83881_ (_33248_, _07260_, \oc8051_golden_model_1.P1 [5]);
  or _83882_ (_33249_, _33248_, _06474_);
  or _83883_ (_33250_, _33249_, _33247_);
  and _83884_ (_33251_, _33250_, _06357_);
  and _83885_ (_33252_, _33251_, _33243_);
  and _83886_ (_33253_, _13593_, \oc8051_golden_model_1.P1 [5]);
  and _83887_ (_33254_, _30873_, _08661_);
  or _83888_ (_33255_, _33254_, _33253_);
  and _83889_ (_33256_, _33255_, _06356_);
  or _83890_ (_33258_, _33256_, _06410_);
  or _83891_ (_33259_, _33258_, _33252_);
  nor _83892_ (_33260_, _08305_, _13585_);
  or _83893_ (_33261_, _33260_, _33237_);
  or _83894_ (_33262_, _33261_, _06772_);
  and _83895_ (_33263_, _33262_, _33259_);
  or _83896_ (_33264_, _33263_, _06417_);
  or _83897_ (_33265_, _33245_, _06426_);
  and _83898_ (_33266_, _33265_, _06353_);
  and _83899_ (_33267_, _33266_, _33264_);
  and _83900_ (_33269_, _30888_, _08661_);
  or _83901_ (_33270_, _33269_, _33253_);
  and _83902_ (_33271_, _33270_, _06352_);
  or _83903_ (_33272_, _33271_, _06345_);
  or _83904_ (_33273_, _33272_, _33267_);
  or _83905_ (_33274_, _33253_, _30895_);
  and _83906_ (_33275_, _33274_, _33255_);
  or _83907_ (_33276_, _33275_, _06346_);
  and _83908_ (_33277_, _33276_, _06340_);
  and _83909_ (_33278_, _33277_, _33273_);
  and _83910_ (_33280_, _30902_, _08661_);
  or _83911_ (_33281_, _33280_, _33253_);
  and _83912_ (_33282_, _33281_, _06339_);
  or _83913_ (_33283_, _33282_, _10153_);
  or _83914_ (_33284_, _33283_, _33278_);
  or _83915_ (_33285_, _33261_, _06327_);
  and _83916_ (_33286_, _33285_, _33284_);
  or _83917_ (_33287_, _33286_, _09572_);
  and _83918_ (_33288_, _09218_, _08029_);
  or _83919_ (_33289_, _33237_, _06333_);
  or _83920_ (_33291_, _33289_, _33288_);
  and _83921_ (_33292_, _33291_, _06313_);
  and _83922_ (_33293_, _33292_, _33287_);
  and _83923_ (_33294_, _30928_, _08029_);
  or _83924_ (_33295_, _33294_, _33237_);
  and _83925_ (_33296_, _33295_, _06037_);
  or _83926_ (_33297_, _33296_, _06277_);
  or _83927_ (_33298_, _33297_, _33293_);
  and _83928_ (_33299_, _08954_, _08029_);
  or _83929_ (_33300_, _33299_, _33237_);
  or _83930_ (_33302_, _33300_, _06278_);
  and _83931_ (_33303_, _33302_, _33298_);
  or _83932_ (_33304_, _33303_, _06502_);
  and _83933_ (_33305_, _30942_, _08029_);
  or _83934_ (_33306_, _33237_, _07334_);
  or _83935_ (_33307_, _33306_, _33305_);
  and _83936_ (_33308_, _33307_, _07337_);
  and _83937_ (_33309_, _33308_, _33304_);
  or _83938_ (_33310_, _33309_, _33240_);
  and _83939_ (_33311_, _33310_, _07339_);
  or _83940_ (_33313_, _33237_, _13359_);
  and _83941_ (_33314_, _33300_, _06507_);
  and _83942_ (_33315_, _33314_, _33313_);
  or _83943_ (_33316_, _33315_, _33311_);
  and _83944_ (_33317_, _33316_, _07331_);
  and _83945_ (_33318_, _33245_, _06610_);
  and _83946_ (_33319_, _33318_, _33313_);
  or _83947_ (_33320_, _33319_, _06509_);
  or _83948_ (_33321_, _33320_, _33317_);
  and _83949_ (_33322_, _30940_, _08029_);
  or _83950_ (_33324_, _33237_, _09107_);
  or _83951_ (_33325_, _33324_, _33322_);
  and _83952_ (_33326_, _33325_, _09112_);
  and _83953_ (_33327_, _33326_, _33321_);
  and _83954_ (_33328_, _30840_, _08029_);
  or _83955_ (_33329_, _33328_, _33237_);
  and _83956_ (_33330_, _33329_, _06602_);
  or _83957_ (_33331_, _33330_, _06639_);
  or _83958_ (_33332_, _33331_, _33327_);
  or _83959_ (_33333_, _33242_, _07048_);
  and _83960_ (_33335_, _33333_, _05990_);
  and _83961_ (_33336_, _33335_, _33332_);
  and _83962_ (_33337_, _33270_, _05989_);
  or _83963_ (_33338_, _33337_, _06646_);
  or _83964_ (_33339_, _33338_, _33336_);
  and _83965_ (_33340_, _30980_, _08029_);
  or _83966_ (_33341_, _33237_, _06651_);
  or _83967_ (_33342_, _33341_, _33340_);
  and _83968_ (_33343_, _33342_, _01442_);
  and _83969_ (_33344_, _33343_, _33339_);
  or _83970_ (_44254_, _33344_, _33236_);
  nor _83971_ (_33346_, \oc8051_golden_model_1.P1 [6], rst);
  nor _83972_ (_33347_, _33346_, _00000_);
  and _83973_ (_33348_, _13585_, \oc8051_golden_model_1.P1 [6]);
  and _83974_ (_33349_, _30992_, _08029_);
  or _83975_ (_33350_, _33349_, _33348_);
  and _83976_ (_33351_, _33350_, _06615_);
  nor _83977_ (_33352_, _08209_, _13585_);
  or _83978_ (_33353_, _33352_, _33348_);
  or _83979_ (_33354_, _33353_, _06327_);
  and _83980_ (_33356_, _13593_, \oc8051_golden_model_1.P1 [6]);
  and _83981_ (_33357_, _31013_, _08661_);
  or _83982_ (_33358_, _33357_, _33356_);
  and _83983_ (_33359_, _33358_, _06352_);
  and _83984_ (_33360_, _31018_, _08029_);
  or _83985_ (_33361_, _33360_, _33348_);
  or _83986_ (_33362_, _33361_, _07275_);
  and _83987_ (_33363_, _08029_, \oc8051_golden_model_1.ACC [6]);
  or _83988_ (_33364_, _33363_, _33348_);
  and _83989_ (_33365_, _33364_, _07259_);
  and _83990_ (_33367_, _07260_, \oc8051_golden_model_1.P1 [6]);
  or _83991_ (_33368_, _33367_, _06474_);
  or _83992_ (_33369_, _33368_, _33365_);
  and _83993_ (_33370_, _33369_, _06357_);
  and _83994_ (_33371_, _33370_, _33362_);
  and _83995_ (_33372_, _31032_, _08661_);
  or _83996_ (_33373_, _33372_, _33356_);
  and _83997_ (_33374_, _33373_, _06356_);
  or _83998_ (_33375_, _33374_, _06410_);
  or _83999_ (_33376_, _33375_, _33371_);
  or _84000_ (_33378_, _33353_, _06772_);
  and _84001_ (_33379_, _33378_, _33376_);
  or _84002_ (_33380_, _33379_, _06417_);
  or _84003_ (_33381_, _33364_, _06426_);
  and _84004_ (_33382_, _33381_, _06353_);
  and _84005_ (_33383_, _33382_, _33380_);
  or _84006_ (_33384_, _33383_, _33359_);
  and _84007_ (_33385_, _33384_, _06346_);
  or _84008_ (_33386_, _33356_, _31049_);
  and _84009_ (_33387_, _33373_, _06345_);
  and _84010_ (_33389_, _33387_, _33386_);
  or _84011_ (_33390_, _33389_, _33385_);
  and _84012_ (_33391_, _33390_, _06340_);
  and _84013_ (_33392_, _31055_, _08661_);
  or _84014_ (_33393_, _33392_, _33356_);
  and _84015_ (_33394_, _33393_, _06339_);
  or _84016_ (_33395_, _33394_, _10153_);
  or _84017_ (_33396_, _33395_, _33391_);
  and _84018_ (_33397_, _33396_, _33354_);
  or _84019_ (_33398_, _33397_, _09572_);
  and _84020_ (_33400_, _09172_, _08029_);
  or _84021_ (_33401_, _33348_, _06333_);
  or _84022_ (_33402_, _33401_, _33400_);
  and _84023_ (_33403_, _33402_, _06313_);
  and _84024_ (_33404_, _33403_, _33398_);
  and _84025_ (_33405_, _31082_, _08029_);
  or _84026_ (_33406_, _33405_, _33348_);
  and _84027_ (_33407_, _33406_, _06037_);
  or _84028_ (_33408_, _33407_, _06277_);
  or _84029_ (_33409_, _33408_, _33404_);
  and _84030_ (_33411_, _15853_, _08029_);
  or _84031_ (_33412_, _33411_, _33348_);
  or _84032_ (_33413_, _33412_, _06278_);
  and _84033_ (_33414_, _33413_, _33409_);
  or _84034_ (_33415_, _33414_, _06502_);
  and _84035_ (_33416_, _31096_, _08029_);
  or _84036_ (_33417_, _33348_, _07334_);
  or _84037_ (_33418_, _33417_, _33416_);
  and _84038_ (_33419_, _33418_, _07337_);
  and _84039_ (_33420_, _33419_, _33415_);
  or _84040_ (_33422_, _33420_, _33351_);
  and _84041_ (_33423_, _33422_, _07339_);
  or _84042_ (_33424_, _33348_, _13358_);
  and _84043_ (_33425_, _33412_, _06507_);
  and _84044_ (_33426_, _33425_, _33424_);
  or _84045_ (_33427_, _33426_, _33423_);
  and _84046_ (_33428_, _33427_, _07331_);
  and _84047_ (_33429_, _33364_, _06610_);
  and _84048_ (_33430_, _33429_, _33424_);
  or _84049_ (_33431_, _33430_, _06509_);
  or _84050_ (_33433_, _33431_, _33428_);
  and _84051_ (_33434_, _31094_, _08029_);
  or _84052_ (_33435_, _33348_, _09107_);
  or _84053_ (_33436_, _33435_, _33434_);
  and _84054_ (_33437_, _33436_, _09112_);
  and _84055_ (_33438_, _33437_, _33433_);
  and _84056_ (_33439_, _30990_, _08029_);
  or _84057_ (_33440_, _33439_, _33348_);
  and _84058_ (_33441_, _33440_, _06602_);
  or _84059_ (_33442_, _33441_, _06639_);
  or _84060_ (_33444_, _33442_, _33438_);
  or _84061_ (_33445_, _33361_, _07048_);
  and _84062_ (_33446_, _33445_, _05990_);
  and _84063_ (_33447_, _33446_, _33444_);
  and _84064_ (_33448_, _33358_, _05989_);
  or _84065_ (_33449_, _33448_, _06646_);
  or _84066_ (_33450_, _33449_, _33447_);
  and _84067_ (_33451_, _31133_, _08029_);
  or _84068_ (_33452_, _33348_, _06651_);
  or _84069_ (_33453_, _33452_, _33451_);
  and _84070_ (_33455_, _33453_, _01442_);
  and _84071_ (_33456_, _33455_, _33450_);
  or _84072_ (_44255_, _33456_, _33347_);
  and _84073_ (_33457_, _01446_, \oc8051_golden_model_1.IP [0]);
  and _84074_ (_33458_, _13693_, \oc8051_golden_model_1.IP [0]);
  nor _84075_ (_33459_, _12622_, _13693_);
  or _84076_ (_33460_, _33459_, _33458_);
  and _84077_ (_33461_, _10577_, _08022_);
  nor _84078_ (_33462_, _33461_, _07337_);
  and _84079_ (_33463_, _33462_, _33460_);
  nor _84080_ (_33465_, _08453_, _13693_);
  or _84081_ (_33466_, _33465_, _33458_);
  or _84082_ (_33467_, _33466_, _07275_);
  and _84083_ (_33468_, _08022_, \oc8051_golden_model_1.ACC [0]);
  or _84084_ (_33469_, _33468_, _33458_);
  and _84085_ (_33470_, _33469_, _07259_);
  and _84086_ (_33471_, _07260_, \oc8051_golden_model_1.IP [0]);
  or _84087_ (_33472_, _33471_, _06474_);
  or _84088_ (_33473_, _33472_, _33470_);
  and _84089_ (_33474_, _33473_, _06357_);
  and _84090_ (_33476_, _33474_, _33467_);
  and _84091_ (_33477_, _13701_, \oc8051_golden_model_1.IP [0]);
  and _84092_ (_33478_, _14581_, _08643_);
  or _84093_ (_33479_, _33478_, _33477_);
  and _84094_ (_33480_, _33479_, _06356_);
  or _84095_ (_33481_, _33480_, _33476_);
  and _84096_ (_33482_, _33481_, _06772_);
  and _84097_ (_33483_, _08022_, _07250_);
  or _84098_ (_33484_, _33483_, _33458_);
  and _84099_ (_33485_, _33484_, _06410_);
  or _84100_ (_33487_, _33485_, _06417_);
  or _84101_ (_33488_, _33487_, _33482_);
  or _84102_ (_33489_, _33469_, _06426_);
  and _84103_ (_33490_, _33489_, _06353_);
  and _84104_ (_33491_, _33490_, _33488_);
  and _84105_ (_33492_, _33458_, _06352_);
  or _84106_ (_33493_, _33492_, _06345_);
  or _84107_ (_33494_, _33493_, _33491_);
  or _84108_ (_33495_, _33466_, _06346_);
  and _84109_ (_33496_, _33495_, _06340_);
  and _84110_ (_33498_, _33496_, _33494_);
  or _84111_ (_33499_, _33477_, _16663_);
  and _84112_ (_33500_, _33499_, _06339_);
  and _84113_ (_33501_, _33500_, _33479_);
  or _84114_ (_33502_, _33501_, _10153_);
  or _84115_ (_33503_, _33502_, _33498_);
  or _84116_ (_33504_, _33484_, _06327_);
  and _84117_ (_33505_, _33504_, _33503_);
  or _84118_ (_33506_, _33505_, _09572_);
  and _84119_ (_33507_, _09447_, _08022_);
  or _84120_ (_33509_, _33458_, _06333_);
  or _84121_ (_33510_, _33509_, _33507_);
  and _84122_ (_33511_, _33510_, _06313_);
  and _84123_ (_33512_, _33511_, _33506_);
  and _84124_ (_33513_, _14666_, _08022_);
  or _84125_ (_33514_, _33513_, _33458_);
  and _84126_ (_33515_, _33514_, _06037_);
  or _84127_ (_33516_, _33515_, _06277_);
  or _84128_ (_33517_, _33516_, _33512_);
  and _84129_ (_33518_, _08022_, _09008_);
  or _84130_ (_33520_, _33518_, _33458_);
  or _84131_ (_33521_, _33520_, _06278_);
  and _84132_ (_33522_, _33521_, _33517_);
  or _84133_ (_33523_, _33522_, _06502_);
  and _84134_ (_33524_, _14566_, _08022_);
  or _84135_ (_33525_, _33458_, _07334_);
  or _84136_ (_33526_, _33525_, _33524_);
  and _84137_ (_33527_, _33526_, _07337_);
  and _84138_ (_33528_, _33527_, _33523_);
  or _84139_ (_33529_, _33528_, _33463_);
  and _84140_ (_33531_, _33529_, _07339_);
  nand _84141_ (_33532_, _33520_, _06507_);
  nor _84142_ (_33533_, _33532_, _33465_);
  or _84143_ (_33534_, _33533_, _06610_);
  or _84144_ (_33535_, _33534_, _33531_);
  or _84145_ (_33536_, _33461_, _33458_);
  or _84146_ (_33537_, _33536_, _07331_);
  and _84147_ (_33538_, _33537_, _33535_);
  or _84148_ (_33539_, _33538_, _06509_);
  and _84149_ (_33540_, _14563_, _08022_);
  or _84150_ (_33542_, _33458_, _09107_);
  or _84151_ (_33543_, _33542_, _33540_);
  and _84152_ (_33544_, _33543_, _09112_);
  and _84153_ (_33545_, _33544_, _33539_);
  and _84154_ (_33546_, _33460_, _06602_);
  or _84155_ (_33547_, _33546_, _06639_);
  or _84156_ (_33548_, _33547_, _33545_);
  or _84157_ (_33549_, _33466_, _07048_);
  and _84158_ (_33550_, _33549_, _33548_);
  or _84159_ (_33551_, _33550_, _05989_);
  or _84160_ (_33553_, _33458_, _05990_);
  and _84161_ (_33554_, _33553_, _33551_);
  or _84162_ (_33555_, _33554_, _06646_);
  or _84163_ (_33556_, _33466_, _06651_);
  and _84164_ (_33557_, _33556_, _01442_);
  and _84165_ (_33558_, _33557_, _33555_);
  or _84166_ (_33559_, _33558_, _33457_);
  and _84167_ (_44257_, _33559_, _43634_);
  and _84168_ (_33560_, _01446_, \oc8051_golden_model_1.IP [1]);
  and _84169_ (_33561_, _13693_, \oc8051_golden_model_1.IP [1]);
  nor _84170_ (_33563_, _10578_, _13693_);
  or _84171_ (_33564_, _33563_, _33561_);
  or _84172_ (_33565_, _33564_, _09112_);
  nand _84173_ (_33566_, _08022_, _07160_);
  or _84174_ (_33567_, _08022_, \oc8051_golden_model_1.IP [1]);
  and _84175_ (_33568_, _33567_, _06277_);
  and _84176_ (_33569_, _33568_, _33566_);
  nor _84177_ (_33570_, _13693_, _07448_);
  or _84178_ (_33571_, _33570_, _33561_);
  or _84179_ (_33572_, _33571_, _06772_);
  and _84180_ (_33574_, _14744_, _08022_);
  not _84181_ (_33575_, _33574_);
  and _84182_ (_33576_, _33575_, _33567_);
  or _84183_ (_33577_, _33576_, _07275_);
  and _84184_ (_33578_, _08022_, \oc8051_golden_model_1.ACC [1]);
  or _84185_ (_33579_, _33578_, _33561_);
  and _84186_ (_33580_, _33579_, _07259_);
  and _84187_ (_33581_, _07260_, \oc8051_golden_model_1.IP [1]);
  or _84188_ (_33582_, _33581_, _06474_);
  or _84189_ (_33583_, _33582_, _33580_);
  and _84190_ (_33585_, _33583_, _06357_);
  and _84191_ (_33586_, _33585_, _33577_);
  and _84192_ (_33587_, _13701_, \oc8051_golden_model_1.IP [1]);
  and _84193_ (_33588_, _14767_, _08643_);
  or _84194_ (_33589_, _33588_, _33587_);
  and _84195_ (_33590_, _33589_, _06356_);
  or _84196_ (_33591_, _33590_, _06410_);
  or _84197_ (_33592_, _33591_, _33586_);
  and _84198_ (_33593_, _33592_, _33572_);
  or _84199_ (_33594_, _33593_, _06417_);
  or _84200_ (_33596_, _33579_, _06426_);
  and _84201_ (_33597_, _33596_, _06353_);
  and _84202_ (_33598_, _33597_, _33594_);
  and _84203_ (_33599_, _14754_, _08643_);
  or _84204_ (_33600_, _33599_, _33587_);
  and _84205_ (_33601_, _33600_, _06352_);
  or _84206_ (_33602_, _33601_, _06345_);
  or _84207_ (_33603_, _33602_, _33598_);
  and _84208_ (_33604_, _33588_, _14782_);
  or _84209_ (_33605_, _33587_, _06346_);
  or _84210_ (_33607_, _33605_, _33604_);
  and _84211_ (_33608_, _33607_, _33603_);
  and _84212_ (_33609_, _33608_, _06340_);
  and _84213_ (_33610_, _14796_, _08643_);
  or _84214_ (_33611_, _33587_, _33610_);
  and _84215_ (_33612_, _33611_, _06339_);
  or _84216_ (_33613_, _33612_, _10153_);
  or _84217_ (_33614_, _33613_, _33609_);
  or _84218_ (_33615_, _33571_, _06327_);
  and _84219_ (_33616_, _33615_, _33614_);
  or _84220_ (_33618_, _33616_, _09572_);
  and _84221_ (_33619_, _09402_, _08022_);
  or _84222_ (_33620_, _33561_, _06333_);
  or _84223_ (_33621_, _33620_, _33619_);
  and _84224_ (_33622_, _33621_, _06313_);
  and _84225_ (_33623_, _33622_, _33618_);
  and _84226_ (_33624_, _14851_, _08022_);
  or _84227_ (_33625_, _33624_, _33561_);
  and _84228_ (_33626_, _33625_, _06037_);
  or _84229_ (_33627_, _33626_, _33623_);
  and _84230_ (_33629_, _33627_, _06278_);
  or _84231_ (_33630_, _33629_, _33569_);
  and _84232_ (_33631_, _33630_, _07334_);
  or _84233_ (_33632_, _14749_, _13693_);
  and _84234_ (_33633_, _33567_, _06502_);
  and _84235_ (_33634_, _33633_, _33632_);
  or _84236_ (_33635_, _33634_, _06615_);
  or _84237_ (_33636_, _33635_, _33631_);
  and _84238_ (_33637_, _10579_, _08022_);
  or _84239_ (_33638_, _33637_, _33561_);
  or _84240_ (_33640_, _33638_, _07337_);
  and _84241_ (_33641_, _33640_, _07339_);
  and _84242_ (_33642_, _33641_, _33636_);
  or _84243_ (_33643_, _14747_, _13693_);
  and _84244_ (_33644_, _33567_, _06507_);
  and _84245_ (_33645_, _33644_, _33643_);
  or _84246_ (_33646_, _33645_, _06610_);
  or _84247_ (_33647_, _33646_, _33642_);
  and _84248_ (_33648_, _33578_, _08404_);
  or _84249_ (_33649_, _33561_, _07331_);
  or _84250_ (_33651_, _33649_, _33648_);
  and _84251_ (_33652_, _33651_, _09107_);
  and _84252_ (_33653_, _33652_, _33647_);
  or _84253_ (_33654_, _33566_, _08404_);
  and _84254_ (_33655_, _33567_, _06509_);
  and _84255_ (_33656_, _33655_, _33654_);
  or _84256_ (_33657_, _33656_, _06602_);
  or _84257_ (_33658_, _33657_, _33653_);
  and _84258_ (_33659_, _33658_, _33565_);
  or _84259_ (_33660_, _33659_, _06639_);
  or _84260_ (_33662_, _33576_, _07048_);
  and _84261_ (_33663_, _33662_, _05990_);
  and _84262_ (_33664_, _33663_, _33660_);
  and _84263_ (_33665_, _33600_, _05989_);
  or _84264_ (_33666_, _33665_, _06646_);
  or _84265_ (_33667_, _33666_, _33664_);
  or _84266_ (_33668_, _33561_, _06651_);
  or _84267_ (_33669_, _33668_, _33574_);
  and _84268_ (_33670_, _33669_, _01442_);
  and _84269_ (_33671_, _33670_, _33667_);
  or _84270_ (_33673_, _33671_, _33560_);
  and _84271_ (_44258_, _33673_, _43634_);
  and _84272_ (_33674_, _01446_, \oc8051_golden_model_1.IP [2]);
  and _84273_ (_33675_, _13693_, \oc8051_golden_model_1.IP [2]);
  nor _84274_ (_33676_, _13693_, _07854_);
  or _84275_ (_33677_, _33676_, _33675_);
  or _84276_ (_33678_, _33677_, _06327_);
  or _84277_ (_33679_, _33677_, _06772_);
  and _84278_ (_33680_, _14959_, _08022_);
  or _84279_ (_33681_, _33680_, _33675_);
  or _84280_ (_33683_, _33681_, _07275_);
  and _84281_ (_33684_, _08022_, \oc8051_golden_model_1.ACC [2]);
  or _84282_ (_33685_, _33684_, _33675_);
  and _84283_ (_33686_, _33685_, _07259_);
  and _84284_ (_33687_, _07260_, \oc8051_golden_model_1.IP [2]);
  or _84285_ (_33688_, _33687_, _06474_);
  or _84286_ (_33689_, _33688_, _33686_);
  and _84287_ (_33690_, _33689_, _06357_);
  and _84288_ (_33691_, _33690_, _33683_);
  and _84289_ (_33692_, _13701_, \oc8051_golden_model_1.IP [2]);
  and _84290_ (_33694_, _14955_, _08643_);
  or _84291_ (_33695_, _33694_, _33692_);
  and _84292_ (_33696_, _33695_, _06356_);
  or _84293_ (_33697_, _33696_, _06410_);
  or _84294_ (_33698_, _33697_, _33691_);
  and _84295_ (_33699_, _33698_, _33679_);
  or _84296_ (_33700_, _33699_, _06417_);
  or _84297_ (_33701_, _33685_, _06426_);
  and _84298_ (_33702_, _33701_, _06353_);
  and _84299_ (_33703_, _33702_, _33700_);
  and _84300_ (_33705_, _14953_, _08643_);
  or _84301_ (_33706_, _33705_, _33692_);
  and _84302_ (_33707_, _33706_, _06352_);
  or _84303_ (_33708_, _33707_, _06345_);
  or _84304_ (_33709_, _33708_, _33703_);
  and _84305_ (_33710_, _33694_, _14986_);
  or _84306_ (_33711_, _33692_, _06346_);
  or _84307_ (_33712_, _33711_, _33710_);
  and _84308_ (_33713_, _33712_, _06340_);
  and _84309_ (_33714_, _33713_, _33709_);
  and _84310_ (_33716_, _15000_, _08643_);
  or _84311_ (_33717_, _33716_, _33692_);
  and _84312_ (_33718_, _33717_, _06339_);
  or _84313_ (_33719_, _33718_, _10153_);
  or _84314_ (_33720_, _33719_, _33714_);
  and _84315_ (_33721_, _33720_, _33678_);
  or _84316_ (_33722_, _33721_, _09572_);
  and _84317_ (_33723_, _09356_, _08022_);
  or _84318_ (_33724_, _33675_, _06333_);
  or _84319_ (_33725_, _33724_, _33723_);
  and _84320_ (_33727_, _33725_, _06313_);
  and _84321_ (_33728_, _33727_, _33722_);
  and _84322_ (_33729_, _15056_, _08022_);
  or _84323_ (_33730_, _33729_, _33675_);
  and _84324_ (_33731_, _33730_, _06037_);
  or _84325_ (_33732_, _33731_, _06277_);
  or _84326_ (_33733_, _33732_, _33728_);
  and _84327_ (_33734_, _08022_, _09057_);
  or _84328_ (_33735_, _33734_, _33675_);
  or _84329_ (_33736_, _33735_, _06278_);
  and _84330_ (_33738_, _33736_, _33733_);
  or _84331_ (_33739_, _33738_, _06502_);
  and _84332_ (_33740_, _14948_, _08022_);
  or _84333_ (_33741_, _33675_, _07334_);
  or _84334_ (_33742_, _33741_, _33740_);
  and _84335_ (_33743_, _33742_, _07337_);
  and _84336_ (_33744_, _33743_, _33739_);
  and _84337_ (_33745_, _10583_, _08022_);
  or _84338_ (_33746_, _33745_, _33675_);
  and _84339_ (_33747_, _33746_, _06615_);
  or _84340_ (_33749_, _33747_, _33744_);
  and _84341_ (_33750_, _33749_, _07339_);
  or _84342_ (_33751_, _33675_, _08503_);
  and _84343_ (_33752_, _33735_, _06507_);
  and _84344_ (_33753_, _33752_, _33751_);
  or _84345_ (_33754_, _33753_, _33750_);
  and _84346_ (_33755_, _33754_, _07331_);
  and _84347_ (_33756_, _33685_, _06610_);
  and _84348_ (_33757_, _33756_, _33751_);
  or _84349_ (_33758_, _33757_, _06509_);
  or _84350_ (_33760_, _33758_, _33755_);
  and _84351_ (_33761_, _14945_, _08022_);
  or _84352_ (_33762_, _33675_, _09107_);
  or _84353_ (_33763_, _33762_, _33761_);
  and _84354_ (_33764_, _33763_, _09112_);
  and _84355_ (_33765_, _33764_, _33760_);
  nor _84356_ (_33766_, _10582_, _13693_);
  or _84357_ (_33767_, _33766_, _33675_);
  and _84358_ (_33768_, _33767_, _06602_);
  or _84359_ (_33769_, _33768_, _06639_);
  or _84360_ (_33771_, _33769_, _33765_);
  or _84361_ (_33772_, _33681_, _07048_);
  and _84362_ (_33773_, _33772_, _05990_);
  and _84363_ (_33774_, _33773_, _33771_);
  and _84364_ (_33775_, _33706_, _05989_);
  or _84365_ (_33776_, _33775_, _06646_);
  or _84366_ (_33777_, _33776_, _33774_);
  and _84367_ (_33778_, _15129_, _08022_);
  or _84368_ (_33779_, _33675_, _06651_);
  or _84369_ (_33780_, _33779_, _33778_);
  and _84370_ (_33782_, _33780_, _01442_);
  and _84371_ (_33783_, _33782_, _33777_);
  or _84372_ (_33784_, _33783_, _33674_);
  and _84373_ (_44259_, _33784_, _43634_);
  and _84374_ (_33785_, _01446_, \oc8051_golden_model_1.IP [3]);
  and _84375_ (_33786_, _13693_, \oc8051_golden_model_1.IP [3]);
  nor _84376_ (_33787_, _13693_, _07680_);
  or _84377_ (_33788_, _33787_, _33786_);
  or _84378_ (_33789_, _33788_, _06327_);
  and _84379_ (_33790_, _15153_, _08022_);
  or _84380_ (_33792_, _33790_, _33786_);
  or _84381_ (_33793_, _33792_, _07275_);
  and _84382_ (_33794_, _08022_, \oc8051_golden_model_1.ACC [3]);
  or _84383_ (_33795_, _33794_, _33786_);
  and _84384_ (_33796_, _33795_, _07259_);
  and _84385_ (_33797_, _07260_, \oc8051_golden_model_1.IP [3]);
  or _84386_ (_33798_, _33797_, _06474_);
  or _84387_ (_33799_, _33798_, _33796_);
  and _84388_ (_33800_, _33799_, _06357_);
  and _84389_ (_33801_, _33800_, _33793_);
  and _84390_ (_33803_, _13701_, \oc8051_golden_model_1.IP [3]);
  and _84391_ (_33804_, _15150_, _08643_);
  or _84392_ (_33805_, _33804_, _33803_);
  and _84393_ (_33806_, _33805_, _06356_);
  or _84394_ (_33807_, _33806_, _06410_);
  or _84395_ (_33808_, _33807_, _33801_);
  or _84396_ (_33809_, _33788_, _06772_);
  and _84397_ (_33810_, _33809_, _33808_);
  or _84398_ (_33811_, _33810_, _06417_);
  or _84399_ (_33812_, _33795_, _06426_);
  and _84400_ (_33814_, _33812_, _06353_);
  and _84401_ (_33815_, _33814_, _33811_);
  and _84402_ (_33816_, _15148_, _08643_);
  or _84403_ (_33817_, _33816_, _33803_);
  and _84404_ (_33818_, _33817_, _06352_);
  or _84405_ (_33819_, _33818_, _06345_);
  or _84406_ (_33820_, _33819_, _33815_);
  or _84407_ (_33821_, _33803_, _15180_);
  and _84408_ (_33822_, _33821_, _33805_);
  or _84409_ (_33823_, _33822_, _06346_);
  and _84410_ (_33825_, _33823_, _06340_);
  and _84411_ (_33826_, _33825_, _33820_);
  and _84412_ (_33827_, _15197_, _08643_);
  or _84413_ (_33828_, _33827_, _33803_);
  and _84414_ (_33829_, _33828_, _06339_);
  or _84415_ (_33830_, _33829_, _10153_);
  or _84416_ (_33831_, _33830_, _33826_);
  and _84417_ (_33832_, _33831_, _33789_);
  or _84418_ (_33833_, _33832_, _09572_);
  and _84419_ (_33834_, _09310_, _08022_);
  or _84420_ (_33836_, _33786_, _06333_);
  or _84421_ (_33837_, _33836_, _33834_);
  and _84422_ (_33838_, _33837_, _06313_);
  and _84423_ (_33839_, _33838_, _33833_);
  and _84424_ (_33840_, _15251_, _08022_);
  or _84425_ (_33841_, _33840_, _33786_);
  and _84426_ (_33842_, _33841_, _06037_);
  or _84427_ (_33843_, _33842_, _06277_);
  or _84428_ (_33844_, _33843_, _33839_);
  and _84429_ (_33845_, _08022_, _09014_);
  or _84430_ (_33846_, _33845_, _33786_);
  or _84431_ (_33847_, _33846_, _06278_);
  and _84432_ (_33848_, _33847_, _33844_);
  or _84433_ (_33849_, _33848_, _06502_);
  and _84434_ (_33850_, _15266_, _08022_);
  or _84435_ (_33851_, _33786_, _07334_);
  or _84436_ (_33852_, _33851_, _33850_);
  and _84437_ (_33853_, _33852_, _07337_);
  and _84438_ (_33854_, _33853_, _33849_);
  and _84439_ (_33855_, _12619_, _08022_);
  or _84440_ (_33857_, _33855_, _33786_);
  and _84441_ (_33858_, _33857_, _06615_);
  or _84442_ (_33859_, _33858_, _33854_);
  and _84443_ (_33860_, _33859_, _07339_);
  or _84444_ (_33861_, _33786_, _08359_);
  and _84445_ (_33862_, _33846_, _06507_);
  and _84446_ (_33863_, _33862_, _33861_);
  or _84447_ (_33864_, _33863_, _33860_);
  and _84448_ (_33865_, _33864_, _07331_);
  and _84449_ (_33866_, _33795_, _06610_);
  and _84450_ (_33868_, _33866_, _33861_);
  or _84451_ (_33869_, _33868_, _06509_);
  or _84452_ (_33870_, _33869_, _33865_);
  and _84453_ (_33871_, _15263_, _08022_);
  or _84454_ (_33872_, _33786_, _09107_);
  or _84455_ (_33873_, _33872_, _33871_);
  and _84456_ (_33874_, _33873_, _09112_);
  and _84457_ (_33875_, _33874_, _33870_);
  nor _84458_ (_33876_, _10574_, _13693_);
  or _84459_ (_33877_, _33876_, _33786_);
  and _84460_ (_33879_, _33877_, _06602_);
  or _84461_ (_33880_, _33879_, _06639_);
  or _84462_ (_33881_, _33880_, _33875_);
  or _84463_ (_33882_, _33792_, _07048_);
  and _84464_ (_33883_, _33882_, _05990_);
  and _84465_ (_33884_, _33883_, _33881_);
  and _84466_ (_33885_, _33817_, _05989_);
  or _84467_ (_33886_, _33885_, _06646_);
  or _84468_ (_33887_, _33886_, _33884_);
  and _84469_ (_33888_, _15321_, _08022_);
  or _84470_ (_33890_, _33786_, _06651_);
  or _84471_ (_33891_, _33890_, _33888_);
  and _84472_ (_33892_, _33891_, _01442_);
  and _84473_ (_33893_, _33892_, _33887_);
  or _84474_ (_33894_, _33893_, _33785_);
  and _84475_ (_44260_, _33894_, _43634_);
  and _84476_ (_33895_, _01446_, \oc8051_golden_model_1.IP [4]);
  and _84477_ (_33896_, _13693_, \oc8051_golden_model_1.IP [4]);
  nor _84478_ (_33897_, _10589_, _13693_);
  or _84479_ (_33898_, _33897_, _33896_);
  and _84480_ (_33900_, _08022_, \oc8051_golden_model_1.ACC [4]);
  nand _84481_ (_33901_, _33900_, _08599_);
  and _84482_ (_33902_, _33901_, _06615_);
  and _84483_ (_33903_, _33902_, _33898_);
  nor _84484_ (_33904_, _08596_, _13693_);
  or _84485_ (_33905_, _33904_, _33896_);
  or _84486_ (_33906_, _33905_, _06327_);
  and _84487_ (_33907_, _13701_, \oc8051_golden_model_1.IP [4]);
  and _84488_ (_33908_, _15348_, _08643_);
  or _84489_ (_33909_, _33908_, _33907_);
  and _84490_ (_33911_, _33909_, _06352_);
  and _84491_ (_33912_, _15367_, _08022_);
  or _84492_ (_33913_, _33912_, _33896_);
  or _84493_ (_33914_, _33913_, _07275_);
  or _84494_ (_33915_, _33900_, _33896_);
  and _84495_ (_33916_, _33915_, _07259_);
  and _84496_ (_33917_, _07260_, \oc8051_golden_model_1.IP [4]);
  or _84497_ (_33918_, _33917_, _06474_);
  or _84498_ (_33919_, _33918_, _33916_);
  and _84499_ (_33920_, _33919_, _06357_);
  and _84500_ (_33922_, _33920_, _33914_);
  and _84501_ (_33923_, _15353_, _08643_);
  or _84502_ (_33924_, _33923_, _33907_);
  and _84503_ (_33925_, _33924_, _06356_);
  or _84504_ (_33926_, _33925_, _06410_);
  or _84505_ (_33927_, _33926_, _33922_);
  or _84506_ (_33928_, _33905_, _06772_);
  and _84507_ (_33929_, _33928_, _33927_);
  or _84508_ (_33930_, _33929_, _06417_);
  or _84509_ (_33931_, _33915_, _06426_);
  and _84510_ (_33933_, _33931_, _06353_);
  and _84511_ (_33934_, _33933_, _33930_);
  or _84512_ (_33935_, _33934_, _33911_);
  and _84513_ (_33936_, _33935_, _06346_);
  and _84514_ (_33937_, _15385_, _08643_);
  or _84515_ (_33938_, _33937_, _33907_);
  and _84516_ (_33939_, _33938_, _06345_);
  or _84517_ (_33940_, _33939_, _33936_);
  and _84518_ (_33941_, _33940_, _06340_);
  and _84519_ (_33942_, _15350_, _08643_);
  or _84520_ (_33944_, _33942_, _33907_);
  and _84521_ (_33945_, _33944_, _06339_);
  or _84522_ (_33946_, _33945_, _10153_);
  or _84523_ (_33947_, _33946_, _33941_);
  and _84524_ (_33948_, _33947_, _33906_);
  or _84525_ (_33949_, _33948_, _09572_);
  and _84526_ (_33950_, _09264_, _08022_);
  or _84527_ (_33951_, _33896_, _06333_);
  or _84528_ (_33952_, _33951_, _33950_);
  and _84529_ (_33953_, _33952_, _06313_);
  and _84530_ (_33955_, _33953_, _33949_);
  and _84531_ (_33956_, _15452_, _08022_);
  or _84532_ (_33957_, _33956_, _33896_);
  and _84533_ (_33958_, _33957_, _06037_);
  or _84534_ (_33959_, _33958_, _06277_);
  or _84535_ (_33960_, _33959_, _33955_);
  and _84536_ (_33961_, _08995_, _08022_);
  or _84537_ (_33962_, _33961_, _33896_);
  or _84538_ (_33963_, _33962_, _06278_);
  and _84539_ (_33964_, _33963_, _33960_);
  or _84540_ (_33966_, _33964_, _06502_);
  and _84541_ (_33967_, _15345_, _08022_);
  or _84542_ (_33968_, _33896_, _07334_);
  or _84543_ (_33969_, _33968_, _33967_);
  and _84544_ (_33970_, _33969_, _07337_);
  and _84545_ (_33971_, _33970_, _33966_);
  or _84546_ (_33972_, _33971_, _33903_);
  and _84547_ (_33973_, _33972_, _07339_);
  or _84548_ (_33974_, _33896_, _08599_);
  and _84549_ (_33975_, _33962_, _06507_);
  and _84550_ (_33977_, _33975_, _33974_);
  or _84551_ (_33978_, _33977_, _33973_);
  and _84552_ (_33979_, _33978_, _07331_);
  and _84553_ (_33980_, _33915_, _06610_);
  and _84554_ (_33981_, _33980_, _33974_);
  or _84555_ (_33982_, _33981_, _06509_);
  or _84556_ (_33983_, _33982_, _33979_);
  and _84557_ (_33984_, _15342_, _08022_);
  or _84558_ (_33985_, _33896_, _09107_);
  or _84559_ (_33986_, _33985_, _33984_);
  and _84560_ (_33988_, _33986_, _09112_);
  and _84561_ (_33989_, _33988_, _33983_);
  and _84562_ (_33990_, _33898_, _06602_);
  or _84563_ (_33991_, _33990_, _06639_);
  or _84564_ (_33992_, _33991_, _33989_);
  or _84565_ (_33993_, _33913_, _07048_);
  and _84566_ (_33994_, _33993_, _05990_);
  and _84567_ (_33995_, _33994_, _33992_);
  and _84568_ (_33996_, _33909_, _05989_);
  or _84569_ (_33997_, _33996_, _06646_);
  or _84570_ (_33999_, _33997_, _33995_);
  and _84571_ (_34000_, _15524_, _08022_);
  or _84572_ (_34001_, _33896_, _06651_);
  or _84573_ (_34002_, _34001_, _34000_);
  and _84574_ (_34003_, _34002_, _01442_);
  and _84575_ (_34004_, _34003_, _33999_);
  or _84576_ (_34005_, _34004_, _33895_);
  and _84577_ (_44261_, _34005_, _43634_);
  and _84578_ (_34006_, _01446_, \oc8051_golden_model_1.IP [5]);
  and _84579_ (_34007_, _13693_, \oc8051_golden_model_1.IP [5]);
  and _84580_ (_34009_, _15550_, _08022_);
  or _84581_ (_34010_, _34009_, _34007_);
  or _84582_ (_34011_, _34010_, _07275_);
  and _84583_ (_34012_, _08022_, \oc8051_golden_model_1.ACC [5]);
  or _84584_ (_34013_, _34012_, _34007_);
  and _84585_ (_34014_, _34013_, _07259_);
  and _84586_ (_34015_, _07260_, \oc8051_golden_model_1.IP [5]);
  or _84587_ (_34016_, _34015_, _06474_);
  or _84588_ (_34017_, _34016_, _34014_);
  and _84589_ (_34018_, _34017_, _06357_);
  and _84590_ (_34020_, _34018_, _34011_);
  and _84591_ (_34021_, _13701_, \oc8051_golden_model_1.IP [5]);
  and _84592_ (_34022_, _15566_, _08643_);
  or _84593_ (_34023_, _34022_, _34021_);
  and _84594_ (_34024_, _34023_, _06356_);
  or _84595_ (_34025_, _34024_, _06410_);
  or _84596_ (_34026_, _34025_, _34020_);
  nor _84597_ (_34027_, _08305_, _13693_);
  or _84598_ (_34028_, _34027_, _34007_);
  or _84599_ (_34029_, _34028_, _06772_);
  and _84600_ (_34031_, _34029_, _34026_);
  or _84601_ (_34032_, _34031_, _06417_);
  or _84602_ (_34033_, _34013_, _06426_);
  and _84603_ (_34034_, _34033_, _06353_);
  and _84604_ (_34035_, _34034_, _34032_);
  and _84605_ (_34036_, _15544_, _08643_);
  or _84606_ (_34037_, _34036_, _34021_);
  and _84607_ (_34038_, _34037_, _06352_);
  or _84608_ (_34039_, _34038_, _06345_);
  or _84609_ (_34040_, _34039_, _34035_);
  or _84610_ (_34042_, _34021_, _15581_);
  and _84611_ (_34043_, _34042_, _34023_);
  or _84612_ (_34044_, _34043_, _06346_);
  and _84613_ (_34045_, _34044_, _06340_);
  and _84614_ (_34046_, _34045_, _34040_);
  and _84615_ (_34047_, _15546_, _08643_);
  or _84616_ (_34048_, _34047_, _34021_);
  and _84617_ (_34049_, _34048_, _06339_);
  or _84618_ (_34050_, _34049_, _10153_);
  or _84619_ (_34051_, _34050_, _34046_);
  or _84620_ (_34053_, _34028_, _06327_);
  and _84621_ (_34054_, _34053_, _34051_);
  or _84622_ (_34055_, _34054_, _09572_);
  and _84623_ (_34056_, _09218_, _08022_);
  or _84624_ (_34057_, _34007_, _06333_);
  or _84625_ (_34058_, _34057_, _34056_);
  and _84626_ (_34059_, _34058_, _06313_);
  and _84627_ (_34060_, _34059_, _34055_);
  and _84628_ (_34061_, _15649_, _08022_);
  or _84629_ (_34062_, _34061_, _34007_);
  and _84630_ (_34064_, _34062_, _06037_);
  or _84631_ (_34065_, _34064_, _06277_);
  or _84632_ (_34066_, _34065_, _34060_);
  and _84633_ (_34067_, _08954_, _08022_);
  or _84634_ (_34068_, _34067_, _34007_);
  or _84635_ (_34069_, _34068_, _06278_);
  and _84636_ (_34070_, _34069_, _34066_);
  or _84637_ (_34071_, _34070_, _06502_);
  and _84638_ (_34072_, _15664_, _08022_);
  or _84639_ (_34073_, _34007_, _07334_);
  or _84640_ (_34075_, _34073_, _34072_);
  and _84641_ (_34076_, _34075_, _07337_);
  and _84642_ (_34077_, _34076_, _34071_);
  and _84643_ (_34078_, _12626_, _08022_);
  or _84644_ (_34079_, _34078_, _34007_);
  and _84645_ (_34080_, _34079_, _06615_);
  or _84646_ (_34081_, _34080_, _34077_);
  and _84647_ (_34082_, _34081_, _07339_);
  or _84648_ (_34083_, _34007_, _08308_);
  and _84649_ (_34084_, _34068_, _06507_);
  and _84650_ (_34086_, _34084_, _34083_);
  or _84651_ (_34087_, _34086_, _34082_);
  and _84652_ (_34088_, _34087_, _07331_);
  and _84653_ (_34089_, _34013_, _06610_);
  and _84654_ (_34090_, _34089_, _34083_);
  or _84655_ (_34091_, _34090_, _06509_);
  or _84656_ (_34092_, _34091_, _34088_);
  and _84657_ (_34093_, _15663_, _08022_);
  or _84658_ (_34094_, _34007_, _09107_);
  or _84659_ (_34095_, _34094_, _34093_);
  and _84660_ (_34097_, _34095_, _09112_);
  and _84661_ (_34098_, _34097_, _34092_);
  nor _84662_ (_34099_, _10570_, _13693_);
  or _84663_ (_34100_, _34099_, _34007_);
  and _84664_ (_34101_, _34100_, _06602_);
  or _84665_ (_34102_, _34101_, _06639_);
  or _84666_ (_34103_, _34102_, _34098_);
  or _84667_ (_34104_, _34010_, _07048_);
  and _84668_ (_34105_, _34104_, _05990_);
  and _84669_ (_34106_, _34105_, _34103_);
  and _84670_ (_34108_, _34037_, _05989_);
  or _84671_ (_34109_, _34108_, _06646_);
  or _84672_ (_34110_, _34109_, _34106_);
  and _84673_ (_34111_, _15721_, _08022_);
  or _84674_ (_34112_, _34007_, _06651_);
  or _84675_ (_34113_, _34112_, _34111_);
  and _84676_ (_34114_, _34113_, _01442_);
  and _84677_ (_34115_, _34114_, _34110_);
  or _84678_ (_34116_, _34115_, _34006_);
  and _84679_ (_44263_, _34116_, _43634_);
  and _84680_ (_34118_, _01446_, \oc8051_golden_model_1.IP [6]);
  and _84681_ (_34119_, _13693_, \oc8051_golden_model_1.IP [6]);
  nor _84682_ (_34120_, _10595_, _13693_);
  or _84683_ (_34121_, _34120_, _34119_);
  and _84684_ (_34122_, _08022_, \oc8051_golden_model_1.ACC [6]);
  nand _84685_ (_34123_, _34122_, _08212_);
  and _84686_ (_34124_, _34123_, _06615_);
  and _84687_ (_34125_, _34124_, _34121_);
  and _84688_ (_34126_, _15759_, _08022_);
  or _84689_ (_34127_, _34126_, _34119_);
  or _84690_ (_34129_, _34127_, _07275_);
  or _84691_ (_34130_, _34122_, _34119_);
  and _84692_ (_34131_, _34130_, _07259_);
  and _84693_ (_34132_, _07260_, \oc8051_golden_model_1.IP [6]);
  or _84694_ (_34133_, _34132_, _06474_);
  or _84695_ (_34134_, _34133_, _34131_);
  and _84696_ (_34135_, _34134_, _06357_);
  and _84697_ (_34136_, _34135_, _34129_);
  and _84698_ (_34138_, _13701_, \oc8051_golden_model_1.IP [6]);
  and _84699_ (_34140_, _15763_, _08643_);
  or _84700_ (_34143_, _34140_, _34138_);
  and _84701_ (_34145_, _34143_, _06356_);
  or _84702_ (_34147_, _34145_, _06410_);
  or _84703_ (_34149_, _34147_, _34136_);
  nor _84704_ (_34151_, _08209_, _13693_);
  or _84705_ (_34153_, _34151_, _34119_);
  or _84706_ (_34155_, _34153_, _06772_);
  and _84707_ (_34157_, _34155_, _34149_);
  or _84708_ (_34158_, _34157_, _06417_);
  or _84709_ (_34159_, _34130_, _06426_);
  and _84710_ (_34161_, _34159_, _06353_);
  and _84711_ (_34162_, _34161_, _34158_);
  and _84712_ (_34163_, _15743_, _08643_);
  or _84713_ (_34164_, _34163_, _34138_);
  and _84714_ (_34165_, _34164_, _06352_);
  or _84715_ (_34166_, _34165_, _06345_);
  or _84716_ (_34167_, _34166_, _34162_);
  or _84717_ (_34168_, _34138_, _15778_);
  and _84718_ (_34169_, _34168_, _34143_);
  or _84719_ (_34170_, _34169_, _06346_);
  and _84720_ (_34172_, _34170_, _06340_);
  and _84721_ (_34173_, _34172_, _34167_);
  and _84722_ (_34174_, _15745_, _08643_);
  or _84723_ (_34175_, _34174_, _34138_);
  and _84724_ (_34176_, _34175_, _06339_);
  or _84725_ (_34177_, _34176_, _10153_);
  or _84726_ (_34178_, _34177_, _34173_);
  or _84727_ (_34179_, _34153_, _06327_);
  and _84728_ (_34180_, _34179_, _34178_);
  or _84729_ (_34181_, _34180_, _09572_);
  and _84730_ (_34183_, _09172_, _08022_);
  or _84731_ (_34184_, _34119_, _06333_);
  or _84732_ (_34185_, _34184_, _34183_);
  and _84733_ (_34186_, _34185_, _06313_);
  and _84734_ (_34187_, _34186_, _34181_);
  and _84735_ (_34188_, _15846_, _08022_);
  or _84736_ (_34189_, _34188_, _34119_);
  and _84737_ (_34190_, _34189_, _06037_);
  or _84738_ (_34191_, _34190_, _06277_);
  or _84739_ (_34192_, _34191_, _34187_);
  and _84740_ (_34194_, _15853_, _08022_);
  or _84741_ (_34195_, _34194_, _34119_);
  or _84742_ (_34196_, _34195_, _06278_);
  and _84743_ (_34197_, _34196_, _34192_);
  or _84744_ (_34198_, _34197_, _06502_);
  and _84745_ (_34199_, _15862_, _08022_);
  or _84746_ (_34200_, _34119_, _07334_);
  or _84747_ (_34201_, _34200_, _34199_);
  and _84748_ (_34202_, _34201_, _07337_);
  and _84749_ (_34203_, _34202_, _34198_);
  or _84750_ (_34205_, _34203_, _34125_);
  and _84751_ (_34206_, _34205_, _07339_);
  or _84752_ (_34207_, _34119_, _08212_);
  and _84753_ (_34208_, _34195_, _06507_);
  and _84754_ (_34209_, _34208_, _34207_);
  or _84755_ (_34210_, _34209_, _34206_);
  and _84756_ (_34211_, _34210_, _07331_);
  and _84757_ (_34212_, _34130_, _06610_);
  and _84758_ (_34213_, _34212_, _34207_);
  or _84759_ (_34214_, _34213_, _06509_);
  or _84760_ (_34216_, _34214_, _34211_);
  and _84761_ (_34217_, _15859_, _08022_);
  or _84762_ (_34218_, _34119_, _09107_);
  or _84763_ (_34219_, _34218_, _34217_);
  and _84764_ (_34220_, _34219_, _09112_);
  and _84765_ (_34221_, _34220_, _34216_);
  and _84766_ (_34222_, _34121_, _06602_);
  or _84767_ (_34223_, _34222_, _06639_);
  or _84768_ (_34224_, _34223_, _34221_);
  or _84769_ (_34225_, _34127_, _07048_);
  and _84770_ (_34227_, _34225_, _05990_);
  and _84771_ (_34228_, _34227_, _34224_);
  and _84772_ (_34229_, _34164_, _05989_);
  or _84773_ (_34230_, _34229_, _06646_);
  or _84774_ (_34231_, _34230_, _34228_);
  and _84775_ (_34232_, _15921_, _08022_);
  or _84776_ (_34233_, _34119_, _06651_);
  or _84777_ (_34234_, _34233_, _34232_);
  and _84778_ (_34235_, _34234_, _01442_);
  and _84779_ (_34236_, _34235_, _34231_);
  or _84780_ (_34238_, _34236_, _34118_);
  and _84781_ (_44264_, _34238_, _43634_);
  and _84782_ (_34239_, _01446_, \oc8051_golden_model_1.IE [0]);
  and _84783_ (_34240_, _13804_, \oc8051_golden_model_1.IE [0]);
  nor _84784_ (_34241_, _12622_, _13804_);
  or _84785_ (_34242_, _34241_, _34240_);
  and _84786_ (_34243_, _10577_, _07986_);
  nor _84787_ (_34244_, _34243_, _07337_);
  and _84788_ (_34245_, _34244_, _34242_);
  nor _84789_ (_34246_, _08453_, _13804_);
  or _84790_ (_34248_, _34246_, _34240_);
  or _84791_ (_34249_, _34248_, _07275_);
  and _84792_ (_34250_, _07986_, \oc8051_golden_model_1.ACC [0]);
  or _84793_ (_34251_, _34250_, _34240_);
  and _84794_ (_34252_, _34251_, _07259_);
  and _84795_ (_34253_, _07260_, \oc8051_golden_model_1.IE [0]);
  or _84796_ (_34254_, _34253_, _06474_);
  or _84797_ (_34255_, _34254_, _34252_);
  and _84798_ (_34256_, _34255_, _06357_);
  and _84799_ (_34257_, _34256_, _34249_);
  and _84800_ (_34259_, _13812_, \oc8051_golden_model_1.IE [0]);
  and _84801_ (_34260_, _14581_, _08652_);
  or _84802_ (_34261_, _34260_, _34259_);
  and _84803_ (_34262_, _34261_, _06356_);
  or _84804_ (_34263_, _34262_, _34257_);
  and _84805_ (_34264_, _34263_, _06772_);
  and _84806_ (_34265_, _07986_, _07250_);
  or _84807_ (_34266_, _34265_, _34240_);
  and _84808_ (_34267_, _34266_, _06410_);
  or _84809_ (_34268_, _34267_, _06417_);
  or _84810_ (_34270_, _34268_, _34264_);
  or _84811_ (_34271_, _34251_, _06426_);
  and _84812_ (_34272_, _34271_, _06353_);
  and _84813_ (_34273_, _34272_, _34270_);
  and _84814_ (_34274_, _34240_, _06352_);
  or _84815_ (_34275_, _34274_, _06345_);
  or _84816_ (_34276_, _34275_, _34273_);
  or _84817_ (_34277_, _34248_, _06346_);
  and _84818_ (_34278_, _34277_, _06340_);
  and _84819_ (_34279_, _34278_, _34276_);
  or _84820_ (_34281_, _34259_, _16663_);
  and _84821_ (_34282_, _34281_, _06339_);
  and _84822_ (_34283_, _34282_, _34261_);
  or _84823_ (_34284_, _34283_, _10153_);
  or _84824_ (_34285_, _34284_, _34279_);
  or _84825_ (_34286_, _34266_, _06327_);
  and _84826_ (_34287_, _34286_, _34285_);
  or _84827_ (_34288_, _34287_, _09572_);
  and _84828_ (_34289_, _09447_, _07986_);
  or _84829_ (_34290_, _34240_, _06333_);
  or _84830_ (_34292_, _34290_, _34289_);
  and _84831_ (_34293_, _34292_, _06313_);
  and _84832_ (_34294_, _34293_, _34288_);
  and _84833_ (_34295_, _14666_, _07986_);
  or _84834_ (_34296_, _34295_, _34240_);
  and _84835_ (_34297_, _34296_, _06037_);
  or _84836_ (_34298_, _34297_, _06277_);
  or _84837_ (_34299_, _34298_, _34294_);
  and _84838_ (_34300_, _07986_, _09008_);
  or _84839_ (_34301_, _34300_, _34240_);
  or _84840_ (_34303_, _34301_, _06278_);
  and _84841_ (_34304_, _34303_, _34299_);
  or _84842_ (_34305_, _34304_, _06502_);
  and _84843_ (_34306_, _14566_, _07986_);
  or _84844_ (_34307_, _34240_, _07334_);
  or _84845_ (_34308_, _34307_, _34306_);
  and _84846_ (_34309_, _34308_, _07337_);
  and _84847_ (_34310_, _34309_, _34305_);
  or _84848_ (_34311_, _34310_, _34245_);
  and _84849_ (_34312_, _34311_, _07339_);
  nand _84850_ (_34314_, _34301_, _06507_);
  nor _84851_ (_34315_, _34314_, _34246_);
  or _84852_ (_34316_, _34315_, _06610_);
  or _84853_ (_34317_, _34316_, _34312_);
  or _84854_ (_34318_, _34243_, _34240_);
  or _84855_ (_34319_, _34318_, _07331_);
  and _84856_ (_34320_, _34319_, _34317_);
  or _84857_ (_34321_, _34320_, _06509_);
  and _84858_ (_34322_, _14563_, _07986_);
  or _84859_ (_34323_, _34240_, _09107_);
  or _84860_ (_34325_, _34323_, _34322_);
  and _84861_ (_34326_, _34325_, _09112_);
  and _84862_ (_34327_, _34326_, _34321_);
  and _84863_ (_34328_, _34242_, _06602_);
  or _84864_ (_34329_, _34328_, _06639_);
  or _84865_ (_34330_, _34329_, _34327_);
  or _84866_ (_34331_, _34248_, _07048_);
  and _84867_ (_34332_, _34331_, _34330_);
  or _84868_ (_34333_, _34332_, _05989_);
  or _84869_ (_34334_, _34240_, _05990_);
  and _84870_ (_34336_, _34334_, _34333_);
  or _84871_ (_34337_, _34336_, _06646_);
  or _84872_ (_34338_, _34248_, _06651_);
  and _84873_ (_34339_, _34338_, _01442_);
  and _84874_ (_34340_, _34339_, _34337_);
  or _84875_ (_34341_, _34340_, _34239_);
  and _84876_ (_44265_, _34341_, _43634_);
  not _84877_ (_34342_, \oc8051_golden_model_1.IE [1]);
  nor _84878_ (_34343_, _01442_, _34342_);
  nor _84879_ (_34344_, _07986_, _34342_);
  nor _84880_ (_34346_, _10578_, _13804_);
  or _84881_ (_34347_, _34346_, _34344_);
  or _84882_ (_34348_, _34347_, _09112_);
  or _84883_ (_34349_, _14851_, _13804_);
  or _84884_ (_34350_, _07986_, \oc8051_golden_model_1.IE [1]);
  and _84885_ (_34351_, _34350_, _06037_);
  and _84886_ (_34352_, _34351_, _34349_);
  nor _84887_ (_34353_, _13804_, _07448_);
  or _84888_ (_34354_, _34353_, _34344_);
  and _84889_ (_34355_, _34354_, _06410_);
  nor _84890_ (_34357_, _08652_, _34342_);
  and _84891_ (_34358_, _14767_, _08652_);
  or _84892_ (_34359_, _34358_, _34357_);
  or _84893_ (_34360_, _34359_, _06357_);
  and _84894_ (_34361_, _14744_, _07986_);
  not _84895_ (_34362_, _34361_);
  and _84896_ (_34363_, _34362_, _34350_);
  and _84897_ (_34364_, _34363_, _06474_);
  nor _84898_ (_34365_, _07259_, _34342_);
  and _84899_ (_34366_, _07986_, \oc8051_golden_model_1.ACC [1]);
  or _84900_ (_34368_, _34366_, _34344_);
  and _84901_ (_34369_, _34368_, _07259_);
  or _84902_ (_34370_, _34369_, _34365_);
  and _84903_ (_34371_, _34370_, _07275_);
  or _84904_ (_34372_, _34371_, _06356_);
  or _84905_ (_34373_, _34372_, _34364_);
  and _84906_ (_34374_, _34373_, _34360_);
  and _84907_ (_34375_, _34374_, _06772_);
  or _84908_ (_34376_, _34375_, _34355_);
  or _84909_ (_34377_, _34376_, _06417_);
  or _84910_ (_34379_, _34368_, _06426_);
  and _84911_ (_34380_, _34379_, _06353_);
  and _84912_ (_34381_, _34380_, _34377_);
  and _84913_ (_34382_, _14754_, _08652_);
  or _84914_ (_34383_, _34382_, _34357_);
  and _84915_ (_34384_, _34383_, _06352_);
  or _84916_ (_34385_, _34384_, _06345_);
  or _84917_ (_34386_, _34385_, _34381_);
  or _84918_ (_34387_, _34357_, _14782_);
  and _84919_ (_34388_, _34387_, _34359_);
  or _84920_ (_34390_, _34388_, _06346_);
  and _84921_ (_34391_, _34390_, _06340_);
  and _84922_ (_34392_, _34391_, _34386_);
  and _84923_ (_34393_, _14796_, _08652_);
  or _84924_ (_34394_, _34393_, _34357_);
  and _84925_ (_34395_, _34394_, _06339_);
  or _84926_ (_34396_, _34395_, _10153_);
  or _84927_ (_34397_, _34396_, _34392_);
  or _84928_ (_34398_, _34354_, _06327_);
  and _84929_ (_34399_, _34398_, _34397_);
  or _84930_ (_34401_, _34399_, _09572_);
  and _84931_ (_34402_, _09402_, _07986_);
  or _84932_ (_34403_, _34344_, _06333_);
  or _84933_ (_34404_, _34403_, _34402_);
  and _84934_ (_34405_, _34404_, _06313_);
  and _84935_ (_34406_, _34405_, _34401_);
  or _84936_ (_34407_, _34406_, _34352_);
  and _84937_ (_34408_, _34407_, _06278_);
  nand _84938_ (_34409_, _07986_, _07160_);
  and _84939_ (_34410_, _34350_, _06277_);
  and _84940_ (_34412_, _34410_, _34409_);
  or _84941_ (_34413_, _34412_, _34408_);
  and _84942_ (_34414_, _34413_, _07334_);
  or _84943_ (_34415_, _14749_, _13804_);
  and _84944_ (_34416_, _34350_, _06502_);
  and _84945_ (_34417_, _34416_, _34415_);
  or _84946_ (_34418_, _34417_, _06615_);
  or _84947_ (_34419_, _34418_, _34414_);
  nand _84948_ (_34420_, _10576_, _07986_);
  and _84949_ (_34421_, _34420_, _34347_);
  or _84950_ (_34423_, _34421_, _07337_);
  and _84951_ (_34424_, _34423_, _07339_);
  and _84952_ (_34425_, _34424_, _34419_);
  or _84953_ (_34426_, _14747_, _13804_);
  and _84954_ (_34427_, _34350_, _06507_);
  and _84955_ (_34428_, _34427_, _34426_);
  or _84956_ (_34429_, _34428_, _06610_);
  or _84957_ (_34430_, _34429_, _34425_);
  nor _84958_ (_34431_, _34344_, _07331_);
  nand _84959_ (_34432_, _34431_, _34420_);
  and _84960_ (_34434_, _34432_, _09107_);
  and _84961_ (_34435_, _34434_, _34430_);
  or _84962_ (_34436_, _34409_, _08404_);
  and _84963_ (_34437_, _34350_, _06509_);
  and _84964_ (_34438_, _34437_, _34436_);
  or _84965_ (_34439_, _34438_, _06602_);
  or _84966_ (_34440_, _34439_, _34435_);
  and _84967_ (_34441_, _34440_, _34348_);
  or _84968_ (_34442_, _34441_, _06639_);
  or _84969_ (_34443_, _34363_, _07048_);
  and _84970_ (_34445_, _34443_, _05990_);
  and _84971_ (_34446_, _34445_, _34442_);
  and _84972_ (_34447_, _34383_, _05989_);
  or _84973_ (_34448_, _34447_, _06646_);
  or _84974_ (_34449_, _34448_, _34446_);
  or _84975_ (_34450_, _34344_, _06651_);
  or _84976_ (_34451_, _34450_, _34361_);
  and _84977_ (_34452_, _34451_, _01442_);
  and _84978_ (_34453_, _34452_, _34449_);
  or _84979_ (_34454_, _34453_, _34343_);
  and _84980_ (_44267_, _34454_, _43634_);
  and _84981_ (_34456_, _01446_, \oc8051_golden_model_1.IE [2]);
  and _84982_ (_34457_, _13804_, \oc8051_golden_model_1.IE [2]);
  nor _84983_ (_34458_, _10582_, _13804_);
  or _84984_ (_34459_, _34458_, _34457_);
  and _84985_ (_34460_, _07986_, \oc8051_golden_model_1.ACC [2]);
  nand _84986_ (_34461_, _34460_, _08503_);
  and _84987_ (_34462_, _34461_, _06615_);
  and _84988_ (_34463_, _34462_, _34459_);
  nor _84989_ (_34464_, _13804_, _07854_);
  or _84990_ (_34466_, _34464_, _34457_);
  or _84991_ (_34467_, _34466_, _06327_);
  or _84992_ (_34468_, _34466_, _06772_);
  and _84993_ (_34469_, _14959_, _07986_);
  or _84994_ (_34470_, _34469_, _34457_);
  or _84995_ (_34471_, _34470_, _07275_);
  or _84996_ (_34472_, _34460_, _34457_);
  and _84997_ (_34473_, _34472_, _07259_);
  and _84998_ (_34474_, _07260_, \oc8051_golden_model_1.IE [2]);
  or _84999_ (_34475_, _34474_, _06474_);
  or _85000_ (_34477_, _34475_, _34473_);
  and _85001_ (_34478_, _34477_, _06357_);
  and _85002_ (_34479_, _34478_, _34471_);
  and _85003_ (_34480_, _13812_, \oc8051_golden_model_1.IE [2]);
  and _85004_ (_34481_, _14955_, _08652_);
  or _85005_ (_34482_, _34481_, _34480_);
  and _85006_ (_34483_, _34482_, _06356_);
  or _85007_ (_34484_, _34483_, _06410_);
  or _85008_ (_34485_, _34484_, _34479_);
  and _85009_ (_34486_, _34485_, _34468_);
  or _85010_ (_34488_, _34486_, _06417_);
  or _85011_ (_34489_, _34472_, _06426_);
  and _85012_ (_34490_, _34489_, _06353_);
  and _85013_ (_34491_, _34490_, _34488_);
  and _85014_ (_34492_, _14953_, _08652_);
  or _85015_ (_34493_, _34492_, _34480_);
  and _85016_ (_34494_, _34493_, _06352_);
  or _85017_ (_34495_, _34494_, _06345_);
  or _85018_ (_34496_, _34495_, _34491_);
  and _85019_ (_34497_, _34481_, _14986_);
  or _85020_ (_34499_, _34480_, _06346_);
  or _85021_ (_34500_, _34499_, _34497_);
  and _85022_ (_34501_, _34500_, _06340_);
  and _85023_ (_34502_, _34501_, _34496_);
  and _85024_ (_34503_, _15000_, _08652_);
  or _85025_ (_34504_, _34503_, _34480_);
  and _85026_ (_34505_, _34504_, _06339_);
  or _85027_ (_34506_, _34505_, _10153_);
  or _85028_ (_34507_, _34506_, _34502_);
  and _85029_ (_34508_, _34507_, _34467_);
  or _85030_ (_34510_, _34508_, _09572_);
  and _85031_ (_34511_, _09356_, _07986_);
  or _85032_ (_34512_, _34457_, _06333_);
  or _85033_ (_34513_, _34512_, _34511_);
  and _85034_ (_34514_, _34513_, _06313_);
  and _85035_ (_34515_, _34514_, _34510_);
  and _85036_ (_34516_, _15056_, _07986_);
  or _85037_ (_34517_, _34516_, _34457_);
  and _85038_ (_34518_, _34517_, _06037_);
  or _85039_ (_34519_, _34518_, _06277_);
  or _85040_ (_34521_, _34519_, _34515_);
  and _85041_ (_34522_, _07986_, _09057_);
  or _85042_ (_34523_, _34522_, _34457_);
  or _85043_ (_34524_, _34523_, _06278_);
  and _85044_ (_34525_, _34524_, _34521_);
  or _85045_ (_34526_, _34525_, _06502_);
  and _85046_ (_34527_, _14948_, _07986_);
  or _85047_ (_34528_, _34457_, _07334_);
  or _85048_ (_34529_, _34528_, _34527_);
  and _85049_ (_34530_, _34529_, _07337_);
  and _85050_ (_34532_, _34530_, _34526_);
  or _85051_ (_34533_, _34532_, _34463_);
  and _85052_ (_34534_, _34533_, _07339_);
  or _85053_ (_34535_, _34457_, _08503_);
  and _85054_ (_34536_, _34523_, _06507_);
  and _85055_ (_34537_, _34536_, _34535_);
  or _85056_ (_34538_, _34537_, _34534_);
  and _85057_ (_34539_, _34538_, _07331_);
  and _85058_ (_34540_, _34472_, _06610_);
  and _85059_ (_34541_, _34540_, _34535_);
  or _85060_ (_34543_, _34541_, _06509_);
  or _85061_ (_34544_, _34543_, _34539_);
  and _85062_ (_34545_, _14945_, _07986_);
  or _85063_ (_34546_, _34457_, _09107_);
  or _85064_ (_34547_, _34546_, _34545_);
  and _85065_ (_34548_, _34547_, _09112_);
  and _85066_ (_34549_, _34548_, _34544_);
  and _85067_ (_34550_, _34459_, _06602_);
  or _85068_ (_34551_, _34550_, _06639_);
  or _85069_ (_34552_, _34551_, _34549_);
  or _85070_ (_34554_, _34470_, _07048_);
  and _85071_ (_34555_, _34554_, _05990_);
  and _85072_ (_34556_, _34555_, _34552_);
  and _85073_ (_34557_, _34493_, _05989_);
  or _85074_ (_34558_, _34557_, _06646_);
  or _85075_ (_34559_, _34558_, _34556_);
  and _85076_ (_34560_, _15129_, _07986_);
  or _85077_ (_34561_, _34457_, _06651_);
  or _85078_ (_34562_, _34561_, _34560_);
  and _85079_ (_34563_, _34562_, _01442_);
  and _85080_ (_34565_, _34563_, _34559_);
  or _85081_ (_34566_, _34565_, _34456_);
  and _85082_ (_44268_, _34566_, _43634_);
  and _85083_ (_34567_, _01446_, \oc8051_golden_model_1.IE [3]);
  and _85084_ (_34568_, _13804_, \oc8051_golden_model_1.IE [3]);
  nor _85085_ (_34569_, _13804_, _07680_);
  or _85086_ (_34570_, _34569_, _34568_);
  or _85087_ (_34571_, _34570_, _06327_);
  and _85088_ (_34572_, _15153_, _07986_);
  or _85089_ (_34573_, _34572_, _34568_);
  or _85090_ (_34575_, _34573_, _07275_);
  and _85091_ (_34576_, _07986_, \oc8051_golden_model_1.ACC [3]);
  or _85092_ (_34577_, _34576_, _34568_);
  and _85093_ (_34578_, _34577_, _07259_);
  and _85094_ (_34579_, _07260_, \oc8051_golden_model_1.IE [3]);
  or _85095_ (_34580_, _34579_, _06474_);
  or _85096_ (_34581_, _34580_, _34578_);
  and _85097_ (_34582_, _34581_, _06357_);
  and _85098_ (_34583_, _34582_, _34575_);
  and _85099_ (_34584_, _13812_, \oc8051_golden_model_1.IE [3]);
  and _85100_ (_34586_, _15150_, _08652_);
  or _85101_ (_34587_, _34586_, _34584_);
  and _85102_ (_34588_, _34587_, _06356_);
  or _85103_ (_34589_, _34588_, _06410_);
  or _85104_ (_34590_, _34589_, _34583_);
  or _85105_ (_34591_, _34570_, _06772_);
  and _85106_ (_34592_, _34591_, _34590_);
  or _85107_ (_34593_, _34592_, _06417_);
  or _85108_ (_34594_, _34577_, _06426_);
  and _85109_ (_34595_, _34594_, _06353_);
  and _85110_ (_34597_, _34595_, _34593_);
  and _85111_ (_34598_, _15148_, _08652_);
  or _85112_ (_34599_, _34598_, _34584_);
  and _85113_ (_34600_, _34599_, _06352_);
  or _85114_ (_34601_, _34600_, _06345_);
  or _85115_ (_34602_, _34601_, _34597_);
  or _85116_ (_34603_, _34584_, _15180_);
  and _85117_ (_34604_, _34603_, _34587_);
  or _85118_ (_34605_, _34604_, _06346_);
  and _85119_ (_34606_, _34605_, _06340_);
  and _85120_ (_34608_, _34606_, _34602_);
  and _85121_ (_34609_, _15197_, _08652_);
  or _85122_ (_34610_, _34609_, _34584_);
  and _85123_ (_34611_, _34610_, _06339_);
  or _85124_ (_34612_, _34611_, _10153_);
  or _85125_ (_34613_, _34612_, _34608_);
  and _85126_ (_34614_, _34613_, _34571_);
  or _85127_ (_34615_, _34614_, _09572_);
  and _85128_ (_34616_, _09310_, _07986_);
  or _85129_ (_34617_, _34568_, _06333_);
  or _85130_ (_34619_, _34617_, _34616_);
  and _85131_ (_34620_, _34619_, _06313_);
  and _85132_ (_34621_, _34620_, _34615_);
  and _85133_ (_34622_, _15251_, _07986_);
  or _85134_ (_34623_, _34622_, _34568_);
  and _85135_ (_34624_, _34623_, _06037_);
  or _85136_ (_34625_, _34624_, _06277_);
  or _85137_ (_34626_, _34625_, _34621_);
  and _85138_ (_34627_, _07986_, _09014_);
  or _85139_ (_34628_, _34627_, _34568_);
  or _85140_ (_34629_, _34628_, _06278_);
  and _85141_ (_34630_, _34629_, _34626_);
  or _85142_ (_34631_, _34630_, _06502_);
  and _85143_ (_34632_, _15266_, _07986_);
  or _85144_ (_34633_, _34568_, _07334_);
  or _85145_ (_34634_, _34633_, _34632_);
  and _85146_ (_34635_, _34634_, _07337_);
  and _85147_ (_34636_, _34635_, _34631_);
  and _85148_ (_34637_, _12619_, _07986_);
  or _85149_ (_34638_, _34637_, _34568_);
  and _85150_ (_34640_, _34638_, _06615_);
  or _85151_ (_34641_, _34640_, _34636_);
  and _85152_ (_34642_, _34641_, _07339_);
  or _85153_ (_34643_, _34568_, _08359_);
  and _85154_ (_34644_, _34628_, _06507_);
  and _85155_ (_34645_, _34644_, _34643_);
  or _85156_ (_34646_, _34645_, _34642_);
  and _85157_ (_34647_, _34646_, _07331_);
  and _85158_ (_34648_, _34577_, _06610_);
  and _85159_ (_34649_, _34648_, _34643_);
  or _85160_ (_34651_, _34649_, _06509_);
  or _85161_ (_34652_, _34651_, _34647_);
  and _85162_ (_34653_, _15263_, _07986_);
  or _85163_ (_34654_, _34568_, _09107_);
  or _85164_ (_34655_, _34654_, _34653_);
  and _85165_ (_34656_, _34655_, _09112_);
  and _85166_ (_34657_, _34656_, _34652_);
  nor _85167_ (_34658_, _10574_, _13804_);
  or _85168_ (_34659_, _34658_, _34568_);
  and _85169_ (_34660_, _34659_, _06602_);
  or _85170_ (_34662_, _34660_, _06639_);
  or _85171_ (_34663_, _34662_, _34657_);
  or _85172_ (_34664_, _34573_, _07048_);
  and _85173_ (_34665_, _34664_, _05990_);
  and _85174_ (_34666_, _34665_, _34663_);
  and _85175_ (_34667_, _34599_, _05989_);
  or _85176_ (_34668_, _34667_, _06646_);
  or _85177_ (_34669_, _34668_, _34666_);
  and _85178_ (_34670_, _15321_, _07986_);
  or _85179_ (_34671_, _34568_, _06651_);
  or _85180_ (_34673_, _34671_, _34670_);
  and _85181_ (_34674_, _34673_, _01442_);
  and _85182_ (_34675_, _34674_, _34669_);
  or _85183_ (_34676_, _34675_, _34567_);
  and _85184_ (_44269_, _34676_, _43634_);
  and _85185_ (_34677_, _01446_, \oc8051_golden_model_1.IE [4]);
  and _85186_ (_34678_, _13804_, \oc8051_golden_model_1.IE [4]);
  nor _85187_ (_34679_, _08596_, _13804_);
  or _85188_ (_34680_, _34679_, _34678_);
  or _85189_ (_34681_, _34680_, _06327_);
  and _85190_ (_34683_, _13812_, \oc8051_golden_model_1.IE [4]);
  and _85191_ (_34684_, _15348_, _08652_);
  or _85192_ (_34685_, _34684_, _34683_);
  and _85193_ (_34686_, _34685_, _06352_);
  and _85194_ (_34687_, _15367_, _07986_);
  or _85195_ (_34688_, _34687_, _34678_);
  or _85196_ (_34689_, _34688_, _07275_);
  and _85197_ (_34690_, _07986_, \oc8051_golden_model_1.ACC [4]);
  or _85198_ (_34691_, _34690_, _34678_);
  and _85199_ (_34692_, _34691_, _07259_);
  and _85200_ (_34694_, _07260_, \oc8051_golden_model_1.IE [4]);
  or _85201_ (_34695_, _34694_, _06474_);
  or _85202_ (_34696_, _34695_, _34692_);
  and _85203_ (_34697_, _34696_, _06357_);
  and _85204_ (_34698_, _34697_, _34689_);
  and _85205_ (_34699_, _15353_, _08652_);
  or _85206_ (_34700_, _34699_, _34683_);
  and _85207_ (_34701_, _34700_, _06356_);
  or _85208_ (_34702_, _34701_, _06410_);
  or _85209_ (_34703_, _34702_, _34698_);
  or _85210_ (_34705_, _34680_, _06772_);
  and _85211_ (_34706_, _34705_, _34703_);
  or _85212_ (_34707_, _34706_, _06417_);
  or _85213_ (_34708_, _34691_, _06426_);
  and _85214_ (_34709_, _34708_, _06353_);
  and _85215_ (_34710_, _34709_, _34707_);
  or _85216_ (_34711_, _34710_, _34686_);
  and _85217_ (_34712_, _34711_, _06346_);
  and _85218_ (_34713_, _15385_, _08652_);
  or _85219_ (_34714_, _34713_, _34683_);
  and _85220_ (_34716_, _34714_, _06345_);
  or _85221_ (_34717_, _34716_, _34712_);
  and _85222_ (_34718_, _34717_, _06340_);
  and _85223_ (_34719_, _15350_, _08652_);
  or _85224_ (_34720_, _34719_, _34683_);
  and _85225_ (_34721_, _34720_, _06339_);
  or _85226_ (_34722_, _34721_, _10153_);
  or _85227_ (_34723_, _34722_, _34718_);
  and _85228_ (_34724_, _34723_, _34681_);
  or _85229_ (_34725_, _34724_, _09572_);
  and _85230_ (_34727_, _09264_, _07986_);
  or _85231_ (_34728_, _34678_, _06333_);
  or _85232_ (_34729_, _34728_, _34727_);
  and _85233_ (_34730_, _34729_, _06313_);
  and _85234_ (_34731_, _34730_, _34725_);
  and _85235_ (_34732_, _15452_, _07986_);
  or _85236_ (_34733_, _34732_, _34678_);
  and _85237_ (_34734_, _34733_, _06037_);
  or _85238_ (_34735_, _34734_, _06277_);
  or _85239_ (_34736_, _34735_, _34731_);
  and _85240_ (_34738_, _08995_, _07986_);
  or _85241_ (_34739_, _34738_, _34678_);
  or _85242_ (_34740_, _34739_, _06278_);
  and _85243_ (_34741_, _34740_, _34736_);
  or _85244_ (_34742_, _34741_, _06502_);
  and _85245_ (_34743_, _15345_, _07986_);
  or _85246_ (_34744_, _34678_, _07334_);
  or _85247_ (_34745_, _34744_, _34743_);
  and _85248_ (_34746_, _34745_, _07337_);
  and _85249_ (_34747_, _34746_, _34742_);
  and _85250_ (_34749_, _10590_, _07986_);
  or _85251_ (_34750_, _34749_, _34678_);
  and _85252_ (_34751_, _34750_, _06615_);
  or _85253_ (_34752_, _34751_, _34747_);
  and _85254_ (_34753_, _34752_, _07339_);
  or _85255_ (_34754_, _34678_, _08599_);
  and _85256_ (_34755_, _34739_, _06507_);
  and _85257_ (_34756_, _34755_, _34754_);
  or _85258_ (_34757_, _34756_, _34753_);
  and _85259_ (_34758_, _34757_, _07331_);
  and _85260_ (_34760_, _34691_, _06610_);
  and _85261_ (_34761_, _34760_, _34754_);
  or _85262_ (_34762_, _34761_, _06509_);
  or _85263_ (_34763_, _34762_, _34758_);
  and _85264_ (_34764_, _15342_, _07986_);
  or _85265_ (_34765_, _34678_, _09107_);
  or _85266_ (_34766_, _34765_, _34764_);
  and _85267_ (_34767_, _34766_, _09112_);
  and _85268_ (_34768_, _34767_, _34763_);
  nor _85269_ (_34769_, _10589_, _13804_);
  or _85270_ (_34771_, _34769_, _34678_);
  and _85271_ (_34772_, _34771_, _06602_);
  or _85272_ (_34773_, _34772_, _06639_);
  or _85273_ (_34774_, _34773_, _34768_);
  or _85274_ (_34775_, _34688_, _07048_);
  and _85275_ (_34776_, _34775_, _05990_);
  and _85276_ (_34777_, _34776_, _34774_);
  and _85277_ (_34778_, _34685_, _05989_);
  or _85278_ (_34779_, _34778_, _06646_);
  or _85279_ (_34780_, _34779_, _34777_);
  and _85280_ (_34782_, _15524_, _07986_);
  or _85281_ (_34783_, _34678_, _06651_);
  or _85282_ (_34784_, _34783_, _34782_);
  and _85283_ (_34785_, _34784_, _01442_);
  and _85284_ (_34786_, _34785_, _34780_);
  or _85285_ (_34787_, _34786_, _34677_);
  and _85286_ (_44270_, _34787_, _43634_);
  and _85287_ (_34788_, _01446_, \oc8051_golden_model_1.IE [5]);
  and _85288_ (_34789_, _13804_, \oc8051_golden_model_1.IE [5]);
  nor _85289_ (_34790_, _10570_, _13804_);
  or _85290_ (_34792_, _34790_, _34789_);
  and _85291_ (_34793_, _07986_, \oc8051_golden_model_1.ACC [5]);
  nand _85292_ (_34794_, _34793_, _08308_);
  and _85293_ (_34795_, _34794_, _06615_);
  and _85294_ (_34796_, _34795_, _34792_);
  and _85295_ (_34797_, _15550_, _07986_);
  or _85296_ (_34798_, _34797_, _34789_);
  or _85297_ (_34799_, _34798_, _07275_);
  or _85298_ (_34800_, _34793_, _34789_);
  and _85299_ (_34801_, _34800_, _07259_);
  and _85300_ (_34803_, _07260_, \oc8051_golden_model_1.IE [5]);
  or _85301_ (_34804_, _34803_, _06474_);
  or _85302_ (_34805_, _34804_, _34801_);
  and _85303_ (_34806_, _34805_, _06357_);
  and _85304_ (_34807_, _34806_, _34799_);
  and _85305_ (_34808_, _13812_, \oc8051_golden_model_1.IE [5]);
  and _85306_ (_34809_, _15566_, _08652_);
  or _85307_ (_34810_, _34809_, _34808_);
  and _85308_ (_34811_, _34810_, _06356_);
  or _85309_ (_34812_, _34811_, _06410_);
  or _85310_ (_34814_, _34812_, _34807_);
  nor _85311_ (_34815_, _08305_, _13804_);
  or _85312_ (_34816_, _34815_, _34789_);
  or _85313_ (_34817_, _34816_, _06772_);
  and _85314_ (_34818_, _34817_, _34814_);
  or _85315_ (_34819_, _34818_, _06417_);
  or _85316_ (_34820_, _34800_, _06426_);
  and _85317_ (_34821_, _34820_, _06353_);
  and _85318_ (_34822_, _34821_, _34819_);
  and _85319_ (_34823_, _15544_, _08652_);
  or _85320_ (_34825_, _34823_, _34808_);
  and _85321_ (_34826_, _34825_, _06352_);
  or _85322_ (_34827_, _34826_, _06345_);
  or _85323_ (_34828_, _34827_, _34822_);
  or _85324_ (_34829_, _34808_, _15581_);
  and _85325_ (_34830_, _34829_, _34810_);
  or _85326_ (_34831_, _34830_, _06346_);
  and _85327_ (_34832_, _34831_, _06340_);
  and _85328_ (_34833_, _34832_, _34828_);
  and _85329_ (_34834_, _15546_, _08652_);
  or _85330_ (_34836_, _34834_, _34808_);
  and _85331_ (_34837_, _34836_, _06339_);
  or _85332_ (_34838_, _34837_, _10153_);
  or _85333_ (_34839_, _34838_, _34833_);
  or _85334_ (_34840_, _34816_, _06327_);
  and _85335_ (_34841_, _34840_, _34839_);
  or _85336_ (_34842_, _34841_, _09572_);
  and _85337_ (_34843_, _09218_, _07986_);
  or _85338_ (_34844_, _34789_, _06333_);
  or _85339_ (_34845_, _34844_, _34843_);
  and _85340_ (_34847_, _34845_, _06313_);
  and _85341_ (_34848_, _34847_, _34842_);
  and _85342_ (_34849_, _15649_, _07986_);
  or _85343_ (_34850_, _34849_, _34789_);
  and _85344_ (_34851_, _34850_, _06037_);
  or _85345_ (_34852_, _34851_, _06277_);
  or _85346_ (_34853_, _34852_, _34848_);
  and _85347_ (_34854_, _08954_, _07986_);
  or _85348_ (_34855_, _34854_, _34789_);
  or _85349_ (_34856_, _34855_, _06278_);
  and _85350_ (_34858_, _34856_, _34853_);
  or _85351_ (_34859_, _34858_, _06502_);
  and _85352_ (_34860_, _15664_, _07986_);
  or _85353_ (_34861_, _34789_, _07334_);
  or _85354_ (_34862_, _34861_, _34860_);
  and _85355_ (_34863_, _34862_, _07337_);
  and _85356_ (_34864_, _34863_, _34859_);
  or _85357_ (_34865_, _34864_, _34796_);
  and _85358_ (_34866_, _34865_, _07339_);
  or _85359_ (_34867_, _34789_, _08308_);
  and _85360_ (_34869_, _34855_, _06507_);
  and _85361_ (_34870_, _34869_, _34867_);
  or _85362_ (_34871_, _34870_, _34866_);
  and _85363_ (_34872_, _34871_, _07331_);
  and _85364_ (_34873_, _34800_, _06610_);
  and _85365_ (_34874_, _34873_, _34867_);
  or _85366_ (_34875_, _34874_, _06509_);
  or _85367_ (_34876_, _34875_, _34872_);
  and _85368_ (_34877_, _15663_, _07986_);
  or _85369_ (_34878_, _34789_, _09107_);
  or _85370_ (_34880_, _34878_, _34877_);
  and _85371_ (_34881_, _34880_, _09112_);
  and _85372_ (_34882_, _34881_, _34876_);
  and _85373_ (_34883_, _34792_, _06602_);
  or _85374_ (_34884_, _34883_, _06639_);
  or _85375_ (_34885_, _34884_, _34882_);
  or _85376_ (_34886_, _34798_, _07048_);
  and _85377_ (_34887_, _34886_, _05990_);
  and _85378_ (_34888_, _34887_, _34885_);
  and _85379_ (_34889_, _34825_, _05989_);
  or _85380_ (_34891_, _34889_, _06646_);
  or _85381_ (_34892_, _34891_, _34888_);
  and _85382_ (_34893_, _15721_, _07986_);
  or _85383_ (_34894_, _34789_, _06651_);
  or _85384_ (_34895_, _34894_, _34893_);
  and _85385_ (_34896_, _34895_, _01442_);
  and _85386_ (_34897_, _34896_, _34892_);
  or _85387_ (_34898_, _34897_, _34788_);
  and _85388_ (_44271_, _34898_, _43634_);
  and _85389_ (_34899_, _01446_, \oc8051_golden_model_1.IE [6]);
  and _85390_ (_34901_, _13804_, \oc8051_golden_model_1.IE [6]);
  and _85391_ (_34902_, _15759_, _07986_);
  or _85392_ (_34903_, _34902_, _34901_);
  or _85393_ (_34904_, _34903_, _07275_);
  and _85394_ (_34905_, _07986_, \oc8051_golden_model_1.ACC [6]);
  or _85395_ (_34906_, _34905_, _34901_);
  and _85396_ (_34907_, _34906_, _07259_);
  and _85397_ (_34908_, _07260_, \oc8051_golden_model_1.IE [6]);
  or _85398_ (_34909_, _34908_, _06474_);
  or _85399_ (_34910_, _34909_, _34907_);
  and _85400_ (_34912_, _34910_, _06357_);
  and _85401_ (_34913_, _34912_, _34904_);
  and _85402_ (_34914_, _13812_, \oc8051_golden_model_1.IE [6]);
  and _85403_ (_34915_, _15763_, _08652_);
  or _85404_ (_34916_, _34915_, _34914_);
  and _85405_ (_34917_, _34916_, _06356_);
  or _85406_ (_34918_, _34917_, _06410_);
  or _85407_ (_34919_, _34918_, _34913_);
  nor _85408_ (_34920_, _08209_, _13804_);
  or _85409_ (_34921_, _34920_, _34901_);
  or _85410_ (_34923_, _34921_, _06772_);
  and _85411_ (_34924_, _34923_, _34919_);
  or _85412_ (_34925_, _34924_, _06417_);
  or _85413_ (_34926_, _34906_, _06426_);
  and _85414_ (_34927_, _34926_, _06353_);
  and _85415_ (_34928_, _34927_, _34925_);
  and _85416_ (_34929_, _15743_, _08652_);
  or _85417_ (_34930_, _34929_, _34914_);
  and _85418_ (_34931_, _34930_, _06352_);
  or _85419_ (_34932_, _34931_, _06345_);
  or _85420_ (_34934_, _34932_, _34928_);
  or _85421_ (_34935_, _34914_, _15778_);
  and _85422_ (_34936_, _34935_, _34916_);
  or _85423_ (_34937_, _34936_, _06346_);
  and _85424_ (_34938_, _34937_, _06340_);
  and _85425_ (_34939_, _34938_, _34934_);
  and _85426_ (_34940_, _15745_, _08652_);
  or _85427_ (_34941_, _34940_, _34914_);
  and _85428_ (_34942_, _34941_, _06339_);
  or _85429_ (_34943_, _34942_, _10153_);
  or _85430_ (_34945_, _34943_, _34939_);
  or _85431_ (_34946_, _34921_, _06327_);
  and _85432_ (_34947_, _34946_, _34945_);
  or _85433_ (_34948_, _34947_, _09572_);
  and _85434_ (_34949_, _09172_, _07986_);
  or _85435_ (_34950_, _34901_, _06333_);
  or _85436_ (_34951_, _34950_, _34949_);
  and _85437_ (_34952_, _34951_, _06313_);
  and _85438_ (_34953_, _34952_, _34948_);
  and _85439_ (_34954_, _15846_, _07986_);
  or _85440_ (_34956_, _34954_, _34901_);
  and _85441_ (_34957_, _34956_, _06037_);
  or _85442_ (_34958_, _34957_, _06277_);
  or _85443_ (_34959_, _34958_, _34953_);
  and _85444_ (_34960_, _15853_, _07986_);
  or _85445_ (_34961_, _34960_, _34901_);
  or _85446_ (_34962_, _34961_, _06278_);
  and _85447_ (_34963_, _34962_, _34959_);
  or _85448_ (_34964_, _34963_, _06502_);
  and _85449_ (_34965_, _15862_, _07986_);
  or _85450_ (_34967_, _34901_, _07334_);
  or _85451_ (_34968_, _34967_, _34965_);
  and _85452_ (_34969_, _34968_, _07337_);
  and _85453_ (_34970_, _34969_, _34964_);
  and _85454_ (_34971_, _10596_, _07986_);
  or _85455_ (_34972_, _34971_, _34901_);
  and _85456_ (_34973_, _34972_, _06615_);
  or _85457_ (_34974_, _34973_, _34970_);
  and _85458_ (_34975_, _34974_, _07339_);
  or _85459_ (_34976_, _34901_, _08212_);
  and _85460_ (_34978_, _34961_, _06507_);
  and _85461_ (_34979_, _34978_, _34976_);
  or _85462_ (_34980_, _34979_, _34975_);
  and _85463_ (_34981_, _34980_, _07331_);
  and _85464_ (_34982_, _34906_, _06610_);
  and _85465_ (_34983_, _34982_, _34976_);
  or _85466_ (_34984_, _34983_, _06509_);
  or _85467_ (_34985_, _34984_, _34981_);
  and _85468_ (_34986_, _15859_, _07986_);
  or _85469_ (_34987_, _34901_, _09107_);
  or _85470_ (_34989_, _34987_, _34986_);
  and _85471_ (_34990_, _34989_, _09112_);
  and _85472_ (_34991_, _34990_, _34985_);
  nor _85473_ (_34992_, _10595_, _13804_);
  or _85474_ (_34993_, _34992_, _34901_);
  and _85475_ (_34994_, _34993_, _06602_);
  or _85476_ (_34995_, _34994_, _06639_);
  or _85477_ (_34996_, _34995_, _34991_);
  or _85478_ (_34997_, _34903_, _07048_);
  and _85479_ (_34998_, _34997_, _05990_);
  and _85480_ (_35000_, _34998_, _34996_);
  and _85481_ (_35001_, _34930_, _05989_);
  or _85482_ (_35002_, _35001_, _06646_);
  or _85483_ (_35003_, _35002_, _35000_);
  and _85484_ (_35004_, _15921_, _07986_);
  or _85485_ (_35005_, _34901_, _06651_);
  or _85486_ (_35006_, _35005_, _35004_);
  and _85487_ (_35007_, _35006_, _01442_);
  and _85488_ (_35008_, _35007_, _35003_);
  or _85489_ (_35009_, _35008_, _34899_);
  and _85490_ (_44272_, _35009_, _43634_);
  and _85491_ (_35011_, _01446_, \oc8051_golden_model_1.SCON [0]);
  and _85492_ (_35012_, _13907_, \oc8051_golden_model_1.SCON [0]);
  nor _85493_ (_35013_, _12622_, _13907_);
  or _85494_ (_35014_, _35013_, _35012_);
  and _85495_ (_35015_, _10577_, _07969_);
  nor _85496_ (_35016_, _35015_, _07337_);
  and _85497_ (_35017_, _35016_, _35014_);
  nor _85498_ (_35018_, _08453_, _13907_);
  or _85499_ (_35019_, _35018_, _35012_);
  or _85500_ (_35021_, _35019_, _07275_);
  and _85501_ (_35022_, _07969_, \oc8051_golden_model_1.ACC [0]);
  or _85502_ (_35023_, _35022_, _35012_);
  and _85503_ (_35024_, _35023_, _07259_);
  and _85504_ (_35025_, _07260_, \oc8051_golden_model_1.SCON [0]);
  or _85505_ (_35026_, _35025_, _06474_);
  or _85506_ (_35027_, _35026_, _35024_);
  and _85507_ (_35028_, _35027_, _06357_);
  and _85508_ (_35029_, _35028_, _35021_);
  and _85509_ (_35030_, _13915_, \oc8051_golden_model_1.SCON [0]);
  and _85510_ (_35032_, _14581_, _08650_);
  or _85511_ (_35033_, _35032_, _35030_);
  and _85512_ (_35034_, _35033_, _06356_);
  or _85513_ (_35035_, _35034_, _35029_);
  and _85514_ (_35036_, _35035_, _06772_);
  and _85515_ (_35037_, _07969_, _07250_);
  or _85516_ (_35038_, _35037_, _35012_);
  and _85517_ (_35039_, _35038_, _06410_);
  or _85518_ (_35040_, _35039_, _06417_);
  or _85519_ (_35041_, _35040_, _35036_);
  or _85520_ (_35043_, _35023_, _06426_);
  and _85521_ (_35044_, _35043_, _06353_);
  and _85522_ (_35045_, _35044_, _35041_);
  and _85523_ (_35046_, _35012_, _06352_);
  or _85524_ (_35047_, _35046_, _06345_);
  or _85525_ (_35048_, _35047_, _35045_);
  or _85526_ (_35049_, _35019_, _06346_);
  and _85527_ (_35050_, _35049_, _06340_);
  and _85528_ (_35051_, _35050_, _35048_);
  or _85529_ (_35052_, _35030_, _16663_);
  and _85530_ (_35054_, _35052_, _06339_);
  and _85531_ (_35055_, _35054_, _35033_);
  or _85532_ (_35056_, _35055_, _10153_);
  or _85533_ (_35057_, _35056_, _35051_);
  or _85534_ (_35058_, _35038_, _06327_);
  and _85535_ (_35059_, _35058_, _35057_);
  or _85536_ (_35060_, _35059_, _09572_);
  and _85537_ (_35061_, _09447_, _07969_);
  or _85538_ (_35062_, _35012_, _06333_);
  or _85539_ (_35063_, _35062_, _35061_);
  and _85540_ (_35065_, _35063_, _06313_);
  and _85541_ (_35066_, _35065_, _35060_);
  and _85542_ (_35067_, _14666_, _07969_);
  or _85543_ (_35068_, _35067_, _35012_);
  and _85544_ (_35069_, _35068_, _06037_);
  or _85545_ (_35070_, _35069_, _06277_);
  or _85546_ (_35071_, _35070_, _35066_);
  and _85547_ (_35072_, _07969_, _09008_);
  or _85548_ (_35073_, _35072_, _35012_);
  or _85549_ (_35074_, _35073_, _06278_);
  and _85550_ (_35076_, _35074_, _35071_);
  or _85551_ (_35077_, _35076_, _06502_);
  and _85552_ (_35078_, _14566_, _07969_);
  or _85553_ (_35079_, _35012_, _07334_);
  or _85554_ (_35080_, _35079_, _35078_);
  and _85555_ (_35081_, _35080_, _07337_);
  and _85556_ (_35082_, _35081_, _35077_);
  or _85557_ (_35083_, _35082_, _35017_);
  and _85558_ (_35084_, _35083_, _07339_);
  nand _85559_ (_35085_, _35073_, _06507_);
  nor _85560_ (_35087_, _35085_, _35018_);
  or _85561_ (_35088_, _35087_, _06610_);
  or _85562_ (_35089_, _35088_, _35084_);
  or _85563_ (_35090_, _35015_, _35012_);
  or _85564_ (_35091_, _35090_, _07331_);
  and _85565_ (_35092_, _35091_, _35089_);
  or _85566_ (_35093_, _35092_, _06509_);
  and _85567_ (_35094_, _14563_, _07969_);
  or _85568_ (_35095_, _35012_, _09107_);
  or _85569_ (_35096_, _35095_, _35094_);
  and _85570_ (_35098_, _35096_, _09112_);
  and _85571_ (_35099_, _35098_, _35093_);
  and _85572_ (_35100_, _35014_, _06602_);
  or _85573_ (_35101_, _35100_, _06639_);
  or _85574_ (_35102_, _35101_, _35099_);
  or _85575_ (_35103_, _35019_, _07048_);
  and _85576_ (_35104_, _35103_, _35102_);
  or _85577_ (_35105_, _35104_, _05989_);
  or _85578_ (_35106_, _35012_, _05990_);
  and _85579_ (_35107_, _35106_, _35105_);
  or _85580_ (_35109_, _35107_, _06646_);
  or _85581_ (_35110_, _35019_, _06651_);
  and _85582_ (_35111_, _35110_, _01442_);
  and _85583_ (_35112_, _35111_, _35109_);
  or _85584_ (_35113_, _35112_, _35011_);
  and _85585_ (_44274_, _35113_, _43634_);
  and _85586_ (_35114_, _01446_, \oc8051_golden_model_1.SCON [1]);
  and _85587_ (_35115_, _13907_, \oc8051_golden_model_1.SCON [1]);
  nor _85588_ (_35116_, _10578_, _13907_);
  or _85589_ (_35117_, _35116_, _35115_);
  or _85590_ (_35119_, _35117_, _09112_);
  nand _85591_ (_35120_, _07969_, _07160_);
  or _85592_ (_35121_, _07969_, \oc8051_golden_model_1.SCON [1]);
  and _85593_ (_35122_, _35121_, _06277_);
  and _85594_ (_35123_, _35122_, _35120_);
  nor _85595_ (_35124_, _13907_, _07448_);
  or _85596_ (_35125_, _35124_, _35115_);
  or _85597_ (_35126_, _35125_, _06772_);
  and _85598_ (_35127_, _14744_, _07969_);
  not _85599_ (_35128_, _35127_);
  and _85600_ (_35130_, _35128_, _35121_);
  or _85601_ (_35131_, _35130_, _07275_);
  and _85602_ (_35132_, _07969_, \oc8051_golden_model_1.ACC [1]);
  or _85603_ (_35133_, _35132_, _35115_);
  and _85604_ (_35134_, _35133_, _07259_);
  and _85605_ (_35135_, _07260_, \oc8051_golden_model_1.SCON [1]);
  or _85606_ (_35136_, _35135_, _06474_);
  or _85607_ (_35137_, _35136_, _35134_);
  and _85608_ (_35138_, _35137_, _06357_);
  and _85609_ (_35139_, _35138_, _35131_);
  and _85610_ (_35141_, _13915_, \oc8051_golden_model_1.SCON [1]);
  and _85611_ (_35142_, _14767_, _08650_);
  or _85612_ (_35143_, _35142_, _35141_);
  and _85613_ (_35144_, _35143_, _06356_);
  or _85614_ (_35145_, _35144_, _06410_);
  or _85615_ (_35146_, _35145_, _35139_);
  and _85616_ (_35147_, _35146_, _35126_);
  or _85617_ (_35148_, _35147_, _06417_);
  or _85618_ (_35149_, _35133_, _06426_);
  and _85619_ (_35150_, _35149_, _06353_);
  and _85620_ (_35152_, _35150_, _35148_);
  and _85621_ (_35153_, _14754_, _08650_);
  or _85622_ (_35154_, _35153_, _35141_);
  and _85623_ (_35155_, _35154_, _06352_);
  or _85624_ (_35156_, _35155_, _06345_);
  or _85625_ (_35157_, _35156_, _35152_);
  and _85626_ (_35158_, _35142_, _14782_);
  or _85627_ (_35159_, _35141_, _06346_);
  or _85628_ (_35160_, _35159_, _35158_);
  and _85629_ (_35161_, _35160_, _35157_);
  and _85630_ (_35163_, _35161_, _06340_);
  and _85631_ (_35164_, _14796_, _08650_);
  or _85632_ (_35165_, _35141_, _35164_);
  and _85633_ (_35166_, _35165_, _06339_);
  or _85634_ (_35167_, _35166_, _10153_);
  or _85635_ (_35168_, _35167_, _35163_);
  or _85636_ (_35169_, _35125_, _06327_);
  and _85637_ (_35170_, _35169_, _35168_);
  or _85638_ (_35171_, _35170_, _09572_);
  and _85639_ (_35172_, _09402_, _07969_);
  or _85640_ (_35174_, _35115_, _06333_);
  or _85641_ (_35175_, _35174_, _35172_);
  and _85642_ (_35176_, _35175_, _06313_);
  and _85643_ (_35177_, _35176_, _35171_);
  and _85644_ (_35178_, _14851_, _07969_);
  or _85645_ (_35179_, _35178_, _35115_);
  and _85646_ (_35180_, _35179_, _06037_);
  or _85647_ (_35181_, _35180_, _35177_);
  and _85648_ (_35182_, _35181_, _06278_);
  or _85649_ (_35183_, _35182_, _35123_);
  and _85650_ (_35185_, _35183_, _07334_);
  or _85651_ (_35186_, _14749_, _13907_);
  and _85652_ (_35187_, _35121_, _06502_);
  and _85653_ (_35188_, _35187_, _35186_);
  or _85654_ (_35189_, _35188_, _06615_);
  or _85655_ (_35190_, _35189_, _35185_);
  and _85656_ (_35191_, _10579_, _07969_);
  or _85657_ (_35192_, _35191_, _35115_);
  or _85658_ (_35193_, _35192_, _07337_);
  and _85659_ (_35194_, _35193_, _07339_);
  and _85660_ (_35196_, _35194_, _35190_);
  or _85661_ (_35197_, _14747_, _13907_);
  and _85662_ (_35198_, _35121_, _06507_);
  and _85663_ (_35199_, _35198_, _35197_);
  or _85664_ (_35200_, _35199_, _06610_);
  or _85665_ (_35201_, _35200_, _35196_);
  and _85666_ (_35202_, _35132_, _08404_);
  or _85667_ (_35203_, _35115_, _07331_);
  or _85668_ (_35204_, _35203_, _35202_);
  and _85669_ (_35205_, _35204_, _09107_);
  and _85670_ (_35207_, _35205_, _35201_);
  or _85671_ (_35208_, _35120_, _08404_);
  and _85672_ (_35209_, _35121_, _06509_);
  and _85673_ (_35210_, _35209_, _35208_);
  or _85674_ (_35211_, _35210_, _06602_);
  or _85675_ (_35212_, _35211_, _35207_);
  and _85676_ (_35213_, _35212_, _35119_);
  or _85677_ (_35214_, _35213_, _06639_);
  or _85678_ (_35215_, _35130_, _07048_);
  and _85679_ (_35216_, _35215_, _05990_);
  and _85680_ (_35218_, _35216_, _35214_);
  and _85681_ (_35219_, _35154_, _05989_);
  or _85682_ (_35220_, _35219_, _06646_);
  or _85683_ (_35221_, _35220_, _35218_);
  or _85684_ (_35222_, _35115_, _06651_);
  or _85685_ (_35223_, _35222_, _35127_);
  and _85686_ (_35224_, _35223_, _01442_);
  and _85687_ (_35225_, _35224_, _35221_);
  or _85688_ (_35226_, _35225_, _35114_);
  and _85689_ (_44275_, _35226_, _43634_);
  and _85690_ (_35228_, _01446_, \oc8051_golden_model_1.SCON [2]);
  and _85691_ (_35229_, _13907_, \oc8051_golden_model_1.SCON [2]);
  nor _85692_ (_35230_, _10582_, _13907_);
  or _85693_ (_35231_, _35230_, _35229_);
  and _85694_ (_35232_, _07969_, \oc8051_golden_model_1.ACC [2]);
  nand _85695_ (_35233_, _35232_, _08503_);
  and _85696_ (_35234_, _35233_, _06615_);
  and _85697_ (_35235_, _35234_, _35231_);
  nor _85698_ (_35236_, _13907_, _07854_);
  or _85699_ (_35237_, _35236_, _35229_);
  or _85700_ (_35239_, _35237_, _06327_);
  or _85701_ (_35240_, _35237_, _06772_);
  and _85702_ (_35241_, _14959_, _07969_);
  or _85703_ (_35242_, _35241_, _35229_);
  or _85704_ (_35243_, _35242_, _07275_);
  or _85705_ (_35244_, _35232_, _35229_);
  and _85706_ (_35245_, _35244_, _07259_);
  and _85707_ (_35246_, _07260_, \oc8051_golden_model_1.SCON [2]);
  or _85708_ (_35247_, _35246_, _06474_);
  or _85709_ (_35248_, _35247_, _35245_);
  and _85710_ (_35250_, _35248_, _06357_);
  and _85711_ (_35251_, _35250_, _35243_);
  and _85712_ (_35252_, _13915_, \oc8051_golden_model_1.SCON [2]);
  and _85713_ (_35253_, _14955_, _08650_);
  or _85714_ (_35254_, _35253_, _35252_);
  and _85715_ (_35255_, _35254_, _06356_);
  or _85716_ (_35256_, _35255_, _06410_);
  or _85717_ (_35257_, _35256_, _35251_);
  and _85718_ (_35258_, _35257_, _35240_);
  or _85719_ (_35259_, _35258_, _06417_);
  or _85720_ (_35261_, _35244_, _06426_);
  and _85721_ (_35262_, _35261_, _06353_);
  and _85722_ (_35263_, _35262_, _35259_);
  and _85723_ (_35264_, _14953_, _08650_);
  or _85724_ (_35265_, _35264_, _35252_);
  and _85725_ (_35266_, _35265_, _06352_);
  or _85726_ (_35267_, _35266_, _06345_);
  or _85727_ (_35268_, _35267_, _35263_);
  and _85728_ (_35269_, _35253_, _14986_);
  or _85729_ (_35270_, _35252_, _06346_);
  or _85730_ (_35272_, _35270_, _35269_);
  and _85731_ (_35273_, _35272_, _06340_);
  and _85732_ (_35274_, _35273_, _35268_);
  and _85733_ (_35275_, _15000_, _08650_);
  or _85734_ (_35276_, _35275_, _35252_);
  and _85735_ (_35277_, _35276_, _06339_);
  or _85736_ (_35278_, _35277_, _10153_);
  or _85737_ (_35279_, _35278_, _35274_);
  and _85738_ (_35280_, _35279_, _35239_);
  or _85739_ (_35281_, _35280_, _09572_);
  and _85740_ (_35283_, _09356_, _07969_);
  or _85741_ (_35284_, _35229_, _06333_);
  or _85742_ (_35285_, _35284_, _35283_);
  and _85743_ (_35286_, _35285_, _06313_);
  and _85744_ (_35287_, _35286_, _35281_);
  and _85745_ (_35288_, _15056_, _07969_);
  or _85746_ (_35289_, _35288_, _35229_);
  and _85747_ (_35290_, _35289_, _06037_);
  or _85748_ (_35291_, _35290_, _06277_);
  or _85749_ (_35292_, _35291_, _35287_);
  and _85750_ (_35294_, _07969_, _09057_);
  or _85751_ (_35295_, _35294_, _35229_);
  or _85752_ (_35296_, _35295_, _06278_);
  and _85753_ (_35297_, _35296_, _35292_);
  or _85754_ (_35298_, _35297_, _06502_);
  and _85755_ (_35299_, _14948_, _07969_);
  or _85756_ (_35300_, _35229_, _07334_);
  or _85757_ (_35301_, _35300_, _35299_);
  and _85758_ (_35302_, _35301_, _07337_);
  and _85759_ (_35303_, _35302_, _35298_);
  or _85760_ (_35305_, _35303_, _35235_);
  and _85761_ (_35306_, _35305_, _07339_);
  or _85762_ (_35307_, _35229_, _08503_);
  and _85763_ (_35308_, _35295_, _06507_);
  and _85764_ (_35309_, _35308_, _35307_);
  or _85765_ (_35310_, _35309_, _35306_);
  and _85766_ (_35311_, _35310_, _07331_);
  and _85767_ (_35312_, _35244_, _06610_);
  and _85768_ (_35313_, _35312_, _35307_);
  or _85769_ (_35314_, _35313_, _06509_);
  or _85770_ (_35316_, _35314_, _35311_);
  and _85771_ (_35317_, _14945_, _07969_);
  or _85772_ (_35318_, _35229_, _09107_);
  or _85773_ (_35319_, _35318_, _35317_);
  and _85774_ (_35320_, _35319_, _09112_);
  and _85775_ (_35321_, _35320_, _35316_);
  and _85776_ (_35322_, _35231_, _06602_);
  or _85777_ (_35323_, _35322_, _06639_);
  or _85778_ (_35324_, _35323_, _35321_);
  or _85779_ (_35325_, _35242_, _07048_);
  and _85780_ (_35326_, _35325_, _05990_);
  and _85781_ (_35327_, _35326_, _35324_);
  and _85782_ (_35328_, _35265_, _05989_);
  or _85783_ (_35329_, _35328_, _06646_);
  or _85784_ (_35330_, _35329_, _35327_);
  and _85785_ (_35331_, _15129_, _07969_);
  or _85786_ (_35332_, _35229_, _06651_);
  or _85787_ (_35333_, _35332_, _35331_);
  and _85788_ (_35334_, _35333_, _01442_);
  and _85789_ (_35335_, _35334_, _35330_);
  or _85790_ (_35337_, _35335_, _35228_);
  and _85791_ (_44276_, _35337_, _43634_);
  and _85792_ (_35338_, _01446_, \oc8051_golden_model_1.SCON [3]);
  and _85793_ (_35339_, _13907_, \oc8051_golden_model_1.SCON [3]);
  nor _85794_ (_35340_, _13907_, _07680_);
  or _85795_ (_35341_, _35340_, _35339_);
  or _85796_ (_35342_, _35341_, _06327_);
  and _85797_ (_35343_, _15153_, _07969_);
  or _85798_ (_35344_, _35343_, _35339_);
  or _85799_ (_35345_, _35344_, _07275_);
  and _85800_ (_35347_, _07969_, \oc8051_golden_model_1.ACC [3]);
  or _85801_ (_35348_, _35347_, _35339_);
  and _85802_ (_35349_, _35348_, _07259_);
  and _85803_ (_35350_, _07260_, \oc8051_golden_model_1.SCON [3]);
  or _85804_ (_35351_, _35350_, _06474_);
  or _85805_ (_35352_, _35351_, _35349_);
  and _85806_ (_35353_, _35352_, _06357_);
  and _85807_ (_35354_, _35353_, _35345_);
  and _85808_ (_35355_, _13915_, \oc8051_golden_model_1.SCON [3]);
  and _85809_ (_35356_, _15150_, _08650_);
  or _85810_ (_35358_, _35356_, _35355_);
  and _85811_ (_35359_, _35358_, _06356_);
  or _85812_ (_35360_, _35359_, _06410_);
  or _85813_ (_35361_, _35360_, _35354_);
  or _85814_ (_35362_, _35341_, _06772_);
  and _85815_ (_35363_, _35362_, _35361_);
  or _85816_ (_35364_, _35363_, _06417_);
  or _85817_ (_35365_, _35348_, _06426_);
  and _85818_ (_35366_, _35365_, _06353_);
  and _85819_ (_35367_, _35366_, _35364_);
  and _85820_ (_35369_, _15148_, _08650_);
  or _85821_ (_35370_, _35369_, _35355_);
  and _85822_ (_35371_, _35370_, _06352_);
  or _85823_ (_35372_, _35371_, _06345_);
  or _85824_ (_35373_, _35372_, _35367_);
  or _85825_ (_35374_, _35355_, _15180_);
  and _85826_ (_35375_, _35374_, _35358_);
  or _85827_ (_35376_, _35375_, _06346_);
  and _85828_ (_35377_, _35376_, _06340_);
  and _85829_ (_35378_, _35377_, _35373_);
  and _85830_ (_35380_, _15197_, _08650_);
  or _85831_ (_35381_, _35380_, _35355_);
  and _85832_ (_35382_, _35381_, _06339_);
  or _85833_ (_35383_, _35382_, _10153_);
  or _85834_ (_35384_, _35383_, _35378_);
  and _85835_ (_35385_, _35384_, _35342_);
  or _85836_ (_35386_, _35385_, _09572_);
  and _85837_ (_35387_, _09310_, _07969_);
  or _85838_ (_35388_, _35339_, _06333_);
  or _85839_ (_35389_, _35388_, _35387_);
  and _85840_ (_35391_, _35389_, _06313_);
  and _85841_ (_35392_, _35391_, _35386_);
  and _85842_ (_35393_, _15251_, _07969_);
  or _85843_ (_35394_, _35393_, _35339_);
  and _85844_ (_35395_, _35394_, _06037_);
  or _85845_ (_35396_, _35395_, _06277_);
  or _85846_ (_35397_, _35396_, _35392_);
  and _85847_ (_35398_, _07969_, _09014_);
  or _85848_ (_35399_, _35398_, _35339_);
  or _85849_ (_35400_, _35399_, _06278_);
  and _85850_ (_35402_, _35400_, _35397_);
  or _85851_ (_35403_, _35402_, _06502_);
  and _85852_ (_35404_, _15266_, _07969_);
  or _85853_ (_35405_, _35339_, _07334_);
  or _85854_ (_35406_, _35405_, _35404_);
  and _85855_ (_35407_, _35406_, _07337_);
  and _85856_ (_35408_, _35407_, _35403_);
  and _85857_ (_35409_, _12619_, _07969_);
  or _85858_ (_35410_, _35409_, _35339_);
  and _85859_ (_35411_, _35410_, _06615_);
  or _85860_ (_35413_, _35411_, _35408_);
  and _85861_ (_35414_, _35413_, _07339_);
  or _85862_ (_35415_, _35339_, _08359_);
  and _85863_ (_35416_, _35399_, _06507_);
  and _85864_ (_35417_, _35416_, _35415_);
  or _85865_ (_35418_, _35417_, _35414_);
  and _85866_ (_35419_, _35418_, _07331_);
  and _85867_ (_35420_, _35348_, _06610_);
  and _85868_ (_35421_, _35420_, _35415_);
  or _85869_ (_35422_, _35421_, _06509_);
  or _85870_ (_35424_, _35422_, _35419_);
  and _85871_ (_35425_, _15263_, _07969_);
  or _85872_ (_35426_, _35339_, _09107_);
  or _85873_ (_35427_, _35426_, _35425_);
  and _85874_ (_35428_, _35427_, _09112_);
  and _85875_ (_35429_, _35428_, _35424_);
  nor _85876_ (_35430_, _10574_, _13907_);
  or _85877_ (_35431_, _35430_, _35339_);
  and _85878_ (_35432_, _35431_, _06602_);
  or _85879_ (_35433_, _35432_, _06639_);
  or _85880_ (_35435_, _35433_, _35429_);
  or _85881_ (_35436_, _35344_, _07048_);
  and _85882_ (_35437_, _35436_, _05990_);
  and _85883_ (_35438_, _35437_, _35435_);
  and _85884_ (_35439_, _35370_, _05989_);
  or _85885_ (_35440_, _35439_, _06646_);
  or _85886_ (_35441_, _35440_, _35438_);
  and _85887_ (_35442_, _15321_, _07969_);
  or _85888_ (_35443_, _35339_, _06651_);
  or _85889_ (_35444_, _35443_, _35442_);
  and _85890_ (_35446_, _35444_, _01442_);
  and _85891_ (_35447_, _35446_, _35441_);
  or _85892_ (_35448_, _35447_, _35338_);
  and _85893_ (_44277_, _35448_, _43634_);
  and _85894_ (_35449_, _01446_, \oc8051_golden_model_1.SCON [4]);
  and _85895_ (_35450_, _13907_, \oc8051_golden_model_1.SCON [4]);
  nor _85896_ (_35451_, _10589_, _13907_);
  or _85897_ (_35452_, _35451_, _35450_);
  and _85898_ (_35453_, _07969_, \oc8051_golden_model_1.ACC [4]);
  nand _85899_ (_35454_, _35453_, _08599_);
  and _85900_ (_35456_, _35454_, _06615_);
  and _85901_ (_35457_, _35456_, _35452_);
  nor _85902_ (_35458_, _08596_, _13907_);
  or _85903_ (_35459_, _35458_, _35450_);
  or _85904_ (_35460_, _35459_, _06327_);
  and _85905_ (_35461_, _13915_, \oc8051_golden_model_1.SCON [4]);
  and _85906_ (_35462_, _15348_, _08650_);
  or _85907_ (_35463_, _35462_, _35461_);
  and _85908_ (_35464_, _35463_, _06352_);
  and _85909_ (_35465_, _15367_, _07969_);
  or _85910_ (_35467_, _35465_, _35450_);
  or _85911_ (_35468_, _35467_, _07275_);
  or _85912_ (_35469_, _35453_, _35450_);
  and _85913_ (_35470_, _35469_, _07259_);
  and _85914_ (_35471_, _07260_, \oc8051_golden_model_1.SCON [4]);
  or _85915_ (_35472_, _35471_, _06474_);
  or _85916_ (_35473_, _35472_, _35470_);
  and _85917_ (_35474_, _35473_, _06357_);
  and _85918_ (_35475_, _35474_, _35468_);
  and _85919_ (_35476_, _15353_, _08650_);
  or _85920_ (_35478_, _35476_, _35461_);
  and _85921_ (_35479_, _35478_, _06356_);
  or _85922_ (_35480_, _35479_, _06410_);
  or _85923_ (_35481_, _35480_, _35475_);
  or _85924_ (_35482_, _35459_, _06772_);
  and _85925_ (_35483_, _35482_, _35481_);
  or _85926_ (_35484_, _35483_, _06417_);
  or _85927_ (_35485_, _35469_, _06426_);
  and _85928_ (_35486_, _35485_, _06353_);
  and _85929_ (_35487_, _35486_, _35484_);
  or _85930_ (_35489_, _35487_, _35464_);
  and _85931_ (_35490_, _35489_, _06346_);
  and _85932_ (_35491_, _15385_, _08650_);
  or _85933_ (_35492_, _35491_, _35461_);
  and _85934_ (_35493_, _35492_, _06345_);
  or _85935_ (_35494_, _35493_, _35490_);
  and _85936_ (_35495_, _35494_, _06340_);
  and _85937_ (_35496_, _15350_, _08650_);
  or _85938_ (_35497_, _35496_, _35461_);
  and _85939_ (_35498_, _35497_, _06339_);
  or _85940_ (_35500_, _35498_, _10153_);
  or _85941_ (_35501_, _35500_, _35495_);
  and _85942_ (_35502_, _35501_, _35460_);
  or _85943_ (_35503_, _35502_, _09572_);
  and _85944_ (_35504_, _09264_, _07969_);
  or _85945_ (_35505_, _35450_, _06333_);
  or _85946_ (_35506_, _35505_, _35504_);
  and _85947_ (_35507_, _35506_, _06313_);
  and _85948_ (_35508_, _35507_, _35503_);
  and _85949_ (_35509_, _15452_, _07969_);
  or _85950_ (_35511_, _35509_, _35450_);
  and _85951_ (_35512_, _35511_, _06037_);
  or _85952_ (_35513_, _35512_, _06277_);
  or _85953_ (_35514_, _35513_, _35508_);
  and _85954_ (_35515_, _08995_, _07969_);
  or _85955_ (_35516_, _35515_, _35450_);
  or _85956_ (_35517_, _35516_, _06278_);
  and _85957_ (_35518_, _35517_, _35514_);
  or _85958_ (_35519_, _35518_, _06502_);
  and _85959_ (_35520_, _15345_, _07969_);
  or _85960_ (_35522_, _35450_, _07334_);
  or _85961_ (_35523_, _35522_, _35520_);
  and _85962_ (_35524_, _35523_, _07337_);
  and _85963_ (_35525_, _35524_, _35519_);
  or _85964_ (_35526_, _35525_, _35457_);
  and _85965_ (_35527_, _35526_, _07339_);
  or _85966_ (_35528_, _35450_, _08599_);
  and _85967_ (_35529_, _35516_, _06507_);
  and _85968_ (_35530_, _35529_, _35528_);
  or _85969_ (_35531_, _35530_, _35527_);
  and _85970_ (_35533_, _35531_, _07331_);
  and _85971_ (_35534_, _35469_, _06610_);
  and _85972_ (_35535_, _35534_, _35528_);
  or _85973_ (_35536_, _35535_, _06509_);
  or _85974_ (_35537_, _35536_, _35533_);
  and _85975_ (_35538_, _15342_, _07969_);
  or _85976_ (_35539_, _35450_, _09107_);
  or _85977_ (_35540_, _35539_, _35538_);
  and _85978_ (_35541_, _35540_, _09112_);
  and _85979_ (_35542_, _35541_, _35537_);
  and _85980_ (_35544_, _35452_, _06602_);
  or _85981_ (_35545_, _35544_, _06639_);
  or _85982_ (_35546_, _35545_, _35542_);
  or _85983_ (_35547_, _35467_, _07048_);
  and _85984_ (_35548_, _35547_, _05990_);
  and _85985_ (_35549_, _35548_, _35546_);
  and _85986_ (_35550_, _35463_, _05989_);
  or _85987_ (_35551_, _35550_, _06646_);
  or _85988_ (_35552_, _35551_, _35549_);
  and _85989_ (_35553_, _15524_, _07969_);
  or _85990_ (_35555_, _35450_, _06651_);
  or _85991_ (_35556_, _35555_, _35553_);
  and _85992_ (_35557_, _35556_, _01442_);
  and _85993_ (_35558_, _35557_, _35552_);
  or _85994_ (_35559_, _35558_, _35449_);
  and _85995_ (_44278_, _35559_, _43634_);
  and _85996_ (_35560_, _01446_, \oc8051_golden_model_1.SCON [5]);
  and _85997_ (_35561_, _13907_, \oc8051_golden_model_1.SCON [5]);
  nor _85998_ (_35562_, _10570_, _13907_);
  or _85999_ (_35563_, _35562_, _35561_);
  and _86000_ (_35565_, _07969_, \oc8051_golden_model_1.ACC [5]);
  nand _86001_ (_35566_, _35565_, _08308_);
  and _86002_ (_35567_, _35566_, _06615_);
  and _86003_ (_35568_, _35567_, _35563_);
  and _86004_ (_35569_, _15550_, _07969_);
  or _86005_ (_35570_, _35569_, _35561_);
  or _86006_ (_35571_, _35570_, _07275_);
  or _86007_ (_35572_, _35565_, _35561_);
  and _86008_ (_35573_, _35572_, _07259_);
  and _86009_ (_35574_, _07260_, \oc8051_golden_model_1.SCON [5]);
  or _86010_ (_35576_, _35574_, _06474_);
  or _86011_ (_35577_, _35576_, _35573_);
  and _86012_ (_35578_, _35577_, _06357_);
  and _86013_ (_35579_, _35578_, _35571_);
  and _86014_ (_35580_, _13915_, \oc8051_golden_model_1.SCON [5]);
  and _86015_ (_35581_, _15566_, _08650_);
  or _86016_ (_35582_, _35581_, _35580_);
  and _86017_ (_35583_, _35582_, _06356_);
  or _86018_ (_35584_, _35583_, _06410_);
  or _86019_ (_35585_, _35584_, _35579_);
  nor _86020_ (_35587_, _08305_, _13907_);
  or _86021_ (_35588_, _35587_, _35561_);
  or _86022_ (_35589_, _35588_, _06772_);
  and _86023_ (_35590_, _35589_, _35585_);
  or _86024_ (_35591_, _35590_, _06417_);
  or _86025_ (_35592_, _35572_, _06426_);
  and _86026_ (_35593_, _35592_, _06353_);
  and _86027_ (_35594_, _35593_, _35591_);
  and _86028_ (_35595_, _15544_, _08650_);
  or _86029_ (_35596_, _35595_, _35580_);
  and _86030_ (_35598_, _35596_, _06352_);
  or _86031_ (_35599_, _35598_, _06345_);
  or _86032_ (_35600_, _35599_, _35594_);
  or _86033_ (_35601_, _35580_, _15581_);
  and _86034_ (_35602_, _35601_, _35582_);
  or _86035_ (_35603_, _35602_, _06346_);
  and _86036_ (_35604_, _35603_, _06340_);
  and _86037_ (_35605_, _35604_, _35600_);
  and _86038_ (_35606_, _15546_, _08650_);
  or _86039_ (_35607_, _35606_, _35580_);
  and _86040_ (_35609_, _35607_, _06339_);
  or _86041_ (_35610_, _35609_, _10153_);
  or _86042_ (_35611_, _35610_, _35605_);
  or _86043_ (_35612_, _35588_, _06327_);
  and _86044_ (_35613_, _35612_, _35611_);
  or _86045_ (_35614_, _35613_, _09572_);
  and _86046_ (_35615_, _09218_, _07969_);
  or _86047_ (_35616_, _35561_, _06333_);
  or _86048_ (_35617_, _35616_, _35615_);
  and _86049_ (_35618_, _35617_, _06313_);
  and _86050_ (_35620_, _35618_, _35614_);
  and _86051_ (_35621_, _15649_, _07969_);
  or _86052_ (_35622_, _35621_, _35561_);
  and _86053_ (_35623_, _35622_, _06037_);
  or _86054_ (_35624_, _35623_, _06277_);
  or _86055_ (_35625_, _35624_, _35620_);
  and _86056_ (_35626_, _08954_, _07969_);
  or _86057_ (_35627_, _35626_, _35561_);
  or _86058_ (_35628_, _35627_, _06278_);
  and _86059_ (_35629_, _35628_, _35625_);
  or _86060_ (_35631_, _35629_, _06502_);
  and _86061_ (_35632_, _15664_, _07969_);
  or _86062_ (_35633_, _35561_, _07334_);
  or _86063_ (_35634_, _35633_, _35632_);
  and _86064_ (_35635_, _35634_, _07337_);
  and _86065_ (_35636_, _35635_, _35631_);
  or _86066_ (_35637_, _35636_, _35568_);
  and _86067_ (_35638_, _35637_, _07339_);
  or _86068_ (_35639_, _35561_, _08308_);
  and _86069_ (_35640_, _35627_, _06507_);
  and _86070_ (_35642_, _35640_, _35639_);
  or _86071_ (_35643_, _35642_, _35638_);
  and _86072_ (_35644_, _35643_, _07331_);
  and _86073_ (_35645_, _35572_, _06610_);
  and _86074_ (_35646_, _35645_, _35639_);
  or _86075_ (_35647_, _35646_, _06509_);
  or _86076_ (_35648_, _35647_, _35644_);
  and _86077_ (_35649_, _15663_, _07969_);
  or _86078_ (_35650_, _35561_, _09107_);
  or _86079_ (_35651_, _35650_, _35649_);
  and _86080_ (_35653_, _35651_, _09112_);
  and _86081_ (_35654_, _35653_, _35648_);
  and _86082_ (_35655_, _35563_, _06602_);
  or _86083_ (_35656_, _35655_, _06639_);
  or _86084_ (_35657_, _35656_, _35654_);
  or _86085_ (_35658_, _35570_, _07048_);
  and _86086_ (_35659_, _35658_, _05990_);
  and _86087_ (_35660_, _35659_, _35657_);
  and _86088_ (_35661_, _35596_, _05989_);
  or _86089_ (_35662_, _35661_, _06646_);
  or _86090_ (_35664_, _35662_, _35660_);
  and _86091_ (_35665_, _15721_, _07969_);
  or _86092_ (_35666_, _35561_, _06651_);
  or _86093_ (_35667_, _35666_, _35665_);
  and _86094_ (_35668_, _35667_, _01442_);
  and _86095_ (_35669_, _35668_, _35664_);
  or _86096_ (_35670_, _35669_, _35560_);
  and _86097_ (_44279_, _35670_, _43634_);
  and _86098_ (_35671_, _01446_, \oc8051_golden_model_1.SCON [6]);
  and _86099_ (_35672_, _13907_, \oc8051_golden_model_1.SCON [6]);
  and _86100_ (_35674_, _15759_, _07969_);
  or _86101_ (_35675_, _35674_, _35672_);
  or _86102_ (_35676_, _35675_, _07275_);
  and _86103_ (_35677_, _07969_, \oc8051_golden_model_1.ACC [6]);
  or _86104_ (_35678_, _35677_, _35672_);
  and _86105_ (_35679_, _35678_, _07259_);
  and _86106_ (_35680_, _07260_, \oc8051_golden_model_1.SCON [6]);
  or _86107_ (_35681_, _35680_, _06474_);
  or _86108_ (_35682_, _35681_, _35679_);
  and _86109_ (_35683_, _35682_, _06357_);
  and _86110_ (_35685_, _35683_, _35676_);
  and _86111_ (_35686_, _13915_, \oc8051_golden_model_1.SCON [6]);
  and _86112_ (_35687_, _15763_, _08650_);
  or _86113_ (_35688_, _35687_, _35686_);
  and _86114_ (_35689_, _35688_, _06356_);
  or _86115_ (_35690_, _35689_, _06410_);
  or _86116_ (_35691_, _35690_, _35685_);
  nor _86117_ (_35692_, _08209_, _13907_);
  or _86118_ (_35693_, _35692_, _35672_);
  or _86119_ (_35694_, _35693_, _06772_);
  and _86120_ (_35696_, _35694_, _35691_);
  or _86121_ (_35697_, _35696_, _06417_);
  or _86122_ (_35698_, _35678_, _06426_);
  and _86123_ (_35699_, _35698_, _06353_);
  and _86124_ (_35700_, _35699_, _35697_);
  and _86125_ (_35701_, _15743_, _08650_);
  or _86126_ (_35702_, _35701_, _35686_);
  and _86127_ (_35703_, _35702_, _06352_);
  or _86128_ (_35704_, _35703_, _06345_);
  or _86129_ (_35705_, _35704_, _35700_);
  or _86130_ (_35707_, _35686_, _15778_);
  and _86131_ (_35708_, _35707_, _35688_);
  or _86132_ (_35709_, _35708_, _06346_);
  and _86133_ (_35710_, _35709_, _06340_);
  and _86134_ (_35711_, _35710_, _35705_);
  and _86135_ (_35712_, _15745_, _08650_);
  or _86136_ (_35713_, _35712_, _35686_);
  and _86137_ (_35714_, _35713_, _06339_);
  or _86138_ (_35715_, _35714_, _10153_);
  or _86139_ (_35716_, _35715_, _35711_);
  or _86140_ (_35718_, _35693_, _06327_);
  and _86141_ (_35719_, _35718_, _35716_);
  or _86142_ (_35720_, _35719_, _09572_);
  and _86143_ (_35721_, _09172_, _07969_);
  or _86144_ (_35722_, _35672_, _06333_);
  or _86145_ (_35723_, _35722_, _35721_);
  and _86146_ (_35724_, _35723_, _06313_);
  and _86147_ (_35725_, _35724_, _35720_);
  and _86148_ (_35726_, _15846_, _07969_);
  or _86149_ (_35727_, _35726_, _35672_);
  and _86150_ (_35729_, _35727_, _06037_);
  or _86151_ (_35730_, _35729_, _06277_);
  or _86152_ (_35731_, _35730_, _35725_);
  and _86153_ (_35732_, _15853_, _07969_);
  or _86154_ (_35733_, _35732_, _35672_);
  or _86155_ (_35734_, _35733_, _06278_);
  and _86156_ (_35735_, _35734_, _35731_);
  or _86157_ (_35736_, _35735_, _06502_);
  and _86158_ (_35737_, _15862_, _07969_);
  or _86159_ (_35738_, _35672_, _07334_);
  or _86160_ (_35740_, _35738_, _35737_);
  and _86161_ (_35741_, _35740_, _07337_);
  and _86162_ (_35742_, _35741_, _35736_);
  and _86163_ (_35743_, _10596_, _07969_);
  or _86164_ (_35744_, _35743_, _35672_);
  and _86165_ (_35745_, _35744_, _06615_);
  or _86166_ (_35746_, _35745_, _35742_);
  and _86167_ (_35747_, _35746_, _07339_);
  or _86168_ (_35748_, _35672_, _08212_);
  and _86169_ (_35749_, _35733_, _06507_);
  and _86170_ (_35751_, _35749_, _35748_);
  or _86171_ (_35752_, _35751_, _35747_);
  and _86172_ (_35753_, _35752_, _07331_);
  and _86173_ (_35754_, _35678_, _06610_);
  and _86174_ (_35755_, _35754_, _35748_);
  or _86175_ (_35756_, _35755_, _06509_);
  or _86176_ (_35757_, _35756_, _35753_);
  and _86177_ (_35758_, _15859_, _07969_);
  or _86178_ (_35759_, _35672_, _09107_);
  or _86179_ (_35760_, _35759_, _35758_);
  and _86180_ (_35762_, _35760_, _09112_);
  and _86181_ (_35763_, _35762_, _35757_);
  nor _86182_ (_35764_, _10595_, _13907_);
  or _86183_ (_35765_, _35764_, _35672_);
  and _86184_ (_35766_, _35765_, _06602_);
  or _86185_ (_35767_, _35766_, _06639_);
  or _86186_ (_35768_, _35767_, _35763_);
  or _86187_ (_35769_, _35675_, _07048_);
  and _86188_ (_35770_, _35769_, _05990_);
  and _86189_ (_35771_, _35770_, _35768_);
  and _86190_ (_35773_, _35702_, _05989_);
  or _86191_ (_35774_, _35773_, _06646_);
  or _86192_ (_35775_, _35774_, _35771_);
  and _86193_ (_35776_, _15921_, _07969_);
  or _86194_ (_35777_, _35672_, _06651_);
  or _86195_ (_35778_, _35777_, _35776_);
  and _86196_ (_35779_, _35778_, _01442_);
  and _86197_ (_35780_, _35779_, _35775_);
  or _86198_ (_35781_, _35780_, _35671_);
  and _86199_ (_44280_, _35781_, _43634_);
  nor _86200_ (_35783_, _01442_, _06342_);
  nor _86201_ (_35784_, _08004_, _06342_);
  nor _86202_ (_35785_, _08453_, _14023_);
  or _86203_ (_35786_, _35785_, _35784_);
  or _86204_ (_35787_, _35786_, _07275_);
  and _86205_ (_35788_, _08004_, \oc8051_golden_model_1.ACC [0]);
  or _86206_ (_35789_, _35788_, _35784_);
  and _86207_ (_35790_, _35789_, _07259_);
  nor _86208_ (_35791_, _07259_, _06342_);
  or _86209_ (_35792_, _35791_, _06474_);
  or _86210_ (_35794_, _35792_, _35790_);
  and _86211_ (_35795_, _35794_, _06772_);
  nand _86212_ (_35796_, _35795_, _35787_);
  nand _86213_ (_35797_, _35796_, _06875_);
  or _86214_ (_35798_, _35789_, _06426_);
  and _86215_ (_35799_, _35798_, _07394_);
  and _86216_ (_35800_, _35799_, _35797_);
  nand _86217_ (_35801_, _06327_, _07301_);
  or _86218_ (_35802_, _35801_, _35800_);
  and _86219_ (_35803_, _08004_, _07250_);
  or _86220_ (_35805_, _35784_, _06327_);
  or _86221_ (_35806_, _35805_, _35803_);
  and _86222_ (_35807_, _35806_, _35802_);
  or _86223_ (_35808_, _35807_, _09572_);
  and _86224_ (_35809_, _09447_, _08004_);
  or _86225_ (_35810_, _35784_, _06333_);
  or _86226_ (_35811_, _35810_, _35809_);
  and _86227_ (_35812_, _35811_, _35808_);
  or _86228_ (_35813_, _35812_, _06037_);
  and _86229_ (_35814_, _14666_, _08004_);
  or _86230_ (_35816_, _35784_, _06313_);
  or _86231_ (_35817_, _35816_, _35814_);
  and _86232_ (_35818_, _35817_, _06278_);
  and _86233_ (_35819_, _35818_, _35813_);
  and _86234_ (_35820_, _08004_, _09008_);
  or _86235_ (_35821_, _35820_, _35784_);
  and _86236_ (_35822_, _35821_, _06277_);
  or _86237_ (_35823_, _35822_, _06502_);
  or _86238_ (_35824_, _35823_, _35819_);
  and _86239_ (_35825_, _14566_, _08004_);
  or _86240_ (_35827_, _35784_, _07334_);
  or _86241_ (_35828_, _35827_, _35825_);
  and _86242_ (_35829_, _35828_, _07337_);
  and _86243_ (_35830_, _35829_, _35824_);
  nor _86244_ (_35831_, _12622_, _14023_);
  or _86245_ (_35832_, _35831_, _35784_);
  and _86246_ (_35833_, _35788_, _08453_);
  nor _86247_ (_35834_, _35833_, _07337_);
  and _86248_ (_35835_, _35834_, _35832_);
  or _86249_ (_35836_, _35835_, _35830_);
  and _86250_ (_35838_, _35836_, _07339_);
  nand _86251_ (_35839_, _35821_, _06507_);
  nor _86252_ (_35840_, _35839_, _35785_);
  or _86253_ (_35841_, _35840_, _06610_);
  or _86254_ (_35842_, _35841_, _35838_);
  or _86255_ (_35843_, _35833_, _35784_);
  or _86256_ (_35844_, _35843_, _07331_);
  and _86257_ (_35845_, _35844_, _35842_);
  or _86258_ (_35846_, _35845_, _06509_);
  and _86259_ (_35847_, _14563_, _08004_);
  or _86260_ (_35849_, _35784_, _09107_);
  or _86261_ (_35850_, _35849_, _35847_);
  and _86262_ (_35851_, _35850_, _09112_);
  and _86263_ (_35852_, _35851_, _35846_);
  and _86264_ (_35853_, _35832_, _06602_);
  or _86265_ (_35854_, _35853_, _19642_);
  or _86266_ (_35855_, _35854_, _35852_);
  or _86267_ (_35856_, _35786_, _19641_);
  and _86268_ (_35857_, _35856_, _01442_);
  and _86269_ (_35858_, _35857_, _35855_);
  or _86270_ (_35860_, _35858_, _35783_);
  and _86271_ (_44282_, _35860_, _43634_);
  nand _86272_ (_35861_, _06621_, \oc8051_golden_model_1.SP [1]);
  or _86273_ (_35862_, _08004_, \oc8051_golden_model_1.SP [1]);
  and _86274_ (_35863_, _14744_, _08004_);
  not _86275_ (_35864_, _35863_);
  and _86276_ (_35865_, _35864_, _35862_);
  or _86277_ (_35866_, _35865_, _07275_);
  nand _86278_ (_35867_, _06816_, \oc8051_golden_model_1.SP [1]);
  nor _86279_ (_35868_, _08004_, _07185_);
  and _86280_ (_35870_, _08004_, \oc8051_golden_model_1.ACC [1]);
  or _86281_ (_35871_, _35870_, _35868_);
  and _86282_ (_35872_, _35871_, _07259_);
  nor _86283_ (_35873_, _07259_, _07185_);
  or _86284_ (_35874_, _35873_, _06816_);
  or _86285_ (_35875_, _35874_, _35872_);
  and _86286_ (_35876_, _35875_, _35867_);
  or _86287_ (_35877_, _35876_, _06474_);
  and _86288_ (_35878_, _35877_, _06052_);
  and _86289_ (_35879_, _35878_, _35866_);
  nor _86290_ (_35881_, _06052_, \oc8051_golden_model_1.SP [1]);
  or _86291_ (_35882_, _35881_, _06410_);
  or _86292_ (_35883_, _35882_, _35879_);
  nand _86293_ (_35884_, _07392_, _06410_);
  and _86294_ (_35885_, _35884_, _35883_);
  or _86295_ (_35886_, _35885_, _06417_);
  or _86296_ (_35887_, _35871_, _06426_);
  and _86297_ (_35888_, _35887_, _07394_);
  and _86298_ (_35889_, _35888_, _35886_);
  or _86299_ (_35890_, _14062_, _07393_);
  or _86300_ (_35892_, _35890_, _35889_);
  nand _86301_ (_35893_, _14062_, \oc8051_golden_model_1.SP [1]);
  and _86302_ (_35894_, _35893_, _06327_);
  and _86303_ (_35895_, _35894_, _35892_);
  nand _86304_ (_35896_, _08004_, _07448_);
  and _86305_ (_35897_, _35862_, _10153_);
  and _86306_ (_35898_, _35897_, _35896_);
  or _86307_ (_35899_, _35898_, _09572_);
  or _86308_ (_35900_, _35899_, _35895_);
  and _86309_ (_35901_, _09402_, _08004_);
  or _86310_ (_35903_, _35868_, _06333_);
  or _86311_ (_35904_, _35903_, _35901_);
  and _86312_ (_35905_, _35904_, _06313_);
  and _86313_ (_35906_, _35905_, _35900_);
  and _86314_ (_35907_, _14851_, _08004_);
  or _86315_ (_35908_, _35907_, _35868_);
  and _86316_ (_35909_, _35908_, _06037_);
  or _86317_ (_35910_, _35909_, _35906_);
  and _86318_ (_35911_, _35910_, _06278_);
  nand _86319_ (_35912_, _08004_, _07160_);
  and _86320_ (_35914_, _35862_, _06277_);
  and _86321_ (_35915_, _35914_, _35912_);
  or _86322_ (_35916_, _35915_, _06275_);
  or _86323_ (_35917_, _35916_, _35911_);
  nor _86324_ (_35918_, _06009_, _07185_);
  nor _86325_ (_35919_, _35918_, _06502_);
  and _86326_ (_35920_, _35919_, _35917_);
  or _86327_ (_35921_, _14749_, _14023_);
  and _86328_ (_35922_, _35862_, _06502_);
  and _86329_ (_35923_, _35922_, _35921_);
  or _86330_ (_35925_, _35923_, _06615_);
  or _86331_ (_35926_, _35925_, _35920_);
  and _86332_ (_35927_, _10579_, _08004_);
  or _86333_ (_35928_, _35927_, _35868_);
  or _86334_ (_35929_, _35928_, _07337_);
  and _86335_ (_35930_, _35929_, _07339_);
  and _86336_ (_35931_, _35930_, _35926_);
  or _86337_ (_35932_, _14747_, _14023_);
  and _86338_ (_35933_, _35862_, _06507_);
  and _86339_ (_35934_, _35933_, _35932_);
  or _86340_ (_35936_, _35934_, _06610_);
  or _86341_ (_35937_, _35936_, _35931_);
  and _86342_ (_35938_, _35870_, _08404_);
  or _86343_ (_35939_, _35938_, _35868_);
  or _86344_ (_35940_, _35939_, _07331_);
  and _86345_ (_35941_, _35940_, _35937_);
  or _86346_ (_35942_, _35941_, _07330_);
  nor _86347_ (_35943_, _06018_, _07185_);
  nor _86348_ (_35944_, _35943_, _06509_);
  and _86349_ (_35945_, _35944_, _35942_);
  or _86350_ (_35947_, _35912_, _08404_);
  and _86351_ (_35948_, _35862_, _06509_);
  and _86352_ (_35949_, _35948_, _35947_);
  or _86353_ (_35950_, _35949_, _35945_);
  and _86354_ (_35951_, _35950_, _09112_);
  nor _86355_ (_35952_, _10578_, _14023_);
  or _86356_ (_35953_, _35952_, _35868_);
  and _86357_ (_35954_, _35953_, _06602_);
  or _86358_ (_35955_, _35954_, _06621_);
  or _86359_ (_35956_, _35955_, _35951_);
  nand _86360_ (_35958_, _35956_, _35861_);
  nor _86361_ (_35959_, _06361_, _07350_);
  nand _86362_ (_35960_, _35959_, _35958_);
  or _86363_ (_35961_, _35959_, _07185_);
  and _86364_ (_35962_, _35961_, _07048_);
  and _86365_ (_35963_, _35962_, _35960_);
  and _86366_ (_35964_, _35865_, _06639_);
  or _86367_ (_35965_, _35964_, _07783_);
  or _86368_ (_35966_, _35965_, _35963_);
  or _86369_ (_35967_, _07367_, _07185_);
  and _86370_ (_35969_, _35967_, _06651_);
  and _86371_ (_35970_, _35969_, _35966_);
  or _86372_ (_35971_, _35868_, _35863_);
  and _86373_ (_35972_, _35971_, _06646_);
  or _86374_ (_35973_, _35972_, _01446_);
  or _86375_ (_35974_, _35973_, _35970_);
  or _86376_ (_35975_, _01442_, \oc8051_golden_model_1.SP [1]);
  and _86377_ (_35976_, _35975_, _43634_);
  and _86378_ (_44283_, _35976_, _35974_);
  nor _86379_ (_35977_, _01442_, _06771_);
  or _86380_ (_35979_, _09521_, _06009_);
  nor _86381_ (_35980_, _14023_, _07854_);
  nor _86382_ (_35981_, _08004_, _06771_);
  or _86383_ (_35982_, _35981_, _06327_);
  or _86384_ (_35983_, _35982_, _35980_);
  and _86385_ (_35984_, _14959_, _08004_);
  or _86386_ (_35985_, _35984_, _35981_);
  or _86387_ (_35986_, _35985_, _07275_);
  and _86388_ (_35987_, _08004_, \oc8051_golden_model_1.ACC [2]);
  or _86389_ (_35988_, _35987_, _35981_);
  or _86390_ (_35990_, _35988_, _07260_);
  or _86391_ (_35991_, _07259_, \oc8051_golden_model_1.SP [2]);
  and _86392_ (_35992_, _35991_, _07564_);
  and _86393_ (_35993_, _35992_, _35990_);
  and _86394_ (_35994_, _09521_, _06816_);
  or _86395_ (_35995_, _35994_, _06474_);
  or _86396_ (_35996_, _35995_, _35993_);
  and _86397_ (_35997_, _35996_, _06052_);
  and _86398_ (_35998_, _35997_, _35986_);
  nor _86399_ (_35999_, _16265_, _06052_);
  or _86400_ (_36001_, _35999_, _06410_);
  or _86401_ (_36002_, _36001_, _35998_);
  nand _86402_ (_36003_, _08716_, _06410_);
  and _86403_ (_36004_, _36003_, _36002_);
  or _86404_ (_36005_, _36004_, _06417_);
  or _86405_ (_36006_, _35988_, _06426_);
  and _86406_ (_36007_, _36006_, _07394_);
  and _86407_ (_36008_, _36007_, _36005_);
  or _86408_ (_36009_, _07808_, _07596_);
  or _86409_ (_36010_, _36009_, _36008_);
  nor _86410_ (_36012_, _09521_, _06049_);
  nor _86411_ (_36013_, _36012_, _06039_);
  and _86412_ (_36014_, _36013_, _36010_);
  nand _86413_ (_36015_, _09521_, _06039_);
  nand _86414_ (_36016_, _36015_, _06327_);
  or _86415_ (_36017_, _36016_, _36014_);
  and _86416_ (_36018_, _36017_, _35983_);
  or _86417_ (_36019_, _36018_, _09572_);
  and _86418_ (_36020_, _09356_, _08004_);
  or _86419_ (_36021_, _35981_, _06333_);
  or _86420_ (_36023_, _36021_, _36020_);
  and _86421_ (_36024_, _36023_, _06313_);
  and _86422_ (_36025_, _36024_, _36019_);
  and _86423_ (_36026_, _15056_, _08004_);
  or _86424_ (_36027_, _36026_, _35981_);
  and _86425_ (_36028_, _36027_, _06037_);
  or _86426_ (_36029_, _36028_, _06277_);
  or _86427_ (_36030_, _36029_, _36025_);
  and _86428_ (_36031_, _08004_, _09057_);
  or _86429_ (_36032_, _36031_, _35981_);
  or _86430_ (_36034_, _36032_, _06278_);
  and _86431_ (_36035_, _36034_, _36030_);
  or _86432_ (_36036_, _36035_, _06275_);
  and _86433_ (_36037_, _36036_, _35979_);
  or _86434_ (_36038_, _36037_, _06502_);
  and _86435_ (_36039_, _14948_, _08004_);
  or _86436_ (_36040_, _35981_, _07334_);
  or _86437_ (_36041_, _36040_, _36039_);
  and _86438_ (_36042_, _36041_, _07337_);
  and _86439_ (_36043_, _36042_, _36038_);
  and _86440_ (_36045_, _10583_, _08004_);
  or _86441_ (_36046_, _36045_, _35981_);
  and _86442_ (_36047_, _36046_, _06615_);
  or _86443_ (_36048_, _36047_, _36043_);
  and _86444_ (_36049_, _36048_, _07339_);
  or _86445_ (_36050_, _35981_, _08503_);
  and _86446_ (_36051_, _36032_, _06507_);
  and _86447_ (_36052_, _36051_, _36050_);
  or _86448_ (_36053_, _36052_, _36049_);
  and _86449_ (_36054_, _36053_, _12805_);
  and _86450_ (_36056_, _35988_, _06610_);
  and _86451_ (_36057_, _36056_, _36050_);
  nor _86452_ (_36058_, _16265_, _06018_);
  or _86453_ (_36059_, _36058_, _06509_);
  or _86454_ (_36060_, _36059_, _36057_);
  or _86455_ (_36061_, _36060_, _36054_);
  and _86456_ (_36062_, _14945_, _08004_);
  or _86457_ (_36063_, _36062_, _35981_);
  or _86458_ (_36064_, _36063_, _09107_);
  and _86459_ (_36065_, _36064_, _36061_);
  or _86460_ (_36067_, _36065_, _06602_);
  nor _86461_ (_36068_, _10582_, _14023_);
  or _86462_ (_36069_, _36068_, _35981_);
  or _86463_ (_36070_, _36069_, _09112_);
  and _86464_ (_36071_, _36070_, _14116_);
  and _86465_ (_36072_, _36071_, _36067_);
  and _86466_ (_36073_, _16265_, _06621_);
  or _86467_ (_36074_, _36073_, _07350_);
  or _86468_ (_36075_, _36074_, _36072_);
  nor _86469_ (_36076_, _09521_, _06016_);
  nor _86470_ (_36078_, _36076_, _06361_);
  and _86471_ (_36079_, _36078_, _36075_);
  and _86472_ (_36080_, _16265_, _06361_);
  or _86473_ (_36081_, _36080_, _06639_);
  or _86474_ (_36082_, _36081_, _36079_);
  or _86475_ (_36083_, _35985_, _07048_);
  and _86476_ (_36084_, _36083_, _07367_);
  and _86477_ (_36085_, _36084_, _36082_);
  nor _86478_ (_36086_, _16265_, _07367_);
  or _86479_ (_36087_, _36086_, _06646_);
  or _86480_ (_36089_, _36087_, _36085_);
  and _86481_ (_36090_, _15129_, _08004_);
  or _86482_ (_36091_, _35981_, _06651_);
  or _86483_ (_36092_, _36091_, _36090_);
  and _86484_ (_36093_, _36092_, _01442_);
  and _86485_ (_36094_, _36093_, _36089_);
  or _86486_ (_36095_, _36094_, _35977_);
  and _86487_ (_44284_, _36095_, _43634_);
  nor _86488_ (_36096_, _01442_, _06409_);
  or _86489_ (_36097_, _09518_, _07367_);
  or _86490_ (_36099_, _09518_, _06016_);
  nor _86491_ (_36100_, _08004_, _06409_);
  nor _86492_ (_36101_, _10574_, _14023_);
  or _86493_ (_36102_, _36101_, _36100_);
  and _86494_ (_36103_, _08004_, \oc8051_golden_model_1.ACC [3]);
  nand _86495_ (_36104_, _36103_, _08359_);
  and _86496_ (_36105_, _36104_, _06615_);
  and _86497_ (_36106_, _36105_, _36102_);
  or _86498_ (_36107_, _09518_, _06009_);
  nor _86499_ (_36108_, _14023_, _07680_);
  or _86500_ (_36110_, _36100_, _14025_);
  or _86501_ (_36111_, _36110_, _36108_);
  and _86502_ (_36112_, _36111_, _14022_);
  and _86503_ (_36113_, _15153_, _08004_);
  or _86504_ (_36114_, _36113_, _36100_);
  or _86505_ (_36115_, _36114_, _07275_);
  or _86506_ (_36116_, _36103_, _36100_);
  or _86507_ (_36117_, _36116_, _07260_);
  or _86508_ (_36118_, _07259_, \oc8051_golden_model_1.SP [3]);
  and _86509_ (_36119_, _36118_, _07564_);
  and _86510_ (_36120_, _36119_, _36117_);
  and _86511_ (_36121_, _09518_, _06816_);
  or _86512_ (_36122_, _36121_, _06474_);
  or _86513_ (_36123_, _36122_, _36120_);
  and _86514_ (_36124_, _36123_, _06052_);
  and _86515_ (_36125_, _36124_, _36115_);
  nor _86516_ (_36126_, _16085_, _06052_);
  or _86517_ (_36127_, _36126_, _06410_);
  or _86518_ (_36128_, _36127_, _36125_);
  nand _86519_ (_36129_, _08701_, _06410_);
  and _86520_ (_36131_, _36129_, _36128_);
  or _86521_ (_36132_, _36131_, _06417_);
  or _86522_ (_36133_, _36116_, _06426_);
  and _86523_ (_36134_, _36133_, _07394_);
  and _86524_ (_36135_, _36134_, _36132_);
  or _86525_ (_36136_, _07731_, _14062_);
  or _86526_ (_36137_, _36136_, _36135_);
  nand _86527_ (_36138_, _16085_, _14062_);
  and _86528_ (_36139_, _36138_, _06327_);
  and _86529_ (_36140_, _36139_, _36137_);
  or _86530_ (_36142_, _36140_, _36112_);
  and _86531_ (_36143_, _09310_, _08004_);
  or _86532_ (_36144_, _36100_, _06333_);
  or _86533_ (_36145_, _36144_, _36143_);
  and _86534_ (_36146_, _36145_, _06313_);
  and _86535_ (_36147_, _36146_, _36142_);
  and _86536_ (_36148_, _15251_, _08004_);
  or _86537_ (_36149_, _36148_, _36100_);
  and _86538_ (_36150_, _36149_, _06037_);
  or _86539_ (_36151_, _36150_, _06277_);
  or _86540_ (_36153_, _36151_, _36147_);
  and _86541_ (_36154_, _08004_, _09014_);
  or _86542_ (_36155_, _36154_, _36100_);
  or _86543_ (_36156_, _36155_, _06278_);
  and _86544_ (_36157_, _36156_, _36153_);
  or _86545_ (_36158_, _36157_, _06275_);
  and _86546_ (_36159_, _36158_, _36107_);
  or _86547_ (_36160_, _36159_, _06502_);
  and _86548_ (_36161_, _15266_, _08004_);
  or _86549_ (_36162_, _36100_, _07334_);
  or _86550_ (_36164_, _36162_, _36161_);
  and _86551_ (_36165_, _36164_, _07337_);
  and _86552_ (_36166_, _36165_, _36160_);
  or _86553_ (_36167_, _36166_, _36106_);
  and _86554_ (_36168_, _36167_, _07339_);
  or _86555_ (_36169_, _36100_, _08359_);
  and _86556_ (_36170_, _36155_, _06507_);
  and _86557_ (_36171_, _36170_, _36169_);
  or _86558_ (_36172_, _36171_, _36168_);
  and _86559_ (_36173_, _36172_, _12805_);
  and _86560_ (_36175_, _36116_, _06610_);
  and _86561_ (_36176_, _36175_, _36169_);
  nor _86562_ (_36177_, _16085_, _06018_);
  or _86563_ (_36178_, _36177_, _06509_);
  or _86564_ (_36179_, _36178_, _36176_);
  or _86565_ (_36180_, _36179_, _36173_);
  and _86566_ (_36181_, _15263_, _08004_);
  or _86567_ (_36182_, _36181_, _36100_);
  or _86568_ (_36183_, _36182_, _09107_);
  and _86569_ (_36184_, _36183_, _36180_);
  or _86570_ (_36186_, _36184_, _06602_);
  or _86571_ (_36187_, _36102_, _09112_);
  and _86572_ (_36188_, _36187_, _14116_);
  and _86573_ (_36189_, _36188_, _36186_);
  nor _86574_ (_36190_, _08698_, _06409_);
  or _86575_ (_36191_, _36190_, _08699_);
  and _86576_ (_36192_, _36191_, _06621_);
  or _86577_ (_36193_, _36192_, _07350_);
  or _86578_ (_36194_, _36193_, _36189_);
  and _86579_ (_36195_, _36194_, _36099_);
  or _86580_ (_36197_, _36195_, _06361_);
  or _86581_ (_36198_, _36191_, _06362_);
  and _86582_ (_36199_, _36198_, _07048_);
  and _86583_ (_36200_, _36199_, _36197_);
  and _86584_ (_36201_, _36114_, _06639_);
  or _86585_ (_36202_, _36201_, _07783_);
  or _86586_ (_36203_, _36202_, _36200_);
  and _86587_ (_36204_, _36203_, _36097_);
  or _86588_ (_36205_, _36204_, _06646_);
  and _86589_ (_36206_, _15321_, _08004_);
  or _86590_ (_36208_, _36100_, _06651_);
  or _86591_ (_36209_, _36208_, _36206_);
  and _86592_ (_36210_, _36209_, _01442_);
  and _86593_ (_36211_, _36210_, _36205_);
  or _86594_ (_36212_, _36211_, _36096_);
  and _86595_ (_44286_, _36212_, _43634_);
  nor _86596_ (_36213_, _01442_, _14048_);
  nor _86597_ (_36214_, _07688_, \oc8051_golden_model_1.SP [4]);
  nor _86598_ (_36215_, _36214_, _14011_);
  or _86599_ (_36216_, _36215_, _07367_);
  nor _86600_ (_36218_, _08004_, _14048_);
  nor _86601_ (_36219_, _10589_, _14023_);
  or _86602_ (_36220_, _36219_, _36218_);
  and _86603_ (_36221_, _08004_, \oc8051_golden_model_1.ACC [4]);
  nand _86604_ (_36222_, _36221_, _08599_);
  and _86605_ (_36223_, _36222_, _06615_);
  and _86606_ (_36224_, _36223_, _36220_);
  nor _86607_ (_36225_, _08596_, _14023_);
  or _86608_ (_36226_, _36218_, _14025_);
  or _86609_ (_36227_, _36226_, _36225_);
  and _86610_ (_36229_, _36227_, _14022_);
  and _86611_ (_36230_, _15367_, _08004_);
  or _86612_ (_36231_, _36230_, _36218_);
  or _86613_ (_36232_, _36231_, _07275_);
  or _86614_ (_36233_, _36221_, _36218_);
  and _86615_ (_36234_, _36233_, _07259_);
  nor _86616_ (_36235_, _07259_, _14048_);
  or _86617_ (_36236_, _36235_, _06816_);
  or _86618_ (_36237_, _36236_, _36234_);
  or _86619_ (_36238_, _36215_, _07564_);
  and _86620_ (_36240_, _36238_, _36237_);
  or _86621_ (_36241_, _36240_, _06474_);
  and _86622_ (_36242_, _36241_, _06052_);
  and _86623_ (_36243_, _36242_, _36232_);
  and _86624_ (_36244_, _36215_, _07692_);
  or _86625_ (_36245_, _36244_, _06410_);
  or _86626_ (_36246_, _36245_, _36243_);
  and _86627_ (_36247_, _14049_, _06342_);
  nor _86628_ (_36248_, _08700_, _14048_);
  nor _86629_ (_36249_, _36248_, _36247_);
  nand _86630_ (_36251_, _36249_, _06410_);
  and _86631_ (_36252_, _36251_, _36246_);
  or _86632_ (_36253_, _36252_, _06417_);
  or _86633_ (_36254_, _36233_, _06426_);
  and _86634_ (_36255_, _36254_, _07394_);
  and _86635_ (_36256_, _36255_, _36253_);
  and _86636_ (_36257_, _07689_, \oc8051_golden_model_1.SP [4]);
  nor _86637_ (_36258_, _07689_, \oc8051_golden_model_1.SP [4]);
  nor _86638_ (_36259_, _36258_, _36257_);
  and _86639_ (_36260_, _36259_, _06351_);
  or _86640_ (_36262_, _36260_, _14062_);
  or _86641_ (_36263_, _36262_, _36256_);
  or _86642_ (_36264_, _36215_, _07597_);
  and _86643_ (_36265_, _36264_, _36263_);
  and _86644_ (_36266_, _36265_, _06327_);
  or _86645_ (_36267_, _36266_, _36229_);
  and _86646_ (_36268_, _09264_, _08004_);
  or _86647_ (_36269_, _36218_, _06333_);
  or _86648_ (_36270_, _36269_, _36268_);
  and _86649_ (_36271_, _36270_, _06313_);
  and _86650_ (_36273_, _36271_, _36267_);
  and _86651_ (_36274_, _15452_, _08004_);
  or _86652_ (_36275_, _36274_, _36218_);
  and _86653_ (_36276_, _36275_, _06037_);
  or _86654_ (_36277_, _36276_, _06277_);
  or _86655_ (_36278_, _36277_, _36273_);
  and _86656_ (_36279_, _08995_, _08004_);
  or _86657_ (_36280_, _36279_, _36218_);
  or _86658_ (_36281_, _36280_, _06278_);
  and _86659_ (_36282_, _36281_, _36278_);
  or _86660_ (_36284_, _36282_, _06275_);
  or _86661_ (_36285_, _36215_, _06009_);
  and _86662_ (_36286_, _36285_, _36284_);
  or _86663_ (_36287_, _36286_, _06502_);
  and _86664_ (_36288_, _15345_, _08004_);
  or _86665_ (_36289_, _36218_, _07334_);
  or _86666_ (_36290_, _36289_, _36288_);
  and _86667_ (_36291_, _36290_, _07337_);
  and _86668_ (_36292_, _36291_, _36287_);
  or _86669_ (_36293_, _36292_, _36224_);
  and _86670_ (_36295_, _36293_, _07339_);
  or _86671_ (_36296_, _36218_, _08599_);
  and _86672_ (_36297_, _36280_, _06507_);
  and _86673_ (_36298_, _36297_, _36296_);
  or _86674_ (_36299_, _36298_, _36295_);
  and _86675_ (_36300_, _36299_, _12805_);
  and _86676_ (_36301_, _36233_, _06610_);
  and _86677_ (_36302_, _36301_, _36296_);
  and _86678_ (_36303_, _36215_, _07330_);
  or _86679_ (_36304_, _36303_, _06509_);
  or _86680_ (_36306_, _36304_, _36302_);
  or _86681_ (_36307_, _36306_, _36300_);
  and _86682_ (_36308_, _15342_, _08004_);
  or _86683_ (_36309_, _36308_, _36218_);
  or _86684_ (_36310_, _36309_, _09107_);
  and _86685_ (_36311_, _36310_, _36307_);
  or _86686_ (_36312_, _36311_, _06602_);
  or _86687_ (_36313_, _36220_, _09112_);
  and _86688_ (_36314_, _36313_, _14116_);
  and _86689_ (_36315_, _36314_, _36312_);
  nor _86690_ (_36317_, _08699_, _14048_);
  or _86691_ (_36318_, _36317_, _14049_);
  and _86692_ (_36319_, _36318_, _06621_);
  or _86693_ (_36320_, _36319_, _07350_);
  or _86694_ (_36321_, _36320_, _36315_);
  or _86695_ (_36322_, _36215_, _06016_);
  and _86696_ (_36323_, _36322_, _36321_);
  or _86697_ (_36324_, _36323_, _06361_);
  or _86698_ (_36325_, _36318_, _06362_);
  and _86699_ (_36326_, _36325_, _07048_);
  and _86700_ (_36328_, _36326_, _36324_);
  and _86701_ (_36329_, _36231_, _06639_);
  or _86702_ (_36330_, _36329_, _07783_);
  or _86703_ (_36331_, _36330_, _36328_);
  and _86704_ (_36332_, _36331_, _36216_);
  or _86705_ (_36333_, _36332_, _06646_);
  and _86706_ (_36334_, _15524_, _08004_);
  or _86707_ (_36335_, _36218_, _06651_);
  or _86708_ (_36336_, _36335_, _36334_);
  and _86709_ (_36337_, _36336_, _01442_);
  and _86710_ (_36339_, _36337_, _36333_);
  or _86711_ (_36340_, _36339_, _36213_);
  and _86712_ (_44287_, _36340_, _43634_);
  nor _86713_ (_36341_, _01442_, _14047_);
  nor _86714_ (_36342_, _14011_, \oc8051_golden_model_1.SP [5]);
  nor _86715_ (_36343_, _36342_, _14012_);
  or _86716_ (_36344_, _36343_, _07367_);
  or _86717_ (_36345_, _36343_, _06016_);
  nor _86718_ (_36346_, _08004_, _14047_);
  nor _86719_ (_36347_, _10570_, _14023_);
  or _86720_ (_36349_, _36347_, _36346_);
  and _86721_ (_36350_, _08004_, \oc8051_golden_model_1.ACC [5]);
  nand _86722_ (_36351_, _36350_, _08308_);
  and _86723_ (_36352_, _36351_, _06615_);
  and _86724_ (_36353_, _36352_, _36349_);
  nor _86725_ (_36354_, _08305_, _14023_);
  or _86726_ (_36355_, _36346_, _14025_);
  or _86727_ (_36356_, _36355_, _36354_);
  and _86728_ (_36357_, _36356_, _14022_);
  and _86729_ (_36358_, _15550_, _08004_);
  or _86730_ (_36360_, _36358_, _36346_);
  or _86731_ (_36361_, _36360_, _07275_);
  or _86732_ (_36362_, _36350_, _36346_);
  or _86733_ (_36363_, _36362_, _07260_);
  or _86734_ (_36364_, _07259_, \oc8051_golden_model_1.SP [5]);
  and _86735_ (_36365_, _36364_, _07564_);
  and _86736_ (_36366_, _36365_, _36363_);
  and _86737_ (_36367_, _36343_, _06816_);
  or _86738_ (_36368_, _36367_, _06474_);
  or _86739_ (_36369_, _36368_, _36366_);
  and _86740_ (_36371_, _36369_, _06052_);
  and _86741_ (_36372_, _36371_, _36361_);
  and _86742_ (_36373_, _36343_, _07692_);
  or _86743_ (_36374_, _36373_, _06410_);
  or _86744_ (_36375_, _36374_, _36372_);
  and _86745_ (_36376_, _14050_, _06342_);
  nor _86746_ (_36377_, _36247_, _14047_);
  nor _86747_ (_36378_, _36377_, _36376_);
  nand _86748_ (_36379_, _36378_, _06410_);
  and _86749_ (_36380_, _36379_, _36375_);
  or _86750_ (_36382_, _36380_, _06417_);
  or _86751_ (_36383_, _36362_, _06426_);
  and _86752_ (_36384_, _36383_, _07394_);
  and _86753_ (_36385_, _36384_, _36382_);
  nor _86754_ (_36386_, _36257_, \oc8051_golden_model_1.SP [5]);
  nor _86755_ (_36387_, _36386_, _14063_);
  and _86756_ (_36388_, _36387_, _06351_);
  or _86757_ (_36389_, _36388_, _14062_);
  or _86758_ (_36390_, _36389_, _36385_);
  or _86759_ (_36391_, _36343_, _07597_);
  and _86760_ (_36393_, _36391_, _36390_);
  and _86761_ (_36394_, _36393_, _06327_);
  or _86762_ (_36395_, _36394_, _36357_);
  and _86763_ (_36396_, _09218_, _08004_);
  or _86764_ (_36397_, _36346_, _06333_);
  or _86765_ (_36398_, _36397_, _36396_);
  and _86766_ (_36399_, _36398_, _06313_);
  and _86767_ (_36400_, _36399_, _36395_);
  and _86768_ (_36401_, _15649_, _08004_);
  or _86769_ (_36402_, _36401_, _36346_);
  and _86770_ (_36404_, _36402_, _06037_);
  or _86771_ (_36405_, _36404_, _06277_);
  or _86772_ (_36406_, _36405_, _36400_);
  and _86773_ (_36407_, _08954_, _08004_);
  or _86774_ (_36408_, _36407_, _36346_);
  or _86775_ (_36409_, _36408_, _06278_);
  and _86776_ (_36410_, _36409_, _36406_);
  or _86777_ (_36411_, _36410_, _06275_);
  or _86778_ (_36412_, _36343_, _06009_);
  and _86779_ (_36413_, _36412_, _36411_);
  or _86780_ (_36415_, _36413_, _06502_);
  and _86781_ (_36416_, _15664_, _08004_);
  or _86782_ (_36417_, _36346_, _07334_);
  or _86783_ (_36418_, _36417_, _36416_);
  and _86784_ (_36419_, _36418_, _07337_);
  and _86785_ (_36420_, _36419_, _36415_);
  or _86786_ (_36421_, _36420_, _36353_);
  and _86787_ (_36422_, _36421_, _07339_);
  or _86788_ (_36423_, _36346_, _08308_);
  and _86789_ (_36424_, _36408_, _06507_);
  and _86790_ (_36426_, _36424_, _36423_);
  or _86791_ (_36427_, _36426_, _36422_);
  and _86792_ (_36428_, _36427_, _12805_);
  and _86793_ (_36429_, _36362_, _06610_);
  and _86794_ (_36430_, _36429_, _36423_);
  and _86795_ (_36431_, _36343_, _07330_);
  or _86796_ (_36432_, _36431_, _06509_);
  or _86797_ (_36433_, _36432_, _36430_);
  or _86798_ (_36434_, _36433_, _36428_);
  and _86799_ (_36435_, _15663_, _08004_);
  or _86800_ (_36437_, _36346_, _09107_);
  or _86801_ (_36438_, _36437_, _36435_);
  and _86802_ (_36439_, _36438_, _36434_);
  or _86803_ (_36440_, _36439_, _06602_);
  or _86804_ (_36441_, _36349_, _09112_);
  and _86805_ (_36442_, _36441_, _14116_);
  and _86806_ (_36443_, _36442_, _36440_);
  nor _86807_ (_36444_, _14049_, _14047_);
  or _86808_ (_36445_, _36444_, _14050_);
  and _86809_ (_36446_, _36445_, _06621_);
  or _86810_ (_36448_, _36446_, _07350_);
  or _86811_ (_36449_, _36448_, _36443_);
  and _86812_ (_36450_, _36449_, _36345_);
  or _86813_ (_36451_, _36450_, _06361_);
  or _86814_ (_36452_, _36445_, _06362_);
  and _86815_ (_36453_, _36452_, _07048_);
  and _86816_ (_36454_, _36453_, _36451_);
  and _86817_ (_36455_, _36360_, _06639_);
  or _86818_ (_36456_, _36455_, _07783_);
  or _86819_ (_36457_, _36456_, _36454_);
  and _86820_ (_36459_, _36457_, _36344_);
  or _86821_ (_36460_, _36459_, _06646_);
  and _86822_ (_36461_, _15721_, _08004_);
  or _86823_ (_36462_, _36346_, _06651_);
  or _86824_ (_36463_, _36462_, _36461_);
  and _86825_ (_36464_, _36463_, _01442_);
  and _86826_ (_36465_, _36464_, _36460_);
  or _86827_ (_36466_, _36465_, _36341_);
  and _86828_ (_44288_, _36466_, _43634_);
  nor _86829_ (_36467_, _01442_, _14046_);
  nor _86830_ (_36469_, _08004_, _14046_);
  and _86831_ (_36470_, _15759_, _08004_);
  or _86832_ (_36471_, _36470_, _36469_);
  or _86833_ (_36472_, _36471_, _07275_);
  and _86834_ (_36473_, _08004_, \oc8051_golden_model_1.ACC [6]);
  or _86835_ (_36474_, _36473_, _36469_);
  or _86836_ (_36475_, _36474_, _07260_);
  or _86837_ (_36476_, _07259_, \oc8051_golden_model_1.SP [6]);
  and _86838_ (_36477_, _36476_, _07564_);
  and _86839_ (_36478_, _36477_, _36475_);
  nor _86840_ (_36480_, _14012_, \oc8051_golden_model_1.SP [6]);
  nor _86841_ (_36481_, _36480_, _14013_);
  and _86842_ (_36482_, _36481_, _06816_);
  or _86843_ (_36483_, _36482_, _06474_);
  or _86844_ (_36484_, _36483_, _36478_);
  and _86845_ (_36485_, _36484_, _06052_);
  and _86846_ (_36486_, _36485_, _36472_);
  and _86847_ (_36487_, _36481_, _07692_);
  or _86848_ (_36488_, _36487_, _06410_);
  or _86849_ (_36489_, _36488_, _36486_);
  nor _86850_ (_36491_, _36376_, _14046_);
  nor _86851_ (_36492_, _36491_, _14052_);
  nand _86852_ (_36493_, _36492_, _06410_);
  and _86853_ (_36494_, _36493_, _36489_);
  or _86854_ (_36495_, _36494_, _06417_);
  or _86855_ (_36496_, _36474_, _06426_);
  and _86856_ (_36497_, _36496_, _07394_);
  and _86857_ (_36498_, _36497_, _36495_);
  nor _86858_ (_36499_, _14063_, \oc8051_golden_model_1.SP [6]);
  nor _86859_ (_36500_, _36499_, _14064_);
  and _86860_ (_36502_, _36500_, _06351_);
  or _86861_ (_36503_, _36502_, _36498_);
  and _86862_ (_36504_, _36503_, _07597_);
  nand _86863_ (_36505_, _36481_, _14062_);
  nand _86864_ (_36506_, _36505_, _06327_);
  or _86865_ (_36507_, _36506_, _36504_);
  nor _86866_ (_36508_, _08209_, _14023_);
  or _86867_ (_36509_, _36469_, _06327_);
  or _86868_ (_36510_, _36509_, _36508_);
  and _86869_ (_36511_, _36510_, _36507_);
  or _86870_ (_36513_, _36511_, _09572_);
  and _86871_ (_36514_, _09172_, _08004_);
  or _86872_ (_36515_, _36469_, _06333_);
  or _86873_ (_36516_, _36515_, _36514_);
  and _86874_ (_36517_, _36516_, _06313_);
  and _86875_ (_36518_, _36517_, _36513_);
  and _86876_ (_36519_, _15846_, _08004_);
  or _86877_ (_36520_, _36519_, _36469_);
  and _86878_ (_36521_, _36520_, _06037_);
  or _86879_ (_36522_, _36521_, _06277_);
  or _86880_ (_36524_, _36522_, _36518_);
  and _86881_ (_36525_, _15853_, _08004_);
  or _86882_ (_36526_, _36525_, _36469_);
  or _86883_ (_36527_, _36526_, _06278_);
  and _86884_ (_36528_, _36527_, _36524_);
  or _86885_ (_36529_, _36528_, _06275_);
  or _86886_ (_36530_, _36481_, _06009_);
  and _86887_ (_36531_, _36530_, _36529_);
  or _86888_ (_36532_, _36531_, _06502_);
  and _86889_ (_36533_, _15862_, _08004_);
  or _86890_ (_36535_, _36469_, _07334_);
  or _86891_ (_36536_, _36535_, _36533_);
  and _86892_ (_36537_, _36536_, _07337_);
  and _86893_ (_36538_, _36537_, _36532_);
  and _86894_ (_36539_, _10596_, _08004_);
  or _86895_ (_36540_, _36539_, _36469_);
  and _86896_ (_36541_, _36540_, _06615_);
  or _86897_ (_36542_, _36541_, _36538_);
  and _86898_ (_36543_, _36542_, _07339_);
  or _86899_ (_36544_, _36469_, _08212_);
  and _86900_ (_36546_, _36526_, _06507_);
  and _86901_ (_36547_, _36546_, _36544_);
  or _86902_ (_36548_, _36547_, _36543_);
  and _86903_ (_36549_, _36548_, _12805_);
  and _86904_ (_36550_, _36474_, _06610_);
  and _86905_ (_36551_, _36550_, _36544_);
  and _86906_ (_36552_, _36481_, _07330_);
  or _86907_ (_36553_, _36552_, _06509_);
  or _86908_ (_36554_, _36553_, _36551_);
  or _86909_ (_36555_, _36554_, _36549_);
  and _86910_ (_36557_, _15859_, _08004_);
  or _86911_ (_36558_, _36469_, _09107_);
  or _86912_ (_36559_, _36558_, _36557_);
  and _86913_ (_36560_, _36559_, _36555_);
  or _86914_ (_36561_, _36560_, _06602_);
  nor _86915_ (_36562_, _10595_, _14023_);
  or _86916_ (_36563_, _36562_, _36469_);
  or _86917_ (_36564_, _36563_, _09112_);
  and _86918_ (_36565_, _36564_, _14116_);
  and _86919_ (_36566_, _36565_, _36561_);
  nor _86920_ (_36568_, _14050_, _14046_);
  or _86921_ (_36569_, _36568_, _14051_);
  and _86922_ (_36570_, _36569_, _06621_);
  or _86923_ (_36571_, _36570_, _07350_);
  or _86924_ (_36572_, _36571_, _36566_);
  nor _86925_ (_36573_, _36481_, _06016_);
  nor _86926_ (_36574_, _36573_, _06361_);
  and _86927_ (_36575_, _36574_, _36572_);
  and _86928_ (_36576_, _36569_, _06361_);
  or _86929_ (_36577_, _36576_, _06639_);
  or _86930_ (_36579_, _36577_, _36575_);
  or _86931_ (_36580_, _36471_, _07048_);
  and _86932_ (_36581_, _36580_, _07367_);
  and _86933_ (_36582_, _36581_, _36579_);
  and _86934_ (_36583_, _36481_, _07783_);
  or _86935_ (_36584_, _36583_, _06646_);
  or _86936_ (_36585_, _36584_, _36582_);
  and _86937_ (_36586_, _15921_, _08004_);
  or _86938_ (_36587_, _36469_, _06651_);
  or _86939_ (_36588_, _36587_, _36586_);
  and _86940_ (_36590_, _36588_, _01442_);
  and _86941_ (_36591_, _36590_, _36585_);
  or _86942_ (_36592_, _36591_, _36467_);
  and _86943_ (_44289_, _36592_, _43634_);
  and _86944_ (_36593_, _01446_, \oc8051_golden_model_1.SBUF [0]);
  and _86945_ (_36594_, _14145_, \oc8051_golden_model_1.SBUF [0]);
  nor _86946_ (_36595_, _08453_, _14145_);
  or _86947_ (_36596_, _36595_, _36594_);
  or _86948_ (_36597_, _36596_, _07275_);
  and _86949_ (_36598_, _07962_, \oc8051_golden_model_1.ACC [0]);
  or _86950_ (_36600_, _36598_, _36594_);
  and _86951_ (_36601_, _36600_, _07259_);
  and _86952_ (_36602_, _07260_, \oc8051_golden_model_1.SBUF [0]);
  or _86953_ (_36603_, _36602_, _06474_);
  or _86954_ (_36604_, _36603_, _36601_);
  and _86955_ (_36605_, _36604_, _06772_);
  and _86956_ (_36606_, _36605_, _36597_);
  and _86957_ (_36607_, _07962_, _07250_);
  or _86958_ (_36608_, _36607_, _36594_);
  and _86959_ (_36609_, _36608_, _06410_);
  or _86960_ (_36611_, _36609_, _36606_);
  and _86961_ (_36612_, _36611_, _06426_);
  and _86962_ (_36613_, _36600_, _06417_);
  or _86963_ (_36614_, _36613_, _10153_);
  or _86964_ (_36615_, _36614_, _36612_);
  or _86965_ (_36616_, _36608_, _06327_);
  and _86966_ (_36617_, _36616_, _36615_);
  or _86967_ (_36618_, _36617_, _09572_);
  and _86968_ (_36619_, _09447_, _07962_);
  or _86969_ (_36620_, _36594_, _06333_);
  or _86970_ (_36622_, _36620_, _36619_);
  and _86971_ (_36623_, _36622_, _36618_);
  or _86972_ (_36624_, _36623_, _06037_);
  and _86973_ (_36625_, _14666_, _07962_);
  or _86974_ (_36626_, _36594_, _06313_);
  or _86975_ (_36627_, _36626_, _36625_);
  and _86976_ (_36628_, _36627_, _06278_);
  and _86977_ (_36629_, _36628_, _36624_);
  and _86978_ (_36630_, _07962_, _09008_);
  or _86979_ (_36631_, _36630_, _36594_);
  and _86980_ (_36633_, _36631_, _06277_);
  or _86981_ (_36634_, _36633_, _06502_);
  or _86982_ (_36635_, _36634_, _36629_);
  and _86983_ (_36636_, _14566_, _07962_);
  or _86984_ (_36637_, _36594_, _07334_);
  or _86985_ (_36638_, _36637_, _36636_);
  and _86986_ (_36639_, _36638_, _07337_);
  and _86987_ (_36640_, _36639_, _36635_);
  nor _86988_ (_36641_, _12622_, _14145_);
  or _86989_ (_36642_, _36641_, _36594_);
  and _86990_ (_36644_, _10577_, _07962_);
  nor _86991_ (_36645_, _36644_, _07337_);
  and _86992_ (_36646_, _36645_, _36642_);
  or _86993_ (_36647_, _36646_, _36640_);
  and _86994_ (_36648_, _36647_, _07339_);
  nand _86995_ (_36649_, _36631_, _06507_);
  nor _86996_ (_36650_, _36649_, _36595_);
  or _86997_ (_36651_, _36650_, _06610_);
  or _86998_ (_36652_, _36651_, _36648_);
  or _86999_ (_36653_, _36644_, _36594_);
  or _87000_ (_36655_, _36653_, _07331_);
  and _87001_ (_36656_, _36655_, _36652_);
  or _87002_ (_36657_, _36656_, _06509_);
  and _87003_ (_36658_, _14563_, _07962_);
  or _87004_ (_36659_, _36594_, _09107_);
  or _87005_ (_36660_, _36659_, _36658_);
  and _87006_ (_36661_, _36660_, _09112_);
  and _87007_ (_36662_, _36661_, _36657_);
  and _87008_ (_36663_, _36642_, _06602_);
  or _87009_ (_36664_, _36663_, _19642_);
  or _87010_ (_36666_, _36664_, _36662_);
  or _87011_ (_36667_, _36596_, _19641_);
  and _87012_ (_36668_, _36667_, _01442_);
  and _87013_ (_36669_, _36668_, _36666_);
  or _87014_ (_36670_, _36669_, _36593_);
  and _87015_ (_44291_, _36670_, _43634_);
  and _87016_ (_36671_, _01446_, \oc8051_golden_model_1.SBUF [1]);
  or _87017_ (_36672_, _14851_, _14145_);
  or _87018_ (_36673_, _07962_, \oc8051_golden_model_1.SBUF [1]);
  and _87019_ (_36674_, _36673_, _06037_);
  and _87020_ (_36676_, _36674_, _36672_);
  and _87021_ (_36677_, _14744_, _07962_);
  not _87022_ (_36678_, _36677_);
  and _87023_ (_36679_, _36678_, _36673_);
  or _87024_ (_36680_, _36679_, _07275_);
  and _87025_ (_36681_, _14145_, \oc8051_golden_model_1.SBUF [1]);
  and _87026_ (_36682_, _07962_, \oc8051_golden_model_1.ACC [1]);
  or _87027_ (_36683_, _36682_, _36681_);
  and _87028_ (_36684_, _36683_, _07259_);
  and _87029_ (_36685_, _07260_, \oc8051_golden_model_1.SBUF [1]);
  or _87030_ (_36687_, _36685_, _06474_);
  or _87031_ (_36688_, _36687_, _36684_);
  and _87032_ (_36689_, _36688_, _06772_);
  and _87033_ (_36690_, _36689_, _36680_);
  nor _87034_ (_36691_, _14145_, _07448_);
  or _87035_ (_36692_, _36691_, _36681_);
  and _87036_ (_36693_, _36692_, _06410_);
  or _87037_ (_36694_, _36693_, _36690_);
  and _87038_ (_36695_, _36694_, _06426_);
  and _87039_ (_36696_, _36683_, _06417_);
  or _87040_ (_36698_, _36696_, _10153_);
  or _87041_ (_36699_, _36698_, _36695_);
  or _87042_ (_36700_, _36692_, _06327_);
  and _87043_ (_36701_, _36700_, _16672_);
  and _87044_ (_36702_, _36701_, _36699_);
  or _87045_ (_36703_, _09402_, _14145_);
  and _87046_ (_36704_, _36673_, _14025_);
  and _87047_ (_36705_, _36704_, _36703_);
  or _87048_ (_36706_, _36705_, _36702_);
  and _87049_ (_36707_, _36706_, _06313_);
  or _87050_ (_36709_, _36707_, _36676_);
  and _87051_ (_36710_, _36709_, _06278_);
  nand _87052_ (_36711_, _07962_, _07160_);
  and _87053_ (_36712_, _36673_, _06277_);
  and _87054_ (_36713_, _36712_, _36711_);
  or _87055_ (_36714_, _36713_, _36710_);
  and _87056_ (_36715_, _36714_, _07334_);
  or _87057_ (_36716_, _14749_, _14145_);
  and _87058_ (_36717_, _36673_, _06502_);
  and _87059_ (_36718_, _36717_, _36716_);
  or _87060_ (_36720_, _36718_, _06615_);
  or _87061_ (_36721_, _36720_, _36715_);
  and _87062_ (_36722_, _10579_, _07962_);
  or _87063_ (_36723_, _36722_, _36681_);
  or _87064_ (_36724_, _36723_, _07337_);
  and _87065_ (_36725_, _36724_, _07339_);
  and _87066_ (_36726_, _36725_, _36721_);
  or _87067_ (_36727_, _14747_, _14145_);
  and _87068_ (_36728_, _36673_, _06507_);
  and _87069_ (_36729_, _36728_, _36727_);
  or _87070_ (_36731_, _36729_, _06610_);
  or _87071_ (_36732_, _36731_, _36726_);
  and _87072_ (_36733_, _36682_, _08404_);
  or _87073_ (_36734_, _36681_, _07331_);
  or _87074_ (_36735_, _36734_, _36733_);
  and _87075_ (_36736_, _36735_, _09107_);
  and _87076_ (_36737_, _36736_, _36732_);
  or _87077_ (_36738_, _36711_, _08404_);
  and _87078_ (_36739_, _36673_, _06509_);
  and _87079_ (_36740_, _36739_, _36738_);
  or _87080_ (_36742_, _36740_, _06602_);
  or _87081_ (_36743_, _36742_, _36737_);
  nor _87082_ (_36744_, _10578_, _14145_);
  or _87083_ (_36745_, _36744_, _36681_);
  or _87084_ (_36746_, _36745_, _09112_);
  and _87085_ (_36747_, _36746_, _07048_);
  and _87086_ (_36748_, _36747_, _36743_);
  and _87087_ (_36749_, _36679_, _06639_);
  or _87088_ (_36750_, _36749_, _06646_);
  or _87089_ (_36751_, _36750_, _36748_);
  or _87090_ (_36753_, _36681_, _06651_);
  or _87091_ (_36754_, _36753_, _36677_);
  and _87092_ (_36755_, _36754_, _01442_);
  and _87093_ (_36756_, _36755_, _36751_);
  or _87094_ (_36757_, _36756_, _36671_);
  and _87095_ (_44292_, _36757_, _43634_);
  and _87096_ (_36758_, _01446_, \oc8051_golden_model_1.SBUF [2]);
  and _87097_ (_36759_, _14145_, \oc8051_golden_model_1.SBUF [2]);
  or _87098_ (_36760_, _36759_, _08503_);
  and _87099_ (_36761_, _07962_, _09057_);
  or _87100_ (_36763_, _36761_, _36759_);
  and _87101_ (_36764_, _36763_, _06507_);
  and _87102_ (_36765_, _36764_, _36760_);
  and _87103_ (_36766_, _09356_, _07962_);
  or _87104_ (_36767_, _36766_, _36759_);
  and _87105_ (_36768_, _36767_, _14025_);
  and _87106_ (_36769_, _14959_, _07962_);
  or _87107_ (_36770_, _36769_, _36759_);
  or _87108_ (_36771_, _36770_, _07275_);
  and _87109_ (_36772_, _07962_, \oc8051_golden_model_1.ACC [2]);
  or _87110_ (_36774_, _36772_, _36759_);
  and _87111_ (_36775_, _36774_, _07259_);
  and _87112_ (_36776_, _07260_, \oc8051_golden_model_1.SBUF [2]);
  or _87113_ (_36777_, _36776_, _06474_);
  or _87114_ (_36778_, _36777_, _36775_);
  and _87115_ (_36779_, _36778_, _06772_);
  and _87116_ (_36780_, _36779_, _36771_);
  nor _87117_ (_36781_, _14145_, _07854_);
  or _87118_ (_36782_, _36781_, _36759_);
  and _87119_ (_36783_, _36782_, _06410_);
  or _87120_ (_36785_, _36783_, _36780_);
  and _87121_ (_36786_, _36785_, _06426_);
  and _87122_ (_36787_, _36774_, _06417_);
  or _87123_ (_36788_, _36787_, _10153_);
  or _87124_ (_36789_, _36788_, _36786_);
  or _87125_ (_36790_, _36782_, _06327_);
  and _87126_ (_36791_, _36790_, _16672_);
  and _87127_ (_36792_, _36791_, _36789_);
  or _87128_ (_36793_, _36792_, _06037_);
  or _87129_ (_36794_, _36793_, _36768_);
  and _87130_ (_36796_, _15056_, _07962_);
  or _87131_ (_36797_, _36759_, _06313_);
  or _87132_ (_36798_, _36797_, _36796_);
  and _87133_ (_36799_, _36798_, _06278_);
  and _87134_ (_36800_, _36799_, _36794_);
  and _87135_ (_36801_, _36763_, _06277_);
  or _87136_ (_36802_, _36801_, _06502_);
  or _87137_ (_36803_, _36802_, _36800_);
  and _87138_ (_36804_, _14948_, _07962_);
  or _87139_ (_36805_, _36759_, _07334_);
  or _87140_ (_36807_, _36805_, _36804_);
  and _87141_ (_36808_, _36807_, _07337_);
  and _87142_ (_36809_, _36808_, _36803_);
  and _87143_ (_36810_, _10583_, _07962_);
  or _87144_ (_36811_, _36810_, _36759_);
  and _87145_ (_36812_, _36811_, _06615_);
  or _87146_ (_36813_, _36812_, _36809_);
  and _87147_ (_36814_, _36813_, _07339_);
  or _87148_ (_36815_, _36814_, _36765_);
  and _87149_ (_36816_, _36815_, _07331_);
  and _87150_ (_36818_, _36774_, _06610_);
  and _87151_ (_36819_, _36818_, _36760_);
  or _87152_ (_36820_, _36819_, _06509_);
  or _87153_ (_36821_, _36820_, _36816_);
  and _87154_ (_36822_, _14945_, _07962_);
  or _87155_ (_36823_, _36759_, _09107_);
  or _87156_ (_36824_, _36823_, _36822_);
  and _87157_ (_36825_, _36824_, _09112_);
  and _87158_ (_36826_, _36825_, _36821_);
  nor _87159_ (_36827_, _10582_, _14145_);
  or _87160_ (_36829_, _36827_, _36759_);
  and _87161_ (_36830_, _36829_, _06602_);
  or _87162_ (_36831_, _36830_, _36826_);
  and _87163_ (_36832_, _36831_, _07048_);
  and _87164_ (_36833_, _36770_, _06639_);
  or _87165_ (_36834_, _36833_, _06646_);
  or _87166_ (_36835_, _36834_, _36832_);
  and _87167_ (_36836_, _15129_, _07962_);
  or _87168_ (_36837_, _36759_, _06651_);
  or _87169_ (_36838_, _36837_, _36836_);
  and _87170_ (_36840_, _36838_, _01442_);
  and _87171_ (_36841_, _36840_, _36835_);
  or _87172_ (_36842_, _36841_, _36758_);
  and _87173_ (_44293_, _36842_, _43634_);
  and _87174_ (_36843_, _14145_, \oc8051_golden_model_1.SBUF [3]);
  or _87175_ (_36844_, _36843_, _08359_);
  and _87176_ (_36845_, _07962_, _09014_);
  or _87177_ (_36846_, _36845_, _36843_);
  and _87178_ (_36847_, _36846_, _06507_);
  and _87179_ (_36848_, _36847_, _36844_);
  nor _87180_ (_36849_, _10574_, _14145_);
  or _87181_ (_36850_, _36849_, _36843_);
  and _87182_ (_36851_, _07962_, \oc8051_golden_model_1.ACC [3]);
  nand _87183_ (_36852_, _36851_, _08359_);
  and _87184_ (_36853_, _36852_, _06615_);
  and _87185_ (_36854_, _36853_, _36850_);
  and _87186_ (_36855_, _15153_, _07962_);
  or _87187_ (_36856_, _36855_, _36843_);
  or _87188_ (_36857_, _36856_, _07275_);
  or _87189_ (_36858_, _36851_, _36843_);
  and _87190_ (_36860_, _36858_, _07259_);
  and _87191_ (_36861_, _07260_, \oc8051_golden_model_1.SBUF [3]);
  or _87192_ (_36862_, _36861_, _06474_);
  or _87193_ (_36863_, _36862_, _36860_);
  and _87194_ (_36864_, _36863_, _06772_);
  and _87195_ (_36865_, _36864_, _36857_);
  nor _87196_ (_36866_, _14145_, _07680_);
  or _87197_ (_36867_, _36866_, _36843_);
  and _87198_ (_36868_, _36867_, _06410_);
  or _87199_ (_36869_, _36868_, _36865_);
  and _87200_ (_36871_, _36869_, _06426_);
  and _87201_ (_36872_, _36858_, _06417_);
  or _87202_ (_36873_, _36872_, _10153_);
  or _87203_ (_36874_, _36873_, _36871_);
  and _87204_ (_36875_, _36867_, _16672_);
  or _87205_ (_36876_, _36875_, _06334_);
  and _87206_ (_36877_, _36876_, _36874_);
  and _87207_ (_36878_, _09310_, _07962_);
  or _87208_ (_36879_, _36878_, _36843_);
  and _87209_ (_36880_, _36879_, _09572_);
  or _87210_ (_36882_, _36880_, _36877_);
  or _87211_ (_36883_, _36882_, _06037_);
  and _87212_ (_36884_, _15251_, _07962_);
  or _87213_ (_36885_, _36843_, _06313_);
  or _87214_ (_36886_, _36885_, _36884_);
  and _87215_ (_36887_, _36886_, _06278_);
  and _87216_ (_36888_, _36887_, _36883_);
  and _87217_ (_36889_, _36846_, _06277_);
  or _87218_ (_36890_, _36889_, _06502_);
  or _87219_ (_36891_, _36890_, _36888_);
  and _87220_ (_36893_, _15266_, _07962_);
  or _87221_ (_36894_, _36843_, _07334_);
  or _87222_ (_36895_, _36894_, _36893_);
  and _87223_ (_36896_, _36895_, _07337_);
  and _87224_ (_36897_, _36896_, _36891_);
  or _87225_ (_36898_, _36897_, _36854_);
  and _87226_ (_36899_, _36898_, _07339_);
  or _87227_ (_36900_, _36899_, _36848_);
  and _87228_ (_36901_, _36900_, _07331_);
  and _87229_ (_36902_, _36858_, _06610_);
  and _87230_ (_36904_, _36902_, _36844_);
  or _87231_ (_36905_, _36904_, _06509_);
  or _87232_ (_36906_, _36905_, _36901_);
  and _87233_ (_36907_, _15263_, _07962_);
  or _87234_ (_36908_, _36843_, _09107_);
  or _87235_ (_36909_, _36908_, _36907_);
  and _87236_ (_36910_, _36909_, _09112_);
  and _87237_ (_36911_, _36910_, _36906_);
  and _87238_ (_36912_, _36850_, _06602_);
  or _87239_ (_36913_, _36912_, _06639_);
  or _87240_ (_36915_, _36913_, _36911_);
  or _87241_ (_36916_, _36856_, _07048_);
  and _87242_ (_36917_, _36916_, _06651_);
  and _87243_ (_36918_, _36917_, _36915_);
  and _87244_ (_36919_, _15321_, _07962_);
  or _87245_ (_36920_, _36919_, _36843_);
  and _87246_ (_36921_, _36920_, _06646_);
  or _87247_ (_36922_, _36921_, _01446_);
  or _87248_ (_36923_, _36922_, _36918_);
  or _87249_ (_36924_, _01442_, \oc8051_golden_model_1.SBUF [3]);
  and _87250_ (_36926_, _36924_, _43634_);
  and _87251_ (_44294_, _36926_, _36923_);
  and _87252_ (_36927_, _14145_, \oc8051_golden_model_1.SBUF [4]);
  or _87253_ (_36928_, _36927_, _08599_);
  and _87254_ (_36929_, _08995_, _07962_);
  or _87255_ (_36930_, _36929_, _36927_);
  and _87256_ (_36931_, _36930_, _06507_);
  and _87257_ (_36932_, _36931_, _36928_);
  and _87258_ (_36933_, _15345_, _07962_);
  or _87259_ (_36934_, _36933_, _36927_);
  and _87260_ (_36936_, _36934_, _06502_);
  and _87261_ (_36937_, _15452_, _07962_);
  or _87262_ (_36938_, _36927_, _06313_);
  or _87263_ (_36939_, _36938_, _36937_);
  and _87264_ (_36940_, _15367_, _07962_);
  or _87265_ (_36941_, _36940_, _36927_);
  or _87266_ (_36942_, _36941_, _07275_);
  and _87267_ (_36943_, _07962_, \oc8051_golden_model_1.ACC [4]);
  or _87268_ (_36944_, _36943_, _36927_);
  and _87269_ (_36945_, _36944_, _07259_);
  and _87270_ (_36947_, _07260_, \oc8051_golden_model_1.SBUF [4]);
  or _87271_ (_36948_, _36947_, _06474_);
  or _87272_ (_36949_, _36948_, _36945_);
  and _87273_ (_36950_, _36949_, _06772_);
  and _87274_ (_36951_, _36950_, _36942_);
  nor _87275_ (_36952_, _08596_, _14145_);
  or _87276_ (_36953_, _36952_, _36927_);
  and _87277_ (_36954_, _36953_, _06410_);
  or _87278_ (_36955_, _36954_, _36951_);
  and _87279_ (_36956_, _36955_, _06426_);
  and _87280_ (_36958_, _36944_, _06417_);
  or _87281_ (_36959_, _36958_, _10153_);
  or _87282_ (_36960_, _36959_, _36956_);
  and _87283_ (_36961_, _36953_, _16672_);
  or _87284_ (_36962_, _36961_, _06334_);
  and _87285_ (_36963_, _36962_, _36960_);
  and _87286_ (_36964_, _09264_, _07962_);
  or _87287_ (_36965_, _36964_, _36927_);
  and _87288_ (_36966_, _36965_, _09572_);
  or _87289_ (_36967_, _36966_, _06037_);
  or _87290_ (_36969_, _36967_, _36963_);
  and _87291_ (_36970_, _36969_, _36939_);
  or _87292_ (_36971_, _36970_, _06277_);
  or _87293_ (_36972_, _36930_, _06278_);
  and _87294_ (_36973_, _36972_, _07334_);
  and _87295_ (_36974_, _36973_, _36971_);
  or _87296_ (_36975_, _36974_, _36936_);
  and _87297_ (_36976_, _36975_, _07337_);
  and _87298_ (_36977_, _10590_, _07962_);
  or _87299_ (_36978_, _36977_, _36927_);
  and _87300_ (_36980_, _36978_, _06615_);
  or _87301_ (_36981_, _36980_, _36976_);
  and _87302_ (_36982_, _36981_, _07339_);
  or _87303_ (_36983_, _36982_, _36932_);
  and _87304_ (_36984_, _36983_, _07331_);
  and _87305_ (_36985_, _36944_, _06610_);
  and _87306_ (_36986_, _36985_, _36928_);
  or _87307_ (_36987_, _36986_, _06509_);
  or _87308_ (_36988_, _36987_, _36984_);
  and _87309_ (_36989_, _15342_, _07962_);
  or _87310_ (_36991_, _36927_, _09107_);
  or _87311_ (_36992_, _36991_, _36989_);
  and _87312_ (_36993_, _36992_, _09112_);
  and _87313_ (_36994_, _36993_, _36988_);
  nor _87314_ (_36995_, _10589_, _14145_);
  or _87315_ (_36996_, _36995_, _36927_);
  and _87316_ (_36997_, _36996_, _06602_);
  or _87317_ (_36998_, _36997_, _06639_);
  or _87318_ (_36999_, _36998_, _36994_);
  or _87319_ (_37000_, _36941_, _07048_);
  and _87320_ (_37002_, _37000_, _06651_);
  and _87321_ (_37003_, _37002_, _36999_);
  and _87322_ (_37004_, _15524_, _07962_);
  or _87323_ (_37005_, _37004_, _36927_);
  and _87324_ (_37006_, _37005_, _06646_);
  or _87325_ (_37007_, _37006_, _01446_);
  or _87326_ (_37008_, _37007_, _37003_);
  or _87327_ (_37009_, _01442_, \oc8051_golden_model_1.SBUF [4]);
  and _87328_ (_37010_, _37009_, _43634_);
  and _87329_ (_44295_, _37010_, _37008_);
  and _87330_ (_37012_, _14145_, \oc8051_golden_model_1.SBUF [5]);
  and _87331_ (_37013_, _15664_, _07962_);
  or _87332_ (_37014_, _37013_, _37012_);
  and _87333_ (_37015_, _37014_, _06502_);
  and _87334_ (_37016_, _15649_, _07962_);
  or _87335_ (_37017_, _37012_, _06313_);
  or _87336_ (_37018_, _37017_, _37016_);
  and _87337_ (_37019_, _15550_, _07962_);
  or _87338_ (_37020_, _37019_, _37012_);
  or _87339_ (_37021_, _37020_, _07275_);
  and _87340_ (_37023_, _07962_, \oc8051_golden_model_1.ACC [5]);
  or _87341_ (_37024_, _37023_, _37012_);
  and _87342_ (_37025_, _37024_, _07259_);
  and _87343_ (_37026_, _07260_, \oc8051_golden_model_1.SBUF [5]);
  or _87344_ (_37027_, _37026_, _06474_);
  or _87345_ (_37028_, _37027_, _37025_);
  and _87346_ (_37029_, _37028_, _06772_);
  and _87347_ (_37030_, _37029_, _37021_);
  nor _87348_ (_37031_, _08305_, _14145_);
  or _87349_ (_37032_, _37031_, _37012_);
  and _87350_ (_37034_, _37032_, _06410_);
  or _87351_ (_37035_, _37034_, _37030_);
  and _87352_ (_37036_, _37035_, _06426_);
  and _87353_ (_37037_, _37024_, _06417_);
  or _87354_ (_37038_, _37037_, _10153_);
  or _87355_ (_37039_, _37038_, _37036_);
  and _87356_ (_37040_, _37032_, _16672_);
  or _87357_ (_37041_, _37040_, _06334_);
  and _87358_ (_37042_, _37041_, _37039_);
  and _87359_ (_37043_, _09218_, _07962_);
  or _87360_ (_37045_, _37043_, _37012_);
  and _87361_ (_37046_, _37045_, _09572_);
  or _87362_ (_37047_, _37046_, _06037_);
  or _87363_ (_37048_, _37047_, _37042_);
  and _87364_ (_37049_, _37048_, _37018_);
  or _87365_ (_37050_, _37049_, _06277_);
  and _87366_ (_37051_, _08954_, _07962_);
  or _87367_ (_37052_, _37051_, _37012_);
  or _87368_ (_37053_, _37052_, _06278_);
  and _87369_ (_37054_, _37053_, _07334_);
  and _87370_ (_37056_, _37054_, _37050_);
  or _87371_ (_37057_, _37056_, _37015_);
  and _87372_ (_37058_, _37057_, _07337_);
  and _87373_ (_37059_, _12626_, _07962_);
  or _87374_ (_37060_, _37059_, _37012_);
  and _87375_ (_37061_, _37060_, _06615_);
  or _87376_ (_37062_, _37061_, _37058_);
  and _87377_ (_37063_, _37062_, _07339_);
  or _87378_ (_37064_, _37012_, _08308_);
  and _87379_ (_37065_, _37052_, _06507_);
  and _87380_ (_37067_, _37065_, _37064_);
  or _87381_ (_37068_, _37067_, _37063_);
  and _87382_ (_37069_, _37068_, _07331_);
  and _87383_ (_37070_, _37024_, _06610_);
  and _87384_ (_37071_, _37070_, _37064_);
  or _87385_ (_37072_, _37071_, _06509_);
  or _87386_ (_37073_, _37072_, _37069_);
  and _87387_ (_37074_, _15663_, _07962_);
  or _87388_ (_37075_, _37012_, _09107_);
  or _87389_ (_37076_, _37075_, _37074_);
  and _87390_ (_37078_, _37076_, _09112_);
  and _87391_ (_37079_, _37078_, _37073_);
  nor _87392_ (_37080_, _10570_, _14145_);
  or _87393_ (_37081_, _37080_, _37012_);
  and _87394_ (_37082_, _37081_, _06602_);
  or _87395_ (_37083_, _37082_, _06639_);
  or _87396_ (_37084_, _37083_, _37079_);
  or _87397_ (_37085_, _37020_, _07048_);
  and _87398_ (_37086_, _37085_, _06651_);
  and _87399_ (_37087_, _37086_, _37084_);
  and _87400_ (_37089_, _15721_, _07962_);
  or _87401_ (_37090_, _37089_, _37012_);
  and _87402_ (_37091_, _37090_, _06646_);
  or _87403_ (_37092_, _37091_, _01446_);
  or _87404_ (_37093_, _37092_, _37087_);
  or _87405_ (_37094_, _01442_, \oc8051_golden_model_1.SBUF [5]);
  and _87406_ (_37095_, _37094_, _43634_);
  and _87407_ (_44296_, _37095_, _37093_);
  and _87408_ (_37096_, _14145_, \oc8051_golden_model_1.SBUF [6]);
  and _87409_ (_37097_, _15862_, _07962_);
  or _87410_ (_37099_, _37097_, _37096_);
  and _87411_ (_37100_, _37099_, _06502_);
  and _87412_ (_37101_, _15846_, _07962_);
  or _87413_ (_37102_, _37096_, _06313_);
  or _87414_ (_37103_, _37102_, _37101_);
  nor _87415_ (_37104_, _08209_, _14145_);
  or _87416_ (_37105_, _37104_, _37096_);
  or _87417_ (_37106_, _37105_, _06327_);
  and _87418_ (_37107_, _15759_, _07962_);
  or _87419_ (_37108_, _37107_, _37096_);
  or _87420_ (_37110_, _37108_, _07275_);
  and _87421_ (_37111_, _07962_, \oc8051_golden_model_1.ACC [6]);
  or _87422_ (_37112_, _37111_, _37096_);
  and _87423_ (_37113_, _37112_, _07259_);
  and _87424_ (_37114_, _07260_, \oc8051_golden_model_1.SBUF [6]);
  or _87425_ (_37115_, _37114_, _06474_);
  or _87426_ (_37116_, _37115_, _37113_);
  and _87427_ (_37117_, _37116_, _06772_);
  and _87428_ (_37118_, _37117_, _37110_);
  and _87429_ (_37119_, _37105_, _06410_);
  or _87430_ (_37121_, _37119_, _37118_);
  and _87431_ (_37122_, _37121_, _06426_);
  and _87432_ (_37123_, _37112_, _06417_);
  or _87433_ (_37124_, _37123_, _10153_);
  or _87434_ (_37125_, _37124_, _37122_);
  and _87435_ (_37126_, _37125_, _06333_);
  and _87436_ (_37127_, _37126_, _37106_);
  and _87437_ (_37128_, _09172_, _07962_);
  or _87438_ (_37129_, _37128_, _37096_);
  and _87439_ (_37130_, _37129_, _09572_);
  or _87440_ (_37132_, _37130_, _06037_);
  or _87441_ (_37133_, _37132_, _37127_);
  and _87442_ (_37134_, _37133_, _37103_);
  or _87443_ (_37135_, _37134_, _06277_);
  and _87444_ (_37136_, _15853_, _07962_);
  or _87445_ (_37137_, _37136_, _37096_);
  or _87446_ (_37138_, _37137_, _06278_);
  and _87447_ (_37139_, _37138_, _07334_);
  and _87448_ (_37140_, _37139_, _37135_);
  or _87449_ (_37141_, _37140_, _37100_);
  and _87450_ (_37143_, _37141_, _07337_);
  nor _87451_ (_37144_, _10595_, _14145_);
  or _87452_ (_37145_, _37144_, _37096_);
  nand _87453_ (_37146_, _37111_, _08212_);
  and _87454_ (_37147_, _37146_, _06615_);
  and _87455_ (_37148_, _37147_, _37145_);
  or _87456_ (_37149_, _37148_, _37143_);
  and _87457_ (_37150_, _37149_, _07339_);
  or _87458_ (_37151_, _37096_, _08212_);
  and _87459_ (_37152_, _37137_, _06507_);
  and _87460_ (_37154_, _37152_, _37151_);
  or _87461_ (_37155_, _37154_, _37150_);
  and _87462_ (_37156_, _37155_, _07331_);
  and _87463_ (_37157_, _37112_, _06610_);
  and _87464_ (_37158_, _37157_, _37151_);
  or _87465_ (_37159_, _37158_, _06509_);
  or _87466_ (_37160_, _37159_, _37156_);
  and _87467_ (_37161_, _15859_, _07962_);
  or _87468_ (_37162_, _37096_, _09107_);
  or _87469_ (_37163_, _37162_, _37161_);
  and _87470_ (_37165_, _37163_, _09112_);
  and _87471_ (_37166_, _37165_, _37160_);
  and _87472_ (_37167_, _37145_, _06602_);
  or _87473_ (_37168_, _37167_, _06639_);
  or _87474_ (_37169_, _37168_, _37166_);
  or _87475_ (_37170_, _37108_, _07048_);
  and _87476_ (_37171_, _37170_, _06651_);
  and _87477_ (_37172_, _37171_, _37169_);
  and _87478_ (_37173_, _15921_, _07962_);
  or _87479_ (_37174_, _37173_, _37096_);
  and _87480_ (_37176_, _37174_, _06646_);
  or _87481_ (_37177_, _37176_, _01446_);
  or _87482_ (_37178_, _37177_, _37172_);
  or _87483_ (_37179_, _01442_, \oc8051_golden_model_1.SBUF [6]);
  and _87484_ (_37180_, _37179_, _43634_);
  and _87485_ (_44297_, _37180_, _37178_);
  and _87486_ (_37181_, _01446_, \oc8051_golden_model_1.PSW [0]);
  and _87487_ (_37182_, _14239_, \oc8051_golden_model_1.PSW [0]);
  nor _87488_ (_37183_, _12622_, _14239_);
  or _87489_ (_37184_, _37183_, _37182_);
  and _87490_ (_37186_, _10577_, _08014_);
  nor _87491_ (_37187_, _37186_, _07337_);
  and _87492_ (_37188_, _37187_, _37184_);
  and _87493_ (_37189_, _14566_, _08014_);
  or _87494_ (_37190_, _37189_, _37182_);
  and _87495_ (_37191_, _37190_, _06502_);
  and _87496_ (_37192_, _14666_, _08014_);
  or _87497_ (_37193_, _37182_, _06313_);
  or _87498_ (_37194_, _37193_, _37192_);
  and _87499_ (_37195_, _09447_, _08014_);
  or _87500_ (_37197_, _37195_, _37182_);
  and _87501_ (_37198_, _37197_, _09572_);
  nor _87502_ (_37199_, _08453_, _14239_);
  or _87503_ (_37200_, _37199_, _37182_);
  or _87504_ (_37201_, _37200_, _07275_);
  and _87505_ (_37202_, _08014_, \oc8051_golden_model_1.ACC [0]);
  or _87506_ (_37203_, _37202_, _37182_);
  and _87507_ (_37204_, _37203_, _07259_);
  and _87508_ (_37205_, _07260_, \oc8051_golden_model_1.PSW [0]);
  or _87509_ (_37206_, _37205_, _06474_);
  or _87510_ (_37208_, _37206_, _37204_);
  and _87511_ (_37209_, _37208_, _06357_);
  and _87512_ (_37210_, _37209_, _37201_);
  not _87513_ (_37211_, _08640_);
  and _87514_ (_37212_, _37211_, \oc8051_golden_model_1.PSW [0]);
  and _87515_ (_37213_, _14581_, _08640_);
  or _87516_ (_37214_, _37213_, _37212_);
  and _87517_ (_37215_, _37214_, _06356_);
  or _87518_ (_37216_, _37215_, _37210_);
  and _87519_ (_37217_, _37216_, _06772_);
  and _87520_ (_37219_, _08014_, _07250_);
  or _87521_ (_37220_, _37219_, _37182_);
  and _87522_ (_37221_, _37220_, _06410_);
  or _87523_ (_37222_, _37221_, _06417_);
  or _87524_ (_37223_, _37222_, _37217_);
  or _87525_ (_37224_, _37203_, _06426_);
  and _87526_ (_37225_, _37224_, _06353_);
  and _87527_ (_37226_, _37225_, _37223_);
  and _87528_ (_37227_, _37182_, _06352_);
  or _87529_ (_37228_, _37227_, _06345_);
  or _87530_ (_37230_, _37228_, _37226_);
  or _87531_ (_37231_, _37200_, _06346_);
  and _87532_ (_37232_, _37231_, _06340_);
  and _87533_ (_37233_, _37232_, _37230_);
  or _87534_ (_37234_, _37212_, _16663_);
  and _87535_ (_37235_, _37234_, _06339_);
  and _87536_ (_37236_, _37235_, _37214_);
  or _87537_ (_37237_, _37236_, _10153_);
  or _87538_ (_37238_, _37237_, _37233_);
  and _87539_ (_37239_, _37220_, _06333_);
  or _87540_ (_37241_, _37239_, _06334_);
  and _87541_ (_37242_, _37241_, _37238_);
  or _87542_ (_37243_, _37242_, _06037_);
  or _87543_ (_37244_, _37243_, _37198_);
  and _87544_ (_37245_, _37244_, _37194_);
  or _87545_ (_37246_, _37245_, _06277_);
  and _87546_ (_37247_, _08014_, _09008_);
  or _87547_ (_37248_, _37247_, _37182_);
  or _87548_ (_37249_, _37248_, _06278_);
  and _87549_ (_37250_, _37249_, _07334_);
  and _87550_ (_37252_, _37250_, _37246_);
  or _87551_ (_37253_, _37252_, _37191_);
  and _87552_ (_37254_, _37253_, _07337_);
  or _87553_ (_37255_, _37254_, _37188_);
  and _87554_ (_37256_, _37255_, _07339_);
  nand _87555_ (_37257_, _37248_, _06507_);
  nor _87556_ (_37258_, _37257_, _37199_);
  or _87557_ (_37259_, _37258_, _06610_);
  or _87558_ (_37260_, _37259_, _37256_);
  or _87559_ (_37261_, _37186_, _37182_);
  or _87560_ (_37263_, _37261_, _07331_);
  and _87561_ (_37264_, _37263_, _37260_);
  or _87562_ (_37265_, _37264_, _06509_);
  and _87563_ (_37266_, _14563_, _08014_);
  or _87564_ (_37267_, _37182_, _09107_);
  or _87565_ (_37268_, _37267_, _37266_);
  and _87566_ (_37269_, _37268_, _09112_);
  and _87567_ (_37270_, _37269_, _37265_);
  and _87568_ (_37271_, _37184_, _06602_);
  or _87569_ (_37272_, _37271_, _06639_);
  or _87570_ (_37274_, _37272_, _37270_);
  or _87571_ (_37275_, _37200_, _07048_);
  and _87572_ (_37276_, _37275_, _37274_);
  or _87573_ (_37277_, _37276_, _05989_);
  or _87574_ (_37278_, _37182_, _05990_);
  and _87575_ (_37279_, _37278_, _37277_);
  or _87576_ (_37280_, _37279_, _06646_);
  or _87577_ (_37281_, _37200_, _06651_);
  and _87578_ (_37282_, _37281_, _01442_);
  and _87579_ (_37283_, _37282_, _37280_);
  or _87580_ (_37285_, _37283_, _37181_);
  and _87581_ (_44299_, _37285_, _43634_);
  not _87582_ (_37286_, \oc8051_golden_model_1.PSW [1]);
  nor _87583_ (_37287_, _01442_, _37286_);
  nor _87584_ (_37288_, _08014_, _37286_);
  nor _87585_ (_37289_, _10578_, _14239_);
  or _87586_ (_37290_, _37289_, _37288_);
  or _87587_ (_37291_, _37290_, _09112_);
  nand _87588_ (_37292_, _08014_, _07160_);
  or _87589_ (_37293_, _08014_, \oc8051_golden_model_1.PSW [1]);
  and _87590_ (_37295_, _37293_, _06277_);
  and _87591_ (_37296_, _37295_, _37292_);
  or _87592_ (_37297_, _14851_, _14239_);
  and _87593_ (_37298_, _37293_, _06037_);
  and _87594_ (_37299_, _37298_, _37297_);
  nor _87595_ (_37300_, _14239_, _07448_);
  or _87596_ (_37301_, _37300_, _37288_);
  or _87597_ (_37302_, _37301_, _06327_);
  and _87598_ (_37303_, _14796_, _08640_);
  nor _87599_ (_37304_, _08640_, _37286_);
  or _87600_ (_37306_, _37304_, _06340_);
  or _87601_ (_37307_, _37306_, _37303_);
  and _87602_ (_37308_, _14754_, _08640_);
  or _87603_ (_37309_, _37308_, _37304_);
  and _87604_ (_37310_, _37309_, _06352_);
  or _87605_ (_37311_, _37301_, _06772_);
  and _87606_ (_37312_, _14744_, _08014_);
  not _87607_ (_37313_, _37312_);
  and _87608_ (_37314_, _37313_, _37293_);
  or _87609_ (_37315_, _37314_, _07275_);
  and _87610_ (_37317_, _08014_, \oc8051_golden_model_1.ACC [1]);
  or _87611_ (_37318_, _37317_, _37288_);
  and _87612_ (_37319_, _37318_, _07259_);
  nor _87613_ (_37320_, _07259_, _37286_);
  or _87614_ (_37321_, _37320_, _06474_);
  or _87615_ (_37322_, _37321_, _37319_);
  and _87616_ (_37323_, _37322_, _06357_);
  and _87617_ (_37324_, _37323_, _37315_);
  and _87618_ (_37325_, _14767_, _08640_);
  or _87619_ (_37326_, _37325_, _37304_);
  and _87620_ (_37328_, _37326_, _06356_);
  or _87621_ (_37329_, _37328_, _06410_);
  or _87622_ (_37330_, _37329_, _37324_);
  and _87623_ (_37331_, _37330_, _37311_);
  or _87624_ (_37332_, _37331_, _06417_);
  or _87625_ (_37333_, _37318_, _06426_);
  and _87626_ (_37334_, _37333_, _06353_);
  and _87627_ (_37335_, _37334_, _37332_);
  or _87628_ (_37336_, _37335_, _37310_);
  and _87629_ (_37337_, _37336_, _06346_);
  and _87630_ (_37339_, _37325_, _14782_);
  or _87631_ (_37340_, _37339_, _37304_);
  and _87632_ (_37341_, _37340_, _06345_);
  or _87633_ (_37342_, _37341_, _06339_);
  or _87634_ (_37343_, _37342_, _37337_);
  and _87635_ (_37344_, _37343_, _37307_);
  or _87636_ (_37345_, _37344_, _10153_);
  and _87637_ (_37346_, _37345_, _37302_);
  or _87638_ (_37347_, _37346_, _09572_);
  and _87639_ (_37348_, _09402_, _08014_);
  or _87640_ (_37350_, _37288_, _06333_);
  or _87641_ (_37351_, _37350_, _37348_);
  and _87642_ (_37352_, _37351_, _06313_);
  and _87643_ (_37353_, _37352_, _37347_);
  or _87644_ (_37354_, _37353_, _37299_);
  and _87645_ (_37355_, _37354_, _06278_);
  or _87646_ (_37356_, _37355_, _37296_);
  and _87647_ (_37357_, _37356_, _07334_);
  or _87648_ (_37358_, _14749_, _14239_);
  and _87649_ (_37359_, _37293_, _06502_);
  and _87650_ (_37361_, _37359_, _37358_);
  or _87651_ (_37362_, _37361_, _06615_);
  or _87652_ (_37363_, _37362_, _37357_);
  nand _87653_ (_37364_, _10576_, _08014_);
  and _87654_ (_37365_, _37364_, _37290_);
  or _87655_ (_37366_, _37365_, _07337_);
  and _87656_ (_37367_, _37366_, _07339_);
  and _87657_ (_37368_, _37367_, _37363_);
  or _87658_ (_37369_, _14747_, _14239_);
  and _87659_ (_37370_, _37293_, _06507_);
  and _87660_ (_37372_, _37370_, _37369_);
  or _87661_ (_37373_, _37372_, _06610_);
  or _87662_ (_37374_, _37373_, _37368_);
  nor _87663_ (_37375_, _37288_, _07331_);
  nand _87664_ (_37376_, _37375_, _37364_);
  and _87665_ (_37377_, _37376_, _09107_);
  and _87666_ (_37378_, _37377_, _37374_);
  or _87667_ (_37379_, _37292_, _08404_);
  and _87668_ (_37380_, _37293_, _06509_);
  and _87669_ (_37381_, _37380_, _37379_);
  or _87670_ (_37383_, _37381_, _06602_);
  or _87671_ (_37384_, _37383_, _37378_);
  and _87672_ (_37385_, _37384_, _37291_);
  or _87673_ (_37386_, _37385_, _06639_);
  or _87674_ (_37387_, _37314_, _07048_);
  and _87675_ (_37388_, _37387_, _05990_);
  and _87676_ (_37389_, _37388_, _37386_);
  and _87677_ (_37390_, _37309_, _05989_);
  or _87678_ (_37391_, _37390_, _06646_);
  or _87679_ (_37392_, _37391_, _37389_);
  or _87680_ (_37394_, _37288_, _06651_);
  or _87681_ (_37395_, _37394_, _37312_);
  and _87682_ (_37396_, _37395_, _01442_);
  and _87683_ (_37397_, _37396_, _37392_);
  or _87684_ (_37398_, _37397_, _37287_);
  and _87685_ (_44300_, _37398_, _43634_);
  and _87686_ (_37399_, _01446_, \oc8051_golden_model_1.PSW [2]);
  not _87687_ (_37400_, _11058_);
  nand _87688_ (_37401_, _11326_, _37400_);
  or _87689_ (_37402_, _11326_, _11057_);
  and _87690_ (_37404_, _37402_, _37401_);
  or _87691_ (_37405_, _37404_, _17691_);
  and _87692_ (_37406_, _10183_, _10179_);
  and _87693_ (_37407_, _37406_, _10166_);
  and _87694_ (_37408_, _14239_, \oc8051_golden_model_1.PSW [2]);
  and _87695_ (_37409_, _09356_, _08014_);
  or _87696_ (_37410_, _37409_, _37408_);
  and _87697_ (_37411_, _37410_, _06332_);
  not _87698_ (_37412_, _10922_);
  nor _87699_ (_37413_, _10857_, _37400_);
  nor _87700_ (_37415_, _10858_, \oc8051_golden_model_1.ACC [7]);
  or _87701_ (_37416_, _37415_, _37413_);
  nor _87702_ (_37417_, _37416_, _14247_);
  and _87703_ (_37418_, _37416_, _14247_);
  nor _87704_ (_37419_, _37418_, _37417_);
  nor _87705_ (_37420_, _37419_, _37412_);
  and _87706_ (_37421_, _37419_, _37412_);
  or _87707_ (_37422_, _37421_, _37420_);
  or _87708_ (_37423_, _37422_, _10854_);
  and _87709_ (_37424_, _37211_, \oc8051_golden_model_1.PSW [2]);
  and _87710_ (_37426_, _14953_, _08640_);
  or _87711_ (_37427_, _37426_, _37424_);
  and _87712_ (_37428_, _37427_, _06352_);
  nor _87713_ (_37429_, _14239_, _07854_);
  or _87714_ (_37430_, _37429_, _37408_);
  or _87715_ (_37431_, _37430_, _06772_);
  and _87716_ (_37432_, _14959_, _08014_);
  or _87717_ (_37433_, _37432_, _37408_);
  or _87718_ (_37434_, _37433_, _07275_);
  and _87719_ (_37435_, _08014_, \oc8051_golden_model_1.ACC [2]);
  or _87720_ (_37437_, _37435_, _37408_);
  and _87721_ (_37438_, _37437_, _07259_);
  and _87722_ (_37439_, _07260_, \oc8051_golden_model_1.PSW [2]);
  or _87723_ (_37440_, _37439_, _06474_);
  or _87724_ (_37441_, _37440_, _37438_);
  and _87725_ (_37442_, _37441_, _06357_);
  and _87726_ (_37443_, _37442_, _37434_);
  and _87727_ (_37444_, _14955_, _08640_);
  or _87728_ (_37445_, _37444_, _37424_);
  and _87729_ (_37446_, _37445_, _06356_);
  or _87730_ (_37448_, _37446_, _06410_);
  or _87731_ (_37449_, _37448_, _37443_);
  and _87732_ (_37450_, _37449_, _37431_);
  or _87733_ (_37451_, _37450_, _06417_);
  or _87734_ (_37452_, _37437_, _06426_);
  and _87735_ (_37453_, _37452_, _06353_);
  and _87736_ (_37454_, _37453_, _37451_);
  or _87737_ (_37455_, _37454_, _37428_);
  and _87738_ (_37456_, _37455_, _06346_);
  and _87739_ (_37457_, _37444_, _14986_);
  or _87740_ (_37459_, _37457_, _37424_);
  and _87741_ (_37460_, _37459_, _06345_);
  or _87742_ (_37461_, _37460_, _37456_);
  and _87743_ (_37462_, _37461_, _09612_);
  or _87744_ (_37463_, _16775_, _16659_);
  or _87745_ (_37464_, _37463_, _16887_);
  or _87746_ (_37465_, _37464_, _17012_);
  or _87747_ (_37466_, _37465_, _17129_);
  or _87748_ (_37467_, _37466_, _17238_);
  or _87749_ (_37468_, _37467_, _10149_);
  or _87750_ (_37470_, _37468_, _17359_);
  and _87751_ (_37471_, _37470_, _09606_);
  or _87752_ (_37472_, _37471_, _12338_);
  or _87753_ (_37473_, _37472_, _37462_);
  not _87754_ (_37474_, _10851_);
  nor _87755_ (_37475_, _10793_, _08107_);
  nor _87756_ (_37476_, _37475_, \oc8051_golden_model_1.ACC [7]);
  not _87757_ (_37477_, _10612_);
  nor _87758_ (_37478_, _10793_, _37477_);
  or _87759_ (_37479_, _37478_, _37476_);
  and _87760_ (_37481_, _37479_, _14401_);
  nor _87761_ (_37482_, _37479_, _14401_);
  nor _87762_ (_37483_, _37482_, _37481_);
  nor _87763_ (_37484_, _37483_, _37474_);
  and _87764_ (_37485_, _37483_, _37474_);
  or _87765_ (_37486_, _37485_, _10784_);
  or _87766_ (_37487_, _37486_, _37484_);
  and _87767_ (_37488_, _37487_, _37473_);
  or _87768_ (_37489_, _37488_, _10853_);
  and _87769_ (_37490_, _37489_, _06458_);
  and _87770_ (_37492_, _37490_, _37423_);
  nor _87771_ (_37493_, _14411_, _14520_);
  nor _87772_ (_37494_, _10626_, \oc8051_golden_model_1.ACC [7]);
  or _87773_ (_37495_, _37494_, _37493_);
  or _87774_ (_37496_, _37495_, _14417_);
  nand _87775_ (_37497_, _37495_, _14417_);
  and _87776_ (_37498_, _37497_, _37496_);
  and _87777_ (_37499_, _37498_, _10690_);
  nor _87778_ (_37500_, _37498_, _10690_);
  or _87779_ (_37501_, _37500_, _37499_);
  and _87780_ (_37503_, _37501_, _06453_);
  or _87781_ (_37504_, _37503_, _37492_);
  or _87782_ (_37505_, _37504_, _10623_);
  nor _87783_ (_37506_, _10929_, _14526_);
  nor _87784_ (_37507_, _10930_, \oc8051_golden_model_1.ACC [7]);
  nor _87785_ (_37508_, _37507_, _37506_);
  not _87786_ (_37509_, _37508_);
  or _87787_ (_37510_, _37509_, _14428_);
  nand _87788_ (_37511_, _37509_, _14428_);
  and _87789_ (_37512_, _37511_, _37510_);
  and _87790_ (_37514_, _37512_, _10996_);
  nor _87791_ (_37515_, _37512_, _10996_);
  or _87792_ (_37516_, _37515_, _37514_);
  or _87793_ (_37517_, _37516_, _10624_);
  and _87794_ (_37518_, _37517_, _06340_);
  and _87795_ (_37519_, _37518_, _37505_);
  and _87796_ (_37520_, _15000_, _08640_);
  or _87797_ (_37521_, _37520_, _37424_);
  and _87798_ (_37522_, _37521_, _06339_);
  or _87799_ (_37523_, _37522_, _10153_);
  or _87800_ (_37525_, _37523_, _37519_);
  nor _87801_ (_37526_, _37430_, _06327_);
  nor _87802_ (_37527_, _37526_, _06332_);
  and _87803_ (_37528_, _37527_, _37525_);
  nor _87804_ (_37529_, _37528_, _37411_);
  nor _87805_ (_37530_, _37529_, _06330_);
  and _87806_ (_37531_, _37410_, _06330_);
  or _87807_ (_37532_, _37531_, _06037_);
  or _87808_ (_37533_, _37532_, _37530_);
  and _87809_ (_37534_, _15056_, _08014_);
  or _87810_ (_37536_, _37408_, _06313_);
  or _87811_ (_37537_, _37536_, _37534_);
  and _87812_ (_37538_, _37537_, _10172_);
  and _87813_ (_37539_, _37538_, _37533_);
  or _87814_ (_37540_, _37539_, _37407_);
  and _87815_ (_37541_, _37540_, _06278_);
  and _87816_ (_37542_, _08014_, _09057_);
  or _87817_ (_37543_, _37542_, _37408_);
  and _87818_ (_37544_, _37543_, _06277_);
  or _87819_ (_37545_, _37544_, _06502_);
  or _87820_ (_37547_, _37545_, _37541_);
  and _87821_ (_37548_, _14948_, _08014_);
  or _87822_ (_37549_, _37408_, _07334_);
  or _87823_ (_37550_, _37549_, _37548_);
  and _87824_ (_37551_, _37550_, _07337_);
  and _87825_ (_37552_, _37551_, _37547_);
  and _87826_ (_37553_, _10583_, _08014_);
  or _87827_ (_37554_, _37553_, _37408_);
  and _87828_ (_37555_, _37554_, _06615_);
  or _87829_ (_37556_, _37555_, _37552_);
  and _87830_ (_37558_, _37556_, _07339_);
  or _87831_ (_37559_, _37408_, _08503_);
  and _87832_ (_37560_, _37543_, _06507_);
  and _87833_ (_37561_, _37560_, _37559_);
  or _87834_ (_37562_, _37561_, _37558_);
  and _87835_ (_37563_, _37562_, _07331_);
  and _87836_ (_37564_, _37437_, _06610_);
  and _87837_ (_37565_, _37564_, _37559_);
  or _87838_ (_37566_, _37565_, _06509_);
  or _87839_ (_37567_, _37566_, _37563_);
  and _87840_ (_37569_, _14945_, _08014_);
  or _87841_ (_37570_, _37408_, _09107_);
  or _87842_ (_37571_, _37570_, _37569_);
  and _87843_ (_37572_, _37571_, _09112_);
  and _87844_ (_37573_, _37572_, _37567_);
  nor _87845_ (_37574_, _10608_, _06015_);
  nor _87846_ (_37575_, _10582_, _14239_);
  or _87847_ (_37576_, _37575_, _37408_);
  and _87848_ (_37577_, _37576_, _06602_);
  or _87849_ (_37578_, _37577_, _37574_);
  or _87850_ (_37580_, _37578_, _37573_);
  not _87851_ (_37581_, _37574_);
  nor _87852_ (_37582_, _37479_, _14229_);
  nor _87853_ (_37583_, _37582_, _37478_);
  and _87854_ (_37584_, _37583_, _11154_);
  and _87855_ (_37585_, _37478_, _11151_);
  or _87856_ (_37586_, _37585_, _37584_);
  or _87857_ (_37587_, _37586_, _37581_);
  and _87858_ (_37588_, _37587_, _37580_);
  nor _87859_ (_37589_, _10708_, _06015_);
  or _87860_ (_37590_, _37589_, _37588_);
  not _87861_ (_37591_, _37589_);
  or _87862_ (_37592_, _37591_, _37586_);
  and _87863_ (_37593_, _37592_, _11158_);
  and _87864_ (_37594_, _37593_, _37590_);
  or _87865_ (_37595_, _37416_, _14485_);
  and _87866_ (_37596_, _37595_, _11182_);
  or _87867_ (_37597_, _37596_, _37413_);
  not _87868_ (_37598_, _37413_);
  or _87869_ (_37599_, _37598_, _11179_);
  and _87870_ (_37601_, _37599_, _11129_);
  and _87871_ (_37602_, _37601_, _37597_);
  or _87872_ (_37603_, _37602_, _11188_);
  or _87873_ (_37604_, _37603_, _37594_);
  nor _87874_ (_37605_, _37495_, _14491_);
  nor _87875_ (_37606_, _37605_, _37493_);
  and _87876_ (_37607_, _37606_, _11212_);
  and _87877_ (_37608_, _37493_, _11209_);
  or _87878_ (_37609_, _37608_, _37607_);
  or _87879_ (_37610_, _37609_, _06601_);
  nor _87880_ (_37612_, _37509_, _14497_);
  nor _87881_ (_37613_, _37612_, _37506_);
  and _87882_ (_37614_, _37613_, _11241_);
  and _87883_ (_37615_, _37506_, _11238_);
  or _87884_ (_37616_, _37615_, _37614_);
  or _87885_ (_37617_, _37616_, _11218_);
  and _87886_ (_37618_, _37617_, _11248_);
  and _87887_ (_37619_, _37618_, _37610_);
  and _87888_ (_37620_, _37619_, _37604_);
  or _87889_ (_37621_, _11284_, _10607_);
  nand _87890_ (_37623_, _11284_, _37477_);
  nand _87891_ (_37624_, _37623_, _37621_);
  nor _87892_ (_37625_, _37624_, _11248_);
  or _87893_ (_37626_, _37625_, _17690_);
  or _87894_ (_37627_, _37626_, _37620_);
  and _87895_ (_37628_, _37627_, _37405_);
  or _87896_ (_37629_, _37628_, _07019_);
  or _87897_ (_37630_, _37404_, _07020_);
  and _87898_ (_37631_, _37630_, _13046_);
  and _87899_ (_37632_, _37631_, _37629_);
  or _87900_ (_37634_, _10598_, _09095_);
  and _87901_ (_37635_, _14522_, _37634_);
  nand _87902_ (_37636_, _11368_, _14526_);
  and _87903_ (_37637_, _37636_, _14528_);
  or _87904_ (_37638_, _37637_, _06639_);
  or _87905_ (_37639_, _37638_, _37635_);
  or _87906_ (_37640_, _37639_, _37632_);
  or _87907_ (_37641_, _37433_, _07048_);
  and _87908_ (_37642_, _37641_, _05990_);
  and _87909_ (_37643_, _37642_, _37640_);
  and _87910_ (_37645_, _37427_, _05989_);
  or _87911_ (_37646_, _37645_, _06646_);
  or _87912_ (_37647_, _37646_, _37643_);
  and _87913_ (_37648_, _15129_, _08014_);
  or _87914_ (_37649_, _37408_, _06651_);
  or _87915_ (_37650_, _37649_, _37648_);
  and _87916_ (_37651_, _37650_, _01442_);
  and _87917_ (_37652_, _37651_, _37647_);
  or _87918_ (_37653_, _37652_, _37399_);
  and _87919_ (_44301_, _37653_, _43634_);
  nor _87920_ (_37655_, _01442_, _06419_);
  nor _87921_ (_37656_, _08640_, _06419_);
  and _87922_ (_37657_, _15148_, _08640_);
  or _87923_ (_37658_, _37657_, _37656_);
  and _87924_ (_37659_, _37658_, _06352_);
  nor _87925_ (_37660_, _08014_, _06419_);
  and _87926_ (_37661_, _15153_, _08014_);
  or _87927_ (_37662_, _37661_, _37660_);
  or _87928_ (_37663_, _37662_, _07275_);
  and _87929_ (_37664_, _08014_, \oc8051_golden_model_1.ACC [3]);
  or _87930_ (_37666_, _37664_, _37660_);
  and _87931_ (_37667_, _37666_, _07259_);
  nor _87932_ (_37668_, _07259_, _06419_);
  or _87933_ (_37669_, _37668_, _06474_);
  or _87934_ (_37670_, _37669_, _37667_);
  and _87935_ (_37671_, _37670_, _06357_);
  and _87936_ (_37672_, _37671_, _37663_);
  and _87937_ (_37673_, _15150_, _08640_);
  or _87938_ (_37674_, _37673_, _37656_);
  and _87939_ (_37675_, _37674_, _06356_);
  or _87940_ (_37677_, _37675_, _06410_);
  or _87941_ (_37678_, _37677_, _37672_);
  nor _87942_ (_37679_, _14239_, _07680_);
  or _87943_ (_37680_, _37679_, _37660_);
  or _87944_ (_37681_, _37680_, _06772_);
  and _87945_ (_37682_, _37681_, _37678_);
  or _87946_ (_37683_, _37682_, _06417_);
  or _87947_ (_37684_, _37666_, _06426_);
  and _87948_ (_37685_, _37684_, _06353_);
  and _87949_ (_37686_, _37685_, _37683_);
  or _87950_ (_37688_, _37686_, _37659_);
  and _87951_ (_37689_, _37688_, _06346_);
  and _87952_ (_37690_, _15181_, _08640_);
  or _87953_ (_37691_, _37690_, _37656_);
  and _87954_ (_37692_, _37691_, _06345_);
  or _87955_ (_37693_, _37692_, _37689_);
  and _87956_ (_37694_, _37693_, _06340_);
  and _87957_ (_37695_, _15197_, _08640_);
  or _87958_ (_37696_, _37695_, _37656_);
  and _87959_ (_37697_, _37696_, _06339_);
  or _87960_ (_37699_, _37697_, _10153_);
  or _87961_ (_37700_, _37699_, _37694_);
  or _87962_ (_37701_, _37680_, _06327_);
  and _87963_ (_37702_, _37701_, _06333_);
  and _87964_ (_37703_, _37702_, _37700_);
  and _87965_ (_37704_, _09310_, _08014_);
  or _87966_ (_37705_, _37704_, _37660_);
  and _87967_ (_37706_, _37705_, _09572_);
  or _87968_ (_37707_, _37706_, _06037_);
  or _87969_ (_37708_, _37707_, _37703_);
  and _87970_ (_37710_, _15251_, _08014_);
  or _87971_ (_37711_, _37660_, _06313_);
  or _87972_ (_37712_, _37711_, _37710_);
  and _87973_ (_37713_, _37712_, _06278_);
  and _87974_ (_37714_, _37713_, _37708_);
  and _87975_ (_37715_, _08014_, _09014_);
  or _87976_ (_37716_, _37715_, _37660_);
  and _87977_ (_37717_, _37716_, _06277_);
  or _87978_ (_37718_, _37717_, _06502_);
  or _87979_ (_37719_, _37718_, _37714_);
  and _87980_ (_37721_, _15266_, _08014_);
  or _87981_ (_37722_, _37660_, _07334_);
  or _87982_ (_37723_, _37722_, _37721_);
  and _87983_ (_37724_, _37723_, _07337_);
  and _87984_ (_37725_, _37724_, _37719_);
  and _87985_ (_37726_, _12619_, _08014_);
  or _87986_ (_37727_, _37726_, _37660_);
  and _87987_ (_37728_, _37727_, _06615_);
  or _87988_ (_37729_, _37728_, _37725_);
  and _87989_ (_37730_, _37729_, _07339_);
  or _87990_ (_37732_, _37660_, _08359_);
  and _87991_ (_37733_, _37716_, _06507_);
  and _87992_ (_37734_, _37733_, _37732_);
  or _87993_ (_37735_, _37734_, _37730_);
  and _87994_ (_37736_, _37735_, _07331_);
  and _87995_ (_37737_, _37666_, _06610_);
  and _87996_ (_37738_, _37737_, _37732_);
  or _87997_ (_37739_, _37738_, _06509_);
  or _87998_ (_37740_, _37739_, _37736_);
  and _87999_ (_37741_, _15263_, _08014_);
  or _88000_ (_37743_, _37660_, _09107_);
  or _88001_ (_37744_, _37743_, _37741_);
  and _88002_ (_37745_, _37744_, _09112_);
  and _88003_ (_37746_, _37745_, _37740_);
  nor _88004_ (_37747_, _10574_, _14239_);
  or _88005_ (_37748_, _37747_, _37660_);
  and _88006_ (_37749_, _37748_, _06602_);
  or _88007_ (_37750_, _37749_, _06639_);
  or _88008_ (_37751_, _37750_, _37746_);
  or _88009_ (_37752_, _37662_, _07048_);
  and _88010_ (_37754_, _37752_, _05990_);
  and _88011_ (_37755_, _37754_, _37751_);
  and _88012_ (_37756_, _37658_, _05989_);
  or _88013_ (_37757_, _37756_, _06646_);
  or _88014_ (_37758_, _37757_, _37755_);
  and _88015_ (_37759_, _15321_, _08014_);
  or _88016_ (_37760_, _37660_, _06651_);
  or _88017_ (_37761_, _37760_, _37759_);
  and _88018_ (_37762_, _37761_, _01442_);
  and _88019_ (_37763_, _37762_, _37758_);
  or _88020_ (_37765_, _37763_, _37655_);
  and _88021_ (_44302_, _37765_, _43634_);
  and _88022_ (_37766_, _01446_, \oc8051_golden_model_1.PSW [4]);
  and _88023_ (_37767_, _14239_, \oc8051_golden_model_1.PSW [4]);
  nor _88024_ (_37768_, _10589_, _14239_);
  or _88025_ (_37769_, _37768_, _37767_);
  and _88026_ (_37770_, _08014_, \oc8051_golden_model_1.ACC [4]);
  nand _88027_ (_37771_, _37770_, _08599_);
  and _88028_ (_37772_, _37771_, _06615_);
  and _88029_ (_37773_, _37772_, _37769_);
  and _88030_ (_37775_, _15367_, _08014_);
  or _88031_ (_37776_, _37775_, _37767_);
  or _88032_ (_37777_, _37776_, _07275_);
  or _88033_ (_37778_, _37770_, _37767_);
  and _88034_ (_37779_, _37778_, _07259_);
  and _88035_ (_37780_, _07260_, \oc8051_golden_model_1.PSW [4]);
  or _88036_ (_37781_, _37780_, _06474_);
  or _88037_ (_37782_, _37781_, _37779_);
  and _88038_ (_37783_, _37782_, _06357_);
  and _88039_ (_37784_, _37783_, _37777_);
  and _88040_ (_37786_, _37211_, \oc8051_golden_model_1.PSW [4]);
  and _88041_ (_37787_, _15353_, _08640_);
  or _88042_ (_37788_, _37787_, _37786_);
  and _88043_ (_37789_, _37788_, _06356_);
  or _88044_ (_37790_, _37789_, _06410_);
  or _88045_ (_37791_, _37790_, _37784_);
  nor _88046_ (_37792_, _08596_, _14239_);
  or _88047_ (_37793_, _37792_, _37767_);
  or _88048_ (_37794_, _37793_, _06772_);
  and _88049_ (_37795_, _37794_, _37791_);
  or _88050_ (_37797_, _37795_, _06417_);
  or _88051_ (_37798_, _37778_, _06426_);
  and _88052_ (_37799_, _37798_, _06353_);
  and _88053_ (_37800_, _37799_, _37797_);
  and _88054_ (_37801_, _15348_, _08640_);
  or _88055_ (_37802_, _37801_, _37786_);
  and _88056_ (_37803_, _37802_, _06352_);
  or _88057_ (_37804_, _37803_, _06345_);
  or _88058_ (_37805_, _37804_, _37800_);
  or _88059_ (_37806_, _37786_, _15384_);
  and _88060_ (_37808_, _37806_, _37788_);
  or _88061_ (_37809_, _37808_, _06346_);
  and _88062_ (_37810_, _37809_, _06340_);
  and _88063_ (_37811_, _37810_, _37805_);
  and _88064_ (_37812_, _15350_, _08640_);
  or _88065_ (_37813_, _37812_, _37786_);
  and _88066_ (_37814_, _37813_, _06339_);
  or _88067_ (_37815_, _37814_, _10153_);
  or _88068_ (_37816_, _37815_, _37811_);
  or _88069_ (_37817_, _37793_, _06327_);
  and _88070_ (_37819_, _37817_, _06333_);
  and _88071_ (_37820_, _37819_, _37816_);
  and _88072_ (_37821_, _09264_, _08014_);
  or _88073_ (_37822_, _37821_, _37767_);
  and _88074_ (_37823_, _37822_, _09572_);
  or _88075_ (_37824_, _37823_, _06037_);
  or _88076_ (_37825_, _37824_, _37820_);
  and _88077_ (_37826_, _15452_, _08014_);
  or _88078_ (_37827_, _37767_, _06313_);
  or _88079_ (_37828_, _37827_, _37826_);
  and _88080_ (_37830_, _37828_, _06278_);
  and _88081_ (_37831_, _37830_, _37825_);
  and _88082_ (_37832_, _08995_, _08014_);
  or _88083_ (_37833_, _37832_, _37767_);
  and _88084_ (_37834_, _37833_, _06277_);
  or _88085_ (_37835_, _37834_, _06502_);
  or _88086_ (_37836_, _37835_, _37831_);
  and _88087_ (_37837_, _15345_, _08014_);
  or _88088_ (_37838_, _37767_, _07334_);
  or _88089_ (_37839_, _37838_, _37837_);
  and _88090_ (_37841_, _37839_, _07337_);
  and _88091_ (_37842_, _37841_, _37836_);
  or _88092_ (_37843_, _37842_, _37773_);
  and _88093_ (_37844_, _37843_, _07339_);
  or _88094_ (_37845_, _37767_, _08599_);
  and _88095_ (_37846_, _37833_, _06507_);
  and _88096_ (_37847_, _37846_, _37845_);
  or _88097_ (_37848_, _37847_, _37844_);
  and _88098_ (_37849_, _37848_, _07331_);
  and _88099_ (_37850_, _37778_, _06610_);
  and _88100_ (_37852_, _37850_, _37845_);
  or _88101_ (_37853_, _37852_, _06509_);
  or _88102_ (_37854_, _37853_, _37849_);
  and _88103_ (_37855_, _15342_, _08014_);
  or _88104_ (_37856_, _37767_, _09107_);
  or _88105_ (_37857_, _37856_, _37855_);
  and _88106_ (_37858_, _37857_, _09112_);
  and _88107_ (_37859_, _37858_, _37854_);
  and _88108_ (_37860_, _37769_, _06602_);
  or _88109_ (_37861_, _37860_, _06639_);
  or _88110_ (_37863_, _37861_, _37859_);
  or _88111_ (_37864_, _37776_, _07048_);
  and _88112_ (_37865_, _37864_, _05990_);
  and _88113_ (_37866_, _37865_, _37863_);
  and _88114_ (_37867_, _37802_, _05989_);
  or _88115_ (_37868_, _37867_, _06646_);
  or _88116_ (_37869_, _37868_, _37866_);
  and _88117_ (_37870_, _15524_, _08014_);
  or _88118_ (_37871_, _37767_, _06651_);
  or _88119_ (_37872_, _37871_, _37870_);
  and _88120_ (_37874_, _37872_, _01442_);
  and _88121_ (_37875_, _37874_, _37869_);
  or _88122_ (_37876_, _37875_, _37766_);
  and _88123_ (_44303_, _37876_, _43634_);
  and _88124_ (_37877_, _01446_, \oc8051_golden_model_1.PSW [5]);
  and _88125_ (_37878_, _14239_, \oc8051_golden_model_1.PSW [5]);
  and _88126_ (_37879_, _15550_, _08014_);
  or _88127_ (_37880_, _37879_, _37878_);
  or _88128_ (_37881_, _37880_, _07275_);
  and _88129_ (_37882_, _08014_, \oc8051_golden_model_1.ACC [5]);
  or _88130_ (_37884_, _37882_, _37878_);
  and _88131_ (_37885_, _37884_, _07259_);
  and _88132_ (_37886_, _07260_, \oc8051_golden_model_1.PSW [5]);
  or _88133_ (_37887_, _37886_, _06474_);
  or _88134_ (_37888_, _37887_, _37885_);
  and _88135_ (_37889_, _37888_, _06357_);
  and _88136_ (_37890_, _37889_, _37881_);
  and _88137_ (_37891_, _37211_, \oc8051_golden_model_1.PSW [5]);
  and _88138_ (_37892_, _15566_, _08640_);
  or _88139_ (_37893_, _37892_, _37891_);
  and _88140_ (_37895_, _37893_, _06356_);
  or _88141_ (_37896_, _37895_, _06410_);
  or _88142_ (_37897_, _37896_, _37890_);
  nor _88143_ (_37898_, _08305_, _14239_);
  or _88144_ (_37899_, _37898_, _37878_);
  or _88145_ (_37900_, _37899_, _06772_);
  and _88146_ (_37901_, _37900_, _37897_);
  or _88147_ (_37902_, _37901_, _06417_);
  or _88148_ (_37903_, _37884_, _06426_);
  and _88149_ (_37904_, _37903_, _06353_);
  and _88150_ (_37906_, _37904_, _37902_);
  and _88151_ (_37907_, _15544_, _08640_);
  or _88152_ (_37908_, _37907_, _37891_);
  and _88153_ (_37909_, _37908_, _06352_);
  or _88154_ (_37910_, _37909_, _06345_);
  or _88155_ (_37911_, _37910_, _37906_);
  or _88156_ (_37912_, _37891_, _15581_);
  and _88157_ (_37913_, _37912_, _37893_);
  or _88158_ (_37914_, _37913_, _06346_);
  and _88159_ (_37915_, _37914_, _06340_);
  and _88160_ (_37917_, _37915_, _37911_);
  and _88161_ (_37918_, _15546_, _08640_);
  or _88162_ (_37919_, _37918_, _37891_);
  and _88163_ (_37920_, _37919_, _06339_);
  or _88164_ (_37921_, _37920_, _10153_);
  or _88165_ (_37922_, _37921_, _37917_);
  or _88166_ (_37923_, _37899_, _06327_);
  and _88167_ (_37924_, _37923_, _06333_);
  and _88168_ (_37925_, _37924_, _37922_);
  and _88169_ (_37926_, _09218_, _08014_);
  or _88170_ (_37928_, _37926_, _37878_);
  and _88171_ (_37929_, _37928_, _09572_);
  or _88172_ (_37930_, _37929_, _06037_);
  or _88173_ (_37931_, _37930_, _37925_);
  and _88174_ (_37932_, _15649_, _08014_);
  or _88175_ (_37933_, _37878_, _06313_);
  or _88176_ (_37934_, _37933_, _37932_);
  and _88177_ (_37935_, _37934_, _06278_);
  and _88178_ (_37936_, _37935_, _37931_);
  and _88179_ (_37937_, _08954_, _08014_);
  or _88180_ (_37939_, _37937_, _37878_);
  and _88181_ (_37940_, _37939_, _06277_);
  or _88182_ (_37941_, _37940_, _06502_);
  or _88183_ (_37942_, _37941_, _37936_);
  and _88184_ (_37943_, _15664_, _08014_);
  or _88185_ (_37944_, _37878_, _07334_);
  or _88186_ (_37945_, _37944_, _37943_);
  and _88187_ (_37946_, _37945_, _07337_);
  and _88188_ (_37947_, _37946_, _37942_);
  and _88189_ (_37948_, _12626_, _08014_);
  or _88190_ (_37950_, _37948_, _37878_);
  and _88191_ (_37951_, _37950_, _06615_);
  or _88192_ (_37952_, _37951_, _37947_);
  and _88193_ (_37953_, _37952_, _07339_);
  or _88194_ (_37954_, _37878_, _08308_);
  and _88195_ (_37955_, _37939_, _06507_);
  and _88196_ (_37956_, _37955_, _37954_);
  or _88197_ (_37957_, _37956_, _37953_);
  and _88198_ (_37958_, _37957_, _07331_);
  and _88199_ (_37959_, _37884_, _06610_);
  and _88200_ (_37961_, _37959_, _37954_);
  or _88201_ (_37962_, _37961_, _06509_);
  or _88202_ (_37963_, _37962_, _37958_);
  and _88203_ (_37964_, _15663_, _08014_);
  or _88204_ (_37965_, _37878_, _09107_);
  or _88205_ (_37966_, _37965_, _37964_);
  and _88206_ (_37967_, _37966_, _09112_);
  and _88207_ (_37968_, _37967_, _37963_);
  nor _88208_ (_37969_, _10570_, _14239_);
  or _88209_ (_37970_, _37969_, _37878_);
  and _88210_ (_37972_, _37970_, _06602_);
  or _88211_ (_37973_, _37972_, _06639_);
  or _88212_ (_37974_, _37973_, _37968_);
  or _88213_ (_37975_, _37880_, _07048_);
  and _88214_ (_37976_, _37975_, _05990_);
  and _88215_ (_37977_, _37976_, _37974_);
  and _88216_ (_37978_, _37908_, _05989_);
  or _88217_ (_37979_, _37978_, _06646_);
  or _88218_ (_37980_, _37979_, _37977_);
  and _88219_ (_37981_, _15721_, _08014_);
  or _88220_ (_37983_, _37878_, _06651_);
  or _88221_ (_37984_, _37983_, _37981_);
  and _88222_ (_37985_, _37984_, _01442_);
  and _88223_ (_37986_, _37985_, _37980_);
  or _88224_ (_37987_, _37986_, _37877_);
  and _88225_ (_44305_, _37987_, _43634_);
  nor _88226_ (_37988_, _01442_, _18384_);
  or _88227_ (_37989_, _11232_, _10927_);
  and _88228_ (_37990_, _37989_, _11186_);
  nor _88229_ (_37991_, _08014_, _18384_);
  nor _88230_ (_37993_, _08209_, _14239_);
  or _88231_ (_37994_, _37993_, _37991_);
  or _88232_ (_37995_, _37994_, _06327_);
  nor _88233_ (_37996_, _08640_, _18384_);
  and _88234_ (_37997_, _15763_, _08640_);
  or _88235_ (_37998_, _37997_, _37996_);
  or _88236_ (_37999_, _37996_, _15778_);
  and _88237_ (_38000_, _37999_, _37998_);
  or _88238_ (_38001_, _38000_, _06346_);
  and _88239_ (_38002_, _15759_, _08014_);
  or _88240_ (_38004_, _38002_, _37991_);
  or _88241_ (_38005_, _38004_, _07275_);
  and _88242_ (_38006_, _08014_, \oc8051_golden_model_1.ACC [6]);
  or _88243_ (_38007_, _38006_, _37991_);
  and _88244_ (_38008_, _38007_, _07259_);
  nor _88245_ (_38009_, _07259_, _18384_);
  or _88246_ (_38010_, _38009_, _06474_);
  or _88247_ (_38011_, _38010_, _38008_);
  and _88248_ (_38012_, _38011_, _06357_);
  and _88249_ (_38013_, _38012_, _38005_);
  and _88250_ (_38015_, _37998_, _06356_);
  or _88251_ (_38016_, _38015_, _06410_);
  or _88252_ (_38017_, _38016_, _38013_);
  or _88253_ (_38018_, _37994_, _06772_);
  and _88254_ (_38019_, _38018_, _38017_);
  or _88255_ (_38020_, _38019_, _06417_);
  or _88256_ (_38021_, _38007_, _06426_);
  and _88257_ (_38022_, _38021_, _06353_);
  and _88258_ (_38023_, _38022_, _38020_);
  and _88259_ (_38024_, _15743_, _08640_);
  or _88260_ (_38026_, _38024_, _37996_);
  and _88261_ (_38027_, _38026_, _06352_);
  or _88262_ (_38028_, _38027_, _06345_);
  or _88263_ (_38029_, _38028_, _38023_);
  and _88264_ (_38030_, _38029_, _38001_);
  and _88265_ (_38031_, _38030_, _10784_);
  or _88266_ (_38032_, _10853_, _10790_);
  or _88267_ (_38033_, _38032_, _10841_);
  and _88268_ (_38034_, _38033_, _12671_);
  or _88269_ (_38035_, _38034_, _38031_);
  or _88270_ (_38037_, _10876_, _10854_);
  or _88271_ (_38038_, _38037_, _10909_);
  and _88272_ (_38039_, _38038_, _38035_);
  or _88273_ (_38040_, _38039_, _12337_);
  or _88274_ (_38041_, _10633_, _06458_);
  or _88275_ (_38042_, _38041_, _10679_);
  or _88276_ (_38043_, _10927_, _10624_);
  or _88277_ (_38044_, _38043_, _10986_);
  and _88278_ (_38045_, _38044_, _06340_);
  and _88279_ (_38046_, _38045_, _38042_);
  and _88280_ (_38048_, _38046_, _38040_);
  and _88281_ (_38049_, _15745_, _08640_);
  or _88282_ (_38050_, _38049_, _37996_);
  and _88283_ (_38051_, _38050_, _06339_);
  or _88284_ (_38052_, _38051_, _10153_);
  or _88285_ (_38053_, _38052_, _38048_);
  and _88286_ (_38054_, _38053_, _37995_);
  or _88287_ (_38055_, _38054_, _09572_);
  and _88288_ (_38056_, _09172_, _08014_);
  or _88289_ (_38057_, _37991_, _06333_);
  or _88290_ (_38059_, _38057_, _38056_);
  and _88291_ (_38060_, _38059_, _06313_);
  and _88292_ (_38061_, _38060_, _38055_);
  and _88293_ (_38062_, _15846_, _08014_);
  or _88294_ (_38063_, _38062_, _37991_);
  and _88295_ (_38064_, _38063_, _06037_);
  or _88296_ (_38065_, _38064_, _06277_);
  or _88297_ (_38066_, _38065_, _38061_);
  and _88298_ (_38067_, _15853_, _08014_);
  or _88299_ (_38068_, _38067_, _37991_);
  or _88300_ (_38070_, _38068_, _06278_);
  and _88301_ (_38071_, _38070_, _38066_);
  or _88302_ (_38072_, _38071_, _06502_);
  and _88303_ (_38073_, _15862_, _08014_);
  or _88304_ (_38074_, _37991_, _07334_);
  or _88305_ (_38075_, _38074_, _38073_);
  and _88306_ (_38076_, _38075_, _07337_);
  and _88307_ (_38077_, _38076_, _38072_);
  and _88308_ (_38078_, _10596_, _08014_);
  or _88309_ (_38079_, _38078_, _37991_);
  and _88310_ (_38081_, _38079_, _06615_);
  or _88311_ (_38082_, _38081_, _38077_);
  and _88312_ (_38083_, _38082_, _07339_);
  or _88313_ (_38084_, _37991_, _08212_);
  and _88314_ (_38085_, _38068_, _06507_);
  and _88315_ (_38086_, _38085_, _38084_);
  or _88316_ (_38087_, _38086_, _38083_);
  and _88317_ (_38088_, _38087_, _07331_);
  and _88318_ (_38089_, _38007_, _06610_);
  and _88319_ (_38090_, _38089_, _38084_);
  or _88320_ (_38092_, _38090_, _06509_);
  or _88321_ (_38093_, _38092_, _38088_);
  and _88322_ (_38094_, _15859_, _08014_);
  or _88323_ (_38095_, _38094_, _37991_);
  or _88324_ (_38096_, _38095_, _09107_);
  and _88325_ (_38097_, _38096_, _38093_);
  or _88326_ (_38098_, _38097_, _06602_);
  nor _88327_ (_38099_, _10595_, _14239_);
  or _88328_ (_38100_, _38099_, _37991_);
  or _88329_ (_38101_, _38100_, _09112_);
  and _88330_ (_38103_, _38101_, _11123_);
  and _88331_ (_38104_, _38103_, _38098_);
  or _88332_ (_38105_, _11145_, _10790_);
  and _88333_ (_38106_, _38105_, _11122_);
  or _88334_ (_38107_, _38106_, _06995_);
  or _88335_ (_38108_, _38107_, _38104_);
  nor _88336_ (_38109_, _38105_, _06996_);
  and _88337_ (_38110_, _06323_, _06511_);
  nor _88338_ (_38111_, _38110_, _38109_);
  and _88339_ (_38112_, _38111_, _38108_);
  and _88340_ (_38114_, _38110_, _38105_);
  or _88341_ (_38115_, _38114_, _11124_);
  or _88342_ (_38116_, _38115_, _38112_);
  not _88343_ (_38117_, _11124_);
  or _88344_ (_38118_, _38105_, _38117_);
  and _88345_ (_38119_, _38118_, _18231_);
  and _88346_ (_38120_, _38119_, _38116_);
  or _88347_ (_38121_, _11173_, _10876_);
  and _88348_ (_38122_, _38121_, _17922_);
  or _88349_ (_38123_, _38122_, _38120_);
  and _88350_ (_38125_, _38123_, _18237_);
  and _88351_ (_38126_, _38121_, _07002_);
  or _88352_ (_38127_, _38126_, _06600_);
  or _88353_ (_38128_, _38127_, _38125_);
  or _88354_ (_38129_, _10633_, _06601_);
  or _88355_ (_38130_, _38129_, _11203_);
  and _88356_ (_38131_, _38130_, _11218_);
  and _88357_ (_38132_, _38131_, _38128_);
  or _88358_ (_38133_, _38132_, _37990_);
  and _88359_ (_38134_, _38133_, _11248_);
  and _88360_ (_38136_, _11277_, _18254_);
  or _88361_ (_38137_, _38136_, _11290_);
  or _88362_ (_38138_, _38137_, _38134_);
  or _88363_ (_38139_, _11320_, _11292_);
  and _88364_ (_38140_, _38139_, _06364_);
  and _88365_ (_38141_, _38140_, _38138_);
  and _88366_ (_38142_, _10588_, _06363_);
  or _88367_ (_38143_, _38142_, _10566_);
  or _88368_ (_38144_, _38143_, _38141_);
  or _88369_ (_38145_, _11362_, _10567_);
  and _88370_ (_38147_, _38145_, _38144_);
  or _88371_ (_38148_, _38147_, _06639_);
  or _88372_ (_38149_, _38004_, _07048_);
  and _88373_ (_38150_, _38149_, _05990_);
  and _88374_ (_38151_, _38150_, _38148_);
  and _88375_ (_38152_, _38026_, _05989_);
  or _88376_ (_38153_, _38152_, _06646_);
  or _88377_ (_38154_, _38153_, _38151_);
  and _88378_ (_38155_, _15921_, _08014_);
  or _88379_ (_38156_, _37991_, _06651_);
  or _88380_ (_38158_, _38156_, _38155_);
  and _88381_ (_38159_, _38158_, _01442_);
  and _88382_ (_38160_, _38159_, _38154_);
  or _88383_ (_38161_, _38160_, _37988_);
  and _88384_ (_44306_, _38161_, _43634_);
  or _88385_ (_38162_, _00000_, \oc8051_golden_model_1.P0INREG [0]);
  or _88386_ (_38163_, _07543_, p0_in[0]);
  and _88387_ (_44307_, _38163_, _38162_);
  or _88388_ (_38164_, _00000_, \oc8051_golden_model_1.P0INREG [1]);
  or _88389_ (_38165_, _07543_, p0_in[1]);
  and _88390_ (_44309_, _38165_, _38164_);
  or _88391_ (_38167_, _00000_, \oc8051_golden_model_1.P0INREG [2]);
  or _88392_ (_38168_, _07543_, p0_in[2]);
  and _88393_ (_44310_, _38168_, _38167_);
  or _88394_ (_38169_, _00000_, \oc8051_golden_model_1.P0INREG [3]);
  or _88395_ (_38170_, _07543_, p0_in[3]);
  and _88396_ (_44311_, _38170_, _38169_);
  or _88397_ (_38171_, _00000_, \oc8051_golden_model_1.P0INREG [4]);
  or _88398_ (_38172_, _07543_, p0_in[4]);
  and _88399_ (_44312_, _38172_, _38171_);
  or _88400_ (_38174_, _00000_, \oc8051_golden_model_1.P0INREG [5]);
  or _88401_ (_38175_, _07543_, p0_in[5]);
  and _88402_ (_44313_, _38175_, _38174_);
  or _88403_ (_38176_, _00000_, \oc8051_golden_model_1.P0INREG [6]);
  or _88404_ (_38177_, _07543_, p0_in[6]);
  and _88405_ (_44314_, _38177_, _38176_);
  or _88406_ (_38178_, _00000_, \oc8051_golden_model_1.P1INREG [0]);
  or _88407_ (_38179_, _07543_, p1_in[0]);
  and _88408_ (_44316_, _38179_, _38178_);
  or _88409_ (_38180_, _00000_, \oc8051_golden_model_1.P1INREG [1]);
  or _88410_ (_38182_, _07543_, p1_in[1]);
  and _88411_ (_44317_, _38182_, _38180_);
  or _88412_ (_38183_, _00000_, \oc8051_golden_model_1.P1INREG [2]);
  or _88413_ (_38184_, _07543_, p1_in[2]);
  and _88414_ (_44318_, _38184_, _38183_);
  or _88415_ (_38185_, _00000_, \oc8051_golden_model_1.P1INREG [3]);
  or _88416_ (_38186_, _07543_, p1_in[3]);
  and _88417_ (_44319_, _38186_, _38185_);
  or _88418_ (_38187_, _00000_, \oc8051_golden_model_1.P1INREG [4]);
  or _88419_ (_38188_, _07543_, p1_in[4]);
  and _88420_ (_44320_, _38188_, _38187_);
  or _88421_ (_38190_, _00000_, \oc8051_golden_model_1.P1INREG [5]);
  or _88422_ (_38191_, _07543_, p1_in[5]);
  and _88423_ (_44321_, _38191_, _38190_);
  or _88424_ (_38192_, _00000_, \oc8051_golden_model_1.P1INREG [6]);
  or _88425_ (_38193_, _07543_, p1_in[6]);
  and _88426_ (_44322_, _38193_, _38192_);
  or _88427_ (_38194_, _00000_, \oc8051_golden_model_1.P2INREG [0]);
  or _88428_ (_38195_, _07543_, p2_in[0]);
  and _88429_ (_44324_, _38195_, _38194_);
  or _88430_ (_38197_, _00000_, \oc8051_golden_model_1.P2INREG [1]);
  or _88431_ (_38198_, _07543_, p2_in[1]);
  and _88432_ (_44325_, _38198_, _38197_);
  or _88433_ (_38199_, _00000_, \oc8051_golden_model_1.P2INREG [2]);
  or _88434_ (_38200_, _07543_, p2_in[2]);
  and _88435_ (_44326_, _38200_, _38199_);
  or _88436_ (_38201_, _00000_, \oc8051_golden_model_1.P2INREG [3]);
  or _88437_ (_38202_, _07543_, p2_in[3]);
  and _88438_ (_44328_, _38202_, _38201_);
  or _88439_ (_38203_, _00000_, \oc8051_golden_model_1.P2INREG [4]);
  or _88440_ (_38205_, _07543_, p2_in[4]);
  and _88441_ (_44329_, _38205_, _38203_);
  or _88442_ (_38206_, _00000_, \oc8051_golden_model_1.P2INREG [5]);
  or _88443_ (_38207_, _07543_, p2_in[5]);
  and _88444_ (_44330_, _38207_, _38206_);
  or _88445_ (_38208_, _00000_, \oc8051_golden_model_1.P2INREG [6]);
  or _88446_ (_38209_, _07543_, p2_in[6]);
  and _88447_ (_44331_, _38209_, _38208_);
  or _88448_ (_38210_, _00000_, \oc8051_golden_model_1.P3INREG [0]);
  or _88449_ (_38211_, _07543_, p3_in[0]);
  and _88450_ (_44333_, _38211_, _38210_);
  or _88451_ (_38213_, _00000_, \oc8051_golden_model_1.P3INREG [1]);
  or _88452_ (_38214_, _07543_, p3_in[1]);
  and _88453_ (_44334_, _38214_, _38213_);
  or _88454_ (_38215_, _00000_, \oc8051_golden_model_1.P3INREG [2]);
  or _88455_ (_38216_, _07543_, p3_in[2]);
  and _88456_ (_44335_, _38216_, _38215_);
  or _88457_ (_38217_, _00000_, \oc8051_golden_model_1.P3INREG [3]);
  or _88458_ (_38218_, _07543_, p3_in[3]);
  and _88459_ (_44336_, _38218_, _38217_);
  or _88460_ (_38220_, _00000_, \oc8051_golden_model_1.P3INREG [4]);
  or _88461_ (_38221_, _07543_, p3_in[4]);
  and _88462_ (_44337_, _38221_, _38220_);
  or _88463_ (_38222_, _00000_, \oc8051_golden_model_1.P3INREG [5]);
  or _88464_ (_38223_, _07543_, p3_in[5]);
  and _88465_ (_44338_, _38223_, _38222_);
  or _88466_ (_38224_, _00000_, \oc8051_golden_model_1.P3INREG [6]);
  or _88467_ (_38225_, _07543_, p3_in[6]);
  and _88468_ (_44339_, _38225_, _38224_);
  and _88469_ (_00005_[6], _03678_, _43634_);
  and _88470_ (_00005_[5], _03645_, _43634_);
  and _88471_ (_00005_[4], _03669_, _43634_);
  and _88472_ (_00005_[3], _03629_, _43634_);
  and _88473_ (_00005_[2], _03685_, _43634_);
  and _88474_ (_00005_[1], _03652_, _43634_);
  and _88475_ (_00005_[0], _03662_, _43634_);
  and _88476_ (_00004_[6], _03769_, _43634_);
  and _88477_ (_00004_[5], _03802_, _43634_);
  and _88478_ (_00004_[4], _03793_, _43634_);
  and _88479_ (_00004_[3], _03753_, _43634_);
  and _88480_ (_00004_[2], _03776_, _43634_);
  and _88481_ (_00004_[1], _03809_, _43634_);
  and _88482_ (_00004_[0], _03786_, _43634_);
  and _88483_ (_00003_[6], _03545_, _43634_);
  and _88484_ (_00003_[5], _03522_, _43634_);
  and _88485_ (_00003_[4], _03496_, _43634_);
  and _88486_ (_00003_[3], _03505_, _43634_);
  and _88487_ (_00003_[2], _03538_, _43634_);
  and _88488_ (_00003_[1], _03529_, _43634_);
  and _88489_ (_00003_[0], _03488_, _43634_);
  and _88490_ (_00002_[6], _03615_, _43634_);
  and _88491_ (_00002_[5], _03592_, _43634_);
  and _88492_ (_00002_[4], _03566_, _43634_);
  and _88493_ (_00002_[3], _03575_, _43634_);
  and _88494_ (_00002_[2], _03608_, _43634_);
  and _88495_ (_00002_[1], _03599_, _43634_);
  and _88496_ (_00002_[0], _03559_, _43634_);
  or _88497_ (_38229_, _05996_, _05989_);
  and _88498_ (_38230_, _38229_, op0_cnst);
  or _88499_ (_00001_, _38230_, rst);
  and _88500_ (_00005_[7], _03636_, _43634_);
  and _88501_ (_00004_[7], _03760_, _43634_);
  and _88502_ (_00003_[7], _03512_, _43634_);
  and _88503_ (_00002_[7], _03582_, _43634_);
  and _88504_ (_38232_, inst_finished_r, op0_cnst);
  not _88505_ (_38233_, word_in[1]);
  and _88506_ (_38234_, _38233_, word_in[0]);
  and _88507_ (_38235_, _38234_, \oc8051_golden_model_1.IRAM[1] [0]);
  nor _88508_ (_38236_, _38233_, word_in[0]);
  and _88509_ (_38237_, _38236_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor _88510_ (_38239_, _38237_, _38235_);
  nor _88511_ (_38240_, word_in[1], word_in[0]);
  and _88512_ (_38241_, _38240_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _88513_ (_38242_, word_in[1], word_in[0]);
  and _88514_ (_38243_, _38242_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor _88515_ (_38244_, _38243_, _38241_);
  and _88516_ (_38245_, _38244_, _38239_);
  nor _88517_ (_38246_, word_in[3], word_in[2]);
  not _88518_ (_38247_, _38246_);
  nor _88519_ (_38248_, _38247_, _38245_);
  and _88520_ (_38250_, _38234_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _88521_ (_38251_, _38236_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor _88522_ (_38252_, _38251_, _38250_);
  and _88523_ (_38253_, _38240_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _88524_ (_38254_, _38242_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor _88525_ (_38255_, _38254_, _38253_);
  and _88526_ (_38256_, _38255_, _38252_);
  and _88527_ (_38257_, word_in[3], word_in[2]);
  not _88528_ (_38258_, _38257_);
  nor _88529_ (_38259_, _38258_, _38256_);
  nor _88530_ (_38261_, _38259_, _38248_);
  and _88531_ (_38262_, _38234_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _88532_ (_38263_, _38236_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor _88533_ (_38264_, _38263_, _38262_);
  and _88534_ (_38265_, _38240_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _88535_ (_38266_, _38242_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor _88536_ (_38267_, _38266_, _38265_);
  and _88537_ (_38268_, _38267_, _38264_);
  not _88538_ (_38269_, word_in[3]);
  and _88539_ (_38270_, _38269_, word_in[2]);
  not _88540_ (_38272_, _38270_);
  nor _88541_ (_38273_, _38272_, _38268_);
  and _88542_ (_38274_, _38234_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _88543_ (_38275_, _38236_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor _88544_ (_38276_, _38275_, _38274_);
  and _88545_ (_38277_, _38240_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _88546_ (_38278_, _38242_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor _88547_ (_38279_, _38278_, _38277_);
  and _88548_ (_38280_, _38279_, _38276_);
  nor _88549_ (_38281_, _38269_, word_in[2]);
  not _88550_ (_38283_, _38281_);
  nor _88551_ (_38284_, _38283_, _38280_);
  nor _88552_ (_38285_, _38284_, _38273_);
  and _88553_ (_38286_, _38285_, _38261_);
  and _88554_ (_38287_, _38281_, _38234_);
  and _88555_ (_38288_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _88556_ (_38289_, _38270_, _38234_);
  and _88557_ (_38290_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _88558_ (_38291_, _38290_, _38288_);
  and _88559_ (_38292_, _38257_, _38242_);
  and _88560_ (_38294_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _88561_ (_38295_, _38270_, _38242_);
  and _88562_ (_38296_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _88563_ (_38297_, _38296_, _38294_);
  and _88564_ (_38298_, _38297_, _38291_);
  and _88565_ (_38299_, _38281_, _38240_);
  and _88566_ (_38300_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and _88567_ (_38301_, _38270_, _38240_);
  and _88568_ (_38302_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _88569_ (_38303_, _38302_, _38300_);
  and _88570_ (_38305_, _38246_, _38240_);
  and _88571_ (_38306_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _88572_ (_38307_, _38246_, _38234_);
  and _88573_ (_38308_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _88574_ (_38309_, _38308_, _38306_);
  and _88575_ (_38310_, _38309_, _38303_);
  and _88576_ (_38311_, _38310_, _38298_);
  and _88577_ (_38312_, _38257_, _38234_);
  and _88578_ (_38313_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _88579_ (_38314_, _38281_, _38236_);
  and _88580_ (_38316_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _88581_ (_38317_, _38316_, _38313_);
  and _88582_ (_38318_, _38270_, _38236_);
  and _88583_ (_38319_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _88584_ (_38320_, _38246_, _38236_);
  and _88585_ (_38321_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _88586_ (_38322_, _38321_, _38319_);
  and _88587_ (_38323_, _38322_, _38317_);
  and _88588_ (_38324_, _38257_, _38236_);
  and _88589_ (_38325_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _88590_ (_38327_, _38281_, _38242_);
  and _88591_ (_38328_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _88592_ (_38329_, _38328_, _38325_);
  and _88593_ (_38330_, _38257_, _38240_);
  and _88594_ (_38331_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and _88595_ (_38332_, _38246_, _38242_);
  and _88596_ (_38333_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _88597_ (_38334_, _38333_, _38331_);
  and _88598_ (_38335_, _38334_, _38329_);
  and _88599_ (_38336_, _38335_, _38323_);
  and _88600_ (_38338_, _38336_, _38311_);
  or _88601_ (_38339_, _38338_, _38286_);
  nand _88602_ (_38340_, _38338_, _38286_);
  and _88603_ (_38341_, _38340_, _38339_);
  and _88604_ (_38342_, _38234_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _88605_ (_38343_, _38236_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor _88606_ (_38344_, _38343_, _38342_);
  and _88607_ (_38345_, _38240_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _88608_ (_38346_, _38242_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor _88609_ (_38347_, _38346_, _38345_);
  and _88610_ (_38349_, _38347_, _38344_);
  nor _88611_ (_38350_, _38349_, _38272_);
  and _88612_ (_38351_, _38234_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _88613_ (_38352_, _38236_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor _88614_ (_38353_, _38352_, _38351_);
  and _88615_ (_38354_, _38240_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _88616_ (_38355_, _38242_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor _88617_ (_38356_, _38355_, _38354_);
  and _88618_ (_38357_, _38356_, _38353_);
  nor _88619_ (_38358_, _38357_, _38258_);
  nor _88620_ (_38360_, _38358_, _38350_);
  and _88621_ (_38361_, _38234_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _88622_ (_38362_, _38236_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor _88623_ (_38363_, _38362_, _38361_);
  and _88624_ (_38364_, _38240_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _88625_ (_38365_, _38242_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor _88626_ (_38366_, _38365_, _38364_);
  and _88627_ (_38367_, _38366_, _38363_);
  nor _88628_ (_38368_, _38367_, _38247_);
  and _88629_ (_38369_, _38234_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _88630_ (_38371_, _38236_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor _88631_ (_38372_, _38371_, _38369_);
  and _88632_ (_38373_, _38240_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _88633_ (_38374_, _38242_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor _88634_ (_38375_, _38374_, _38373_);
  and _88635_ (_38376_, _38375_, _38372_);
  nor _88636_ (_38377_, _38376_, _38283_);
  nor _88637_ (_38378_, _38377_, _38368_);
  and _88638_ (_38379_, _38378_, _38360_);
  and _88639_ (_38380_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _88640_ (_38382_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _88641_ (_38383_, _38382_, _38380_);
  and _88642_ (_38384_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _88643_ (_38385_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _88644_ (_38386_, _38385_, _38384_);
  and _88645_ (_38387_, _38386_, _38383_);
  and _88646_ (_38388_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _88647_ (_38389_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _88648_ (_38390_, _38389_, _38388_);
  and _88649_ (_38391_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _88650_ (_38393_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _88651_ (_38394_, _38393_, _38391_);
  and _88652_ (_38395_, _38394_, _38390_);
  and _88653_ (_38396_, _38395_, _38387_);
  and _88654_ (_38397_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and _88655_ (_38398_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _88656_ (_38399_, _38398_, _38397_);
  and _88657_ (_38400_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _88658_ (_38401_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _88659_ (_38402_, _38401_, _38400_);
  and _88660_ (_38404_, _38402_, _38399_);
  and _88661_ (_38405_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _88662_ (_38406_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _88663_ (_38407_, _38406_, _38405_);
  and _88664_ (_38408_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _88665_ (_38409_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _88666_ (_38410_, _38409_, _38408_);
  and _88667_ (_38411_, _38410_, _38407_);
  and _88668_ (_38412_, _38411_, _38404_);
  and _88669_ (_38413_, _38412_, _38396_);
  nand _88670_ (_38415_, _38413_, _38379_);
  or _88671_ (_38416_, _38413_, _38379_);
  and _88672_ (_38417_, _38416_, _38415_);
  or _88673_ (_38418_, _38417_, _38341_);
  and _88674_ (_38419_, _38234_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _88675_ (_38420_, _38236_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor _88676_ (_38421_, _38420_, _38419_);
  and _88677_ (_38422_, _38240_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _88678_ (_38423_, _38242_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor _88679_ (_38424_, _38423_, _38422_);
  and _88680_ (_38426_, _38424_, _38421_);
  nor _88681_ (_38427_, _38426_, _38272_);
  and _88682_ (_38428_, _38234_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _88683_ (_38429_, _38236_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor _88684_ (_38430_, _38429_, _38428_);
  and _88685_ (_38431_, _38240_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _88686_ (_38432_, _38242_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor _88687_ (_38433_, _38432_, _38431_);
  and _88688_ (_38434_, _38433_, _38430_);
  nor _88689_ (_38435_, _38434_, _38283_);
  nor _88690_ (_38437_, _38435_, _38427_);
  and _88691_ (_38438_, _38234_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _88692_ (_38439_, _38236_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor _88693_ (_38440_, _38439_, _38438_);
  and _88694_ (_38441_, _38240_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _88695_ (_38442_, _38242_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor _88696_ (_38443_, _38442_, _38441_);
  and _88697_ (_38444_, _38443_, _38440_);
  nor _88698_ (_38445_, _38444_, _38247_);
  and _88699_ (_38446_, _38234_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _88700_ (_38448_, _38236_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor _88701_ (_38449_, _38448_, _38446_);
  and _88702_ (_38450_, _38240_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _88703_ (_38451_, _38242_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor _88704_ (_38452_, _38451_, _38450_);
  and _88705_ (_38453_, _38452_, _38449_);
  nor _88706_ (_38454_, _38453_, _38258_);
  nor _88707_ (_38455_, _38454_, _38445_);
  and _88708_ (_38456_, _38455_, _38437_);
  not _88709_ (_38457_, _38456_);
  and _88710_ (_38459_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _88711_ (_38460_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _88712_ (_38461_, _38460_, _38459_);
  and _88713_ (_38462_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _88714_ (_38463_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _88715_ (_38464_, _38463_, _38462_);
  and _88716_ (_38465_, _38464_, _38461_);
  and _88717_ (_38466_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _88718_ (_38467_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _88719_ (_38468_, _38467_, _38466_);
  and _88720_ (_38470_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _88721_ (_38471_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _88722_ (_38472_, _38471_, _38470_);
  and _88723_ (_38473_, _38472_, _38468_);
  and _88724_ (_38474_, _38473_, _38465_);
  and _88725_ (_38475_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and _88726_ (_38476_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _88727_ (_38477_, _38476_, _38475_);
  and _88728_ (_38478_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _88729_ (_38479_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _88730_ (_38481_, _38479_, _38478_);
  and _88731_ (_38482_, _38481_, _38477_);
  and _88732_ (_38483_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _88733_ (_38484_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _88734_ (_38485_, _38484_, _38483_);
  and _88735_ (_38486_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _88736_ (_38487_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _88737_ (_38488_, _38487_, _38486_);
  and _88738_ (_38489_, _38488_, _38485_);
  and _88739_ (_38490_, _38489_, _38482_);
  and _88740_ (_38492_, _38490_, _38474_);
  nor _88741_ (_38493_, _38492_, _38457_);
  and _88742_ (_38494_, _38492_, _38457_);
  or _88743_ (_38495_, _38494_, _38493_);
  and _88744_ (_38496_, _38234_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _88745_ (_38497_, _38236_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor _88746_ (_38498_, _38497_, _38496_);
  and _88747_ (_38499_, _38240_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _88748_ (_38500_, _38242_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor _88749_ (_38501_, _38500_, _38499_);
  and _88750_ (_38503_, _38501_, _38498_);
  nor _88751_ (_38504_, _38503_, _38247_);
  and _88752_ (_38505_, _38234_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _88753_ (_38506_, _38236_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor _88754_ (_38507_, _38506_, _38505_);
  and _88755_ (_38508_, _38240_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _88756_ (_38509_, _38242_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor _88757_ (_38510_, _38509_, _38508_);
  and _88758_ (_38511_, _38510_, _38507_);
  nor _88759_ (_38512_, _38511_, _38283_);
  nor _88760_ (_38514_, _38512_, _38504_);
  and _88761_ (_38515_, _38234_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _88762_ (_38516_, _38236_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor _88763_ (_38517_, _38516_, _38515_);
  and _88764_ (_38518_, _38240_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _88765_ (_38519_, _38242_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor _88766_ (_38520_, _38519_, _38518_);
  and _88767_ (_38521_, _38520_, _38517_);
  nor _88768_ (_38522_, _38521_, _38272_);
  and _88769_ (_38523_, _38234_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _88770_ (_38525_, _38236_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor _88771_ (_38526_, _38525_, _38523_);
  and _88772_ (_38527_, _38240_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _88773_ (_38528_, _38242_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor _88774_ (_38529_, _38528_, _38527_);
  and _88775_ (_38530_, _38529_, _38526_);
  nor _88776_ (_38531_, _38530_, _38258_);
  nor _88777_ (_38532_, _38531_, _38522_);
  and _88778_ (_38533_, _38532_, _38514_);
  and _88779_ (_38534_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _88780_ (_38536_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _88781_ (_38537_, _38536_, _38534_);
  and _88782_ (_38538_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _88783_ (_38539_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _88784_ (_38540_, _38539_, _38538_);
  and _88785_ (_38541_, _38540_, _38537_);
  and _88786_ (_38542_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _88787_ (_38543_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _88788_ (_38544_, _38543_, _38542_);
  and _88789_ (_38545_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _88790_ (_38547_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _88791_ (_38548_, _38547_, _38545_);
  and _88792_ (_38549_, _38548_, _38544_);
  and _88793_ (_38550_, _38549_, _38541_);
  and _88794_ (_38551_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _88795_ (_38552_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _88796_ (_38553_, _38552_, _38551_);
  and _88797_ (_38554_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _88798_ (_38555_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _88799_ (_38556_, _38555_, _38554_);
  and _88800_ (_38558_, _38556_, _38553_);
  and _88801_ (_38559_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and _88802_ (_38560_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _88803_ (_38561_, _38560_, _38559_);
  and _88804_ (_38562_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _88805_ (_38563_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _88806_ (_38564_, _38563_, _38562_);
  and _88807_ (_38565_, _38564_, _38561_);
  and _88808_ (_38566_, _38565_, _38558_);
  and _88809_ (_38567_, _38566_, _38550_);
  nand _88810_ (_38569_, _38567_, _38533_);
  or _88811_ (_38570_, _38567_, _38533_);
  and _88812_ (_38571_, _38570_, _38569_);
  or _88813_ (_38572_, _38571_, _38495_);
  or _88814_ (_38573_, _38572_, _38418_);
  and _88815_ (_38574_, _38234_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _88816_ (_38575_, _38236_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor _88817_ (_38576_, _38575_, _38574_);
  and _88818_ (_38577_, _38240_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _88819_ (_38578_, _38242_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor _88820_ (_38580_, _38578_, _38577_);
  and _88821_ (_38581_, _38580_, _38576_);
  nor _88822_ (_38582_, _38581_, _38272_);
  and _88823_ (_38583_, _38234_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _88824_ (_38584_, _38236_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor _88825_ (_38585_, _38584_, _38583_);
  and _88826_ (_38586_, _38240_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _88827_ (_38587_, _38242_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor _88828_ (_38588_, _38587_, _38586_);
  and _88829_ (_38589_, _38588_, _38585_);
  nor _88830_ (_38591_, _38589_, _38283_);
  nor _88831_ (_38592_, _38591_, _38582_);
  and _88832_ (_38593_, _38234_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _88833_ (_38594_, _38236_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor _88834_ (_38595_, _38594_, _38593_);
  and _88835_ (_38596_, _38240_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _88836_ (_38597_, _38242_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor _88837_ (_38598_, _38597_, _38596_);
  and _88838_ (_38599_, _38598_, _38595_);
  nor _88839_ (_38600_, _38599_, _38247_);
  and _88840_ (_38602_, _38234_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _88841_ (_38603_, _38236_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor _88842_ (_38604_, _38603_, _38602_);
  and _88843_ (_38605_, _38240_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _88844_ (_38606_, _38242_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor _88845_ (_38607_, _38606_, _38605_);
  and _88846_ (_38608_, _38607_, _38604_);
  nor _88847_ (_38609_, _38608_, _38258_);
  nor _88848_ (_38610_, _38609_, _38600_);
  and _88849_ (_38611_, _38610_, _38592_);
  and _88850_ (_38613_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and _88851_ (_38614_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _88852_ (_38615_, _38614_, _38613_);
  and _88853_ (_38616_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _88854_ (_38617_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _88855_ (_38618_, _38617_, _38616_);
  and _88856_ (_38619_, _38618_, _38615_);
  and _88857_ (_38620_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _88858_ (_38621_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _88859_ (_38622_, _38621_, _38620_);
  and _88860_ (_38624_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _88861_ (_38625_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _88862_ (_38626_, _38625_, _38624_);
  and _88863_ (_38627_, _38626_, _38622_);
  and _88864_ (_38628_, _38627_, _38619_);
  and _88865_ (_38629_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _88866_ (_38630_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _88867_ (_38631_, _38630_, _38629_);
  and _88868_ (_38632_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _88869_ (_38633_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _88870_ (_38635_, _38633_, _38632_);
  and _88871_ (_38636_, _38635_, _38631_);
  and _88872_ (_38637_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _88873_ (_38638_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _88874_ (_38639_, _38638_, _38637_);
  and _88875_ (_38640_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _88876_ (_38641_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _88877_ (_38642_, _38641_, _38640_);
  and _88878_ (_38643_, _38642_, _38639_);
  and _88879_ (_38644_, _38643_, _38636_);
  and _88880_ (_38646_, _38644_, _38628_);
  or _88881_ (_38647_, _38646_, _38611_);
  nand _88882_ (_38648_, _38646_, _38611_);
  and _88883_ (_38649_, _38648_, _38647_);
  and _88884_ (_38650_, _38234_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _88885_ (_38651_, _38236_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor _88886_ (_38652_, _38651_, _38650_);
  and _88887_ (_38653_, _38240_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _88888_ (_38654_, _38242_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor _88889_ (_38655_, _38654_, _38653_);
  and _88890_ (_38657_, _38655_, _38652_);
  nor _88891_ (_38658_, _38657_, _38272_);
  and _88892_ (_38659_, _38234_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _88893_ (_38660_, _38236_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor _88894_ (_38661_, _38660_, _38659_);
  and _88895_ (_38662_, _38240_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _88896_ (_38663_, _38242_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor _88897_ (_38664_, _38663_, _38662_);
  and _88898_ (_38665_, _38664_, _38661_);
  nor _88899_ (_38666_, _38665_, _38258_);
  nor _88900_ (_38668_, _38666_, _38658_);
  and _88901_ (_38669_, _38234_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _88902_ (_38670_, _38236_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor _88903_ (_38671_, _38670_, _38669_);
  and _88904_ (_38672_, _38240_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _88905_ (_38673_, _38242_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor _88906_ (_38674_, _38673_, _38672_);
  and _88907_ (_38675_, _38674_, _38671_);
  nor _88908_ (_38676_, _38675_, _38247_);
  and _88909_ (_38677_, _38234_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _88910_ (_38679_, _38236_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor _88911_ (_38680_, _38679_, _38677_);
  and _88912_ (_38681_, _38240_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _88913_ (_38682_, _38242_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor _88914_ (_38683_, _38682_, _38681_);
  and _88915_ (_38684_, _38683_, _38680_);
  nor _88916_ (_38685_, _38684_, _38283_);
  nor _88917_ (_38686_, _38685_, _38676_);
  and _88918_ (_38687_, _38686_, _38668_);
  and _88919_ (_38688_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _88920_ (_38690_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _88921_ (_38691_, _38690_, _38688_);
  and _88922_ (_38692_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _88923_ (_38693_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _88924_ (_38694_, _38693_, _38692_);
  and _88925_ (_38695_, _38694_, _38691_);
  and _88926_ (_38696_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _88927_ (_38697_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _88928_ (_38698_, _38697_, _38696_);
  and _88929_ (_38699_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _88930_ (_38701_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _88931_ (_38702_, _38701_, _38699_);
  and _88932_ (_38703_, _38702_, _38698_);
  and _88933_ (_38704_, _38703_, _38695_);
  and _88934_ (_38705_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and _88935_ (_38706_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _88936_ (_38707_, _38706_, _38705_);
  and _88937_ (_38708_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _88938_ (_38709_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _88939_ (_38710_, _38709_, _38708_);
  and _88940_ (_38712_, _38710_, _38707_);
  and _88941_ (_38713_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _88942_ (_38714_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _88943_ (_38715_, _38714_, _38713_);
  and _88944_ (_38716_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _88945_ (_38717_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _88946_ (_38718_, _38717_, _38716_);
  and _88947_ (_38719_, _38718_, _38715_);
  and _88948_ (_38720_, _38719_, _38712_);
  and _88949_ (_38721_, _38720_, _38704_);
  nand _88950_ (_38723_, _38721_, _38687_);
  or _88951_ (_38724_, _38721_, _38687_);
  and _88952_ (_38725_, _38724_, _38723_);
  or _88953_ (_38726_, _38725_, _38649_);
  and _88954_ (_38727_, _38234_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _88955_ (_38728_, _38236_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor _88956_ (_38729_, _38728_, _38727_);
  and _88957_ (_38730_, _38240_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _88958_ (_38731_, _38242_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor _88959_ (_38732_, _38731_, _38730_);
  and _88960_ (_38734_, _38732_, _38729_);
  nor _88961_ (_38735_, _38734_, _38272_);
  and _88962_ (_38736_, _38234_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _88963_ (_38737_, _38236_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor _88964_ (_38738_, _38737_, _38736_);
  and _88965_ (_38739_, _38240_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _88966_ (_38740_, _38242_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor _88967_ (_38741_, _38740_, _38739_);
  and _88968_ (_38742_, _38741_, _38738_);
  nor _88969_ (_38743_, _38742_, _38258_);
  nor _88970_ (_38745_, _38743_, _38735_);
  and _88971_ (_38746_, _38234_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _88972_ (_38747_, _38236_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _88973_ (_38748_, _38747_, _38746_);
  and _88974_ (_38749_, _38240_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _88975_ (_38750_, _38242_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor _88976_ (_38751_, _38750_, _38749_);
  and _88977_ (_38752_, _38751_, _38748_);
  nor _88978_ (_38753_, _38752_, _38247_);
  and _88979_ (_38754_, _38234_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _88980_ (_38756_, _38236_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor _88981_ (_38757_, _38756_, _38754_);
  and _88982_ (_38758_, _38240_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _88983_ (_38759_, _38242_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor _88984_ (_38760_, _38759_, _38758_);
  and _88985_ (_38761_, _38760_, _38757_);
  nor _88986_ (_38762_, _38761_, _38283_);
  nor _88987_ (_38763_, _38762_, _38753_);
  and _88988_ (_38764_, _38763_, _38745_);
  and _88989_ (_38765_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _88990_ (_38767_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor _88991_ (_38768_, _38767_, _38765_);
  and _88992_ (_38769_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _88993_ (_38770_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _88994_ (_38771_, _38770_, _38769_);
  and _88995_ (_38772_, _38771_, _38768_);
  and _88996_ (_38773_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and _88997_ (_38774_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _88998_ (_38775_, _38774_, _38773_);
  and _88999_ (_38776_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _89000_ (_38778_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _89001_ (_38779_, _38778_, _38776_);
  and _89002_ (_38780_, _38779_, _38775_);
  and _89003_ (_38781_, _38780_, _38772_);
  and _89004_ (_38782_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _89005_ (_38783_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _89006_ (_38784_, _38783_, _38782_);
  and _89007_ (_38785_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _89008_ (_38786_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _89009_ (_38787_, _38786_, _38785_);
  and _89010_ (_38789_, _38787_, _38784_);
  and _89011_ (_38790_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _89012_ (_38791_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor _89013_ (_38792_, _38791_, _38790_);
  and _89014_ (_38793_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and _89015_ (_38794_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _89016_ (_38795_, _38794_, _38793_);
  and _89017_ (_38796_, _38795_, _38792_);
  and _89018_ (_38797_, _38796_, _38789_);
  and _89019_ (_38798_, _38797_, _38781_);
  nand _89020_ (_38800_, _38798_, _38764_);
  or _89021_ (_38801_, _38798_, _38764_);
  and _89022_ (_38802_, _38801_, _38800_);
  and _89023_ (_38803_, _38234_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _89024_ (_38804_, _38236_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor _89025_ (_38805_, _38804_, _38803_);
  and _89026_ (_38806_, _38240_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _89027_ (_38807_, _38242_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor _89028_ (_38808_, _38807_, _38806_);
  and _89029_ (_38809_, _38808_, _38805_);
  nor _89030_ (_38811_, _38809_, _38247_);
  and _89031_ (_38812_, _38234_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _89032_ (_38813_, _38236_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor _89033_ (_38814_, _38813_, _38812_);
  and _89034_ (_38815_, _38240_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _89035_ (_38816_, _38242_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor _89036_ (_38817_, _38816_, _38815_);
  and _89037_ (_38818_, _38817_, _38814_);
  nor _89038_ (_38819_, _38818_, _38283_);
  nor _89039_ (_38820_, _38819_, _38811_);
  and _89040_ (_38822_, _38234_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _89041_ (_38823_, _38236_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor _89042_ (_38824_, _38823_, _38822_);
  and _89043_ (_38825_, _38240_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _89044_ (_38826_, _38242_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor _89045_ (_38827_, _38826_, _38825_);
  and _89046_ (_38828_, _38827_, _38824_);
  nor _89047_ (_38829_, _38828_, _38272_);
  and _89048_ (_38830_, _38234_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _89049_ (_38831_, _38236_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor _89050_ (_38833_, _38831_, _38830_);
  and _89051_ (_38834_, _38240_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _89052_ (_38835_, _38242_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor _89053_ (_38836_, _38835_, _38834_);
  and _89054_ (_38837_, _38836_, _38833_);
  nor _89055_ (_38838_, _38837_, _38258_);
  nor _89056_ (_38839_, _38838_, _38829_);
  and _89057_ (_38840_, _38839_, _38820_);
  and _89058_ (_38841_, _38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _89059_ (_38842_, _38327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _89060_ (_38844_, _38842_, _38841_);
  and _89061_ (_38845_, _38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _89062_ (_38846_, _38301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _89063_ (_38847_, _38846_, _38845_);
  and _89064_ (_38848_, _38847_, _38844_);
  and _89065_ (_38849_, _38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _89066_ (_38850_, _38287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _89067_ (_38851_, _38850_, _38849_);
  and _89068_ (_38852_, _38324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _89069_ (_38853_, _38330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _89070_ (_38855_, _38853_, _38852_);
  and _89071_ (_38856_, _38855_, _38851_);
  and _89072_ (_38857_, _38856_, _38848_);
  and _89073_ (_38858_, _38305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and _89074_ (_38859_, _38320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _89075_ (_38860_, _38859_, _38858_);
  and _89076_ (_38861_, _38295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _89077_ (_38862_, _38289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _89078_ (_38863_, _38862_, _38861_);
  and _89079_ (_38864_, _38863_, _38860_);
  and _89080_ (_38866_, _38292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _89081_ (_38867_, _38299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _89082_ (_38868_, _38867_, _38866_);
  and _89083_ (_38869_, _38332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _89084_ (_38870_, _38307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _89085_ (_38871_, _38870_, _38869_);
  and _89086_ (_38872_, _38871_, _38868_);
  and _89087_ (_38873_, _38872_, _38864_);
  and _89088_ (_38874_, _38873_, _38857_);
  not _89089_ (_38875_, _38874_);
  nor _89090_ (_38877_, _38875_, _38840_);
  and _89091_ (_38878_, _38875_, _38840_);
  or _89092_ (_38879_, _38878_, _38877_);
  or _89093_ (_38880_, _38879_, _38802_);
  or _89094_ (_38881_, _38880_, _38726_);
  or _89095_ (_38882_, _38881_, _38573_);
  and _89096_ (property_invalid_iram, _38882_, _38232_);
  and _89097_ (_38883_, \oc8051_golden_model_1.ACC [2], _39990_);
  and _89098_ (_38884_, _10280_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _89099_ (_38885_, _38884_, _38883_);
  nand _89100_ (_38887_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _89101_ (_38888_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _89102_ (_38889_, _38888_, _38887_);
  or _89103_ (_38890_, _38889_, _38885_);
  and _89104_ (_38891_, _06097_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _89105_ (_38892_, \oc8051_golden_model_1.ACC [1], _39970_);
  or _89106_ (_38893_, _38892_, _38891_);
  and _89107_ (_38894_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _89108_ (_38895_, \oc8051_golden_model_1.ACC [0], _39951_);
  or _89109_ (_38896_, _38895_, _38894_);
  or _89110_ (_38898_, _38896_, _38893_);
  or _89111_ (_38899_, _38898_, _38890_);
  or _89112_ (_38900_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _89113_ (_38901_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _89114_ (_38902_, _38901_, _38900_);
  or _89115_ (_38903_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _89116_ (_38904_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _89117_ (_38905_, _38904_, _38903_);
  or _89118_ (_38906_, _38905_, _38902_);
  nand _89119_ (_38907_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _89120_ (_38909_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _89121_ (_38910_, _38909_, _38907_);
  and _89122_ (_38911_, _08688_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _89123_ (_38912_, _08688_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _89124_ (_38913_, _38912_, _38911_);
  or _89125_ (_38914_, _38913_, _38910_);
  or _89126_ (_38915_, _38914_, _38906_);
  or _89127_ (_38916_, _38915_, _38899_);
  and _89128_ (property_invalid_acc, _38916_, _38232_);
  and _89129_ (_38917_, _38230_, _01442_);
  nor _89130_ (_38919_, _25815_, _02061_);
  and _89131_ (_38920_, _25815_, _02061_);
  and _89132_ (_38921_, _26175_, _02065_);
  nor _89133_ (_38922_, _26175_, _02065_);
  nor _89134_ (_38923_, _26878_, _02073_);
  and _89135_ (_38924_, _26878_, _02073_);
  or _89136_ (_38925_, _38924_, _38923_);
  and _89137_ (_38926_, _27576_, _02081_);
  nand _89138_ (_38927_, _28581_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _89139_ (_38928_, _28581_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _89140_ (_38930_, _38928_, _38927_);
  nand _89141_ (_38931_, _28254_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _89142_ (_38932_, _28254_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _89143_ (_38933_, _38932_, _38931_);
  and _89144_ (_38934_, _28881_, _39397_);
  nor _89145_ (_38935_, _28881_, _39397_);
  or _89146_ (_38936_, _38935_, _38934_);
  nor _89147_ (_38937_, _13112_, _39414_);
  and _89148_ (_38938_, _13112_, _39414_);
  or _89149_ (_38939_, _38938_, _38937_);
  or _89150_ (_38941_, _38939_, _38936_);
  and _89151_ (_38942_, _29185_, _39382_);
  nor _89152_ (_38943_, _29185_, _39382_);
  or _89153_ (_38944_, _38943_, _38942_);
  nor _89154_ (_38945_, _29793_, _39378_);
  and _89155_ (_38946_, _29793_, _39378_);
  nor _89156_ (_38947_, _29488_, _39403_);
  and _89157_ (_38948_, _29488_, _39403_);
  or _89158_ (_38949_, _38948_, _38947_);
  and _89159_ (_38950_, _30091_, _39409_);
  or _89160_ (_38952_, _25424_, _02057_);
  nand _89161_ (_38953_, _25424_, _02057_);
  and _89162_ (_38954_, _38953_, _38952_);
  nor _89163_ (_38955_, _30091_, _39409_);
  or _89164_ (_38956_, _38955_, _38954_);
  or _89165_ (_38957_, _38956_, _38950_);
  or _89166_ (_38958_, _38957_, _38949_);
  or _89167_ (_38959_, _38958_, _38946_);
  or _89168_ (_38960_, _38959_, _38945_);
  or _89169_ (_38961_, _38960_, _38944_);
  or _89170_ (_38963_, _38961_, _38941_);
  or _89171_ (_38964_, _38963_, _38933_);
  or _89172_ (_38965_, _38964_, _38930_);
  or _89173_ (_38966_, _38965_, _38926_);
  and _89174_ (_38967_, _26523_, _02069_);
  nor _89175_ (_38968_, _27233_, _02077_);
  or _89176_ (_38969_, _38968_, _38967_);
  or _89177_ (_38970_, _38969_, _38966_);
  or _89178_ (_38971_, _38970_, _38925_);
  and _89179_ (_38972_, _27929_, _02085_);
  nor _89180_ (_38974_, _27929_, _02085_);
  and _89181_ (_38975_, _27233_, _02077_);
  nor _89182_ (_38976_, _26523_, _02069_);
  nor _89183_ (_38977_, _27576_, _02081_);
  or _89184_ (_38978_, _38977_, _38976_);
  or _89185_ (_38979_, _38978_, _38975_);
  or _89186_ (_38980_, _38979_, _38974_);
  or _89187_ (_38981_, _38980_, _38972_);
  or _89188_ (_38982_, _38981_, _38971_);
  or _89189_ (_38983_, _38982_, _38922_);
  or _89190_ (_38985_, _38983_, _38921_);
  or _89191_ (_38986_, _38985_, _38920_);
  or _89192_ (_38987_, _38986_, _38919_);
  and _89193_ (property_invalid_pc, _38987_, _38917_);
  buf _89194_ (_00550_, _43637_);
  buf _89195_ (_05099_, _43634_);
  buf _89196_ (_05150_, _43634_);
  buf _89197_ (_05202_, _43634_);
  buf _89198_ (_05254_, _43634_);
  buf _89199_ (_05305_, _43634_);
  buf _89200_ (_05357_, _43634_);
  buf _89201_ (_05408_, _43634_);
  buf _89202_ (_05460_, _43634_);
  buf _89203_ (_05512_, _43634_);
  buf _89204_ (_05563_, _43634_);
  buf _89205_ (_05615_, _43634_);
  buf _89206_ (_05666_, _43634_);
  buf _89207_ (_05719_, _43634_);
  buf _89208_ (_05772_, _43634_);
  buf _89209_ (_05825_, _43634_);
  buf _89210_ (_05878_, _43634_);
  buf _89211_ (_39793_, _39696_);
  buf _89212_ (_39795_, _39698_);
  buf _89213_ (_39808_, _39696_);
  buf _89214_ (_39809_, _39698_);
  buf _89215_ (_40122_, _39714_);
  buf _89216_ (_40123_, _39715_);
  buf _89217_ (_40124_, _39717_);
  buf _89218_ (_40125_, _39718_);
  buf _89219_ (_40126_, _39719_);
  buf _89220_ (_40127_, _39720_);
  buf _89221_ (_40128_, _39721_);
  buf _89222_ (_40129_, _39722_);
  buf _89223_ (_40130_, _39723_);
  buf _89224_ (_40132_, _39724_);
  buf _89225_ (_40133_, _39725_);
  buf _89226_ (_40134_, _39726_);
  buf _89227_ (_40135_, _39728_);
  buf _89228_ (_40136_, _39729_);
  buf _89229_ (_40188_, _39714_);
  buf _89230_ (_40189_, _39715_);
  buf _89231_ (_40190_, _39717_);
  buf _89232_ (_40191_, _39718_);
  buf _89233_ (_40192_, _39719_);
  buf _89234_ (_40193_, _39720_);
  buf _89235_ (_40194_, _39721_);
  buf _89236_ (_40195_, _39722_);
  buf _89237_ (_40196_, _39723_);
  buf _89238_ (_40198_, _39724_);
  buf _89239_ (_40199_, _39725_);
  buf _89240_ (_40200_, _39726_);
  buf _89241_ (_40201_, _39728_);
  buf _89242_ (_40202_, _39729_);
  buf _89243_ (_40596_, _40499_);
  buf _89244_ (_40753_, _40499_);
  dff _89245_ (p0in_reg[0], _00002_[0], clk);
  dff _89246_ (p0in_reg[1], _00002_[1], clk);
  dff _89247_ (p0in_reg[2], _00002_[2], clk);
  dff _89248_ (p0in_reg[3], _00002_[3], clk);
  dff _89249_ (p0in_reg[4], _00002_[4], clk);
  dff _89250_ (p0in_reg[5], _00002_[5], clk);
  dff _89251_ (p0in_reg[6], _00002_[6], clk);
  dff _89252_ (p0in_reg[7], _00002_[7], clk);
  dff _89253_ (p1in_reg[0], _00003_[0], clk);
  dff _89254_ (p1in_reg[1], _00003_[1], clk);
  dff _89255_ (p1in_reg[2], _00003_[2], clk);
  dff _89256_ (p1in_reg[3], _00003_[3], clk);
  dff _89257_ (p1in_reg[4], _00003_[4], clk);
  dff _89258_ (p1in_reg[5], _00003_[5], clk);
  dff _89259_ (p1in_reg[6], _00003_[6], clk);
  dff _89260_ (p1in_reg[7], _00003_[7], clk);
  dff _89261_ (p2in_reg[0], _00004_[0], clk);
  dff _89262_ (p2in_reg[1], _00004_[1], clk);
  dff _89263_ (p2in_reg[2], _00004_[2], clk);
  dff _89264_ (p2in_reg[3], _00004_[3], clk);
  dff _89265_ (p2in_reg[4], _00004_[4], clk);
  dff _89266_ (p2in_reg[5], _00004_[5], clk);
  dff _89267_ (p2in_reg[6], _00004_[6], clk);
  dff _89268_ (p2in_reg[7], _00004_[7], clk);
  dff _89269_ (p3in_reg[0], _00005_[0], clk);
  dff _89270_ (p3in_reg[1], _00005_[1], clk);
  dff _89271_ (p3in_reg[2], _00005_[2], clk);
  dff _89272_ (p3in_reg[3], _00005_[3], clk);
  dff _89273_ (p3in_reg[4], _00005_[4], clk);
  dff _89274_ (p3in_reg[5], _00005_[5], clk);
  dff _89275_ (p3in_reg[6], _00005_[6], clk);
  dff _89276_ (p3in_reg[7], _00005_[7], clk);
  dff _89277_ (op0_cnst, _00001_, clk);
  dff _89278_ (inst_finished_r, _00000_, clk);
  dff _89279_ (\oc8051_gm_cxrom_1.cell0.data [0], _05103_, clk);
  dff _89280_ (\oc8051_gm_cxrom_1.cell0.data [1], _05107_, clk);
  dff _89281_ (\oc8051_gm_cxrom_1.cell0.data [2], _05111_, clk);
  dff _89282_ (\oc8051_gm_cxrom_1.cell0.data [3], _05115_, clk);
  dff _89283_ (\oc8051_gm_cxrom_1.cell0.data [4], _05118_, clk);
  dff _89284_ (\oc8051_gm_cxrom_1.cell0.data [5], _05122_, clk);
  dff _89285_ (\oc8051_gm_cxrom_1.cell0.data [6], _05126_, clk);
  dff _89286_ (\oc8051_gm_cxrom_1.cell0.data [7], _05096_, clk);
  dff _89287_ (\oc8051_gm_cxrom_1.cell0.valid , _05099_, clk);
  dff _89288_ (\oc8051_gm_cxrom_1.cell1.data [0], _05154_, clk);
  dff _89289_ (\oc8051_gm_cxrom_1.cell1.data [1], _05158_, clk);
  dff _89290_ (\oc8051_gm_cxrom_1.cell1.data [2], _05162_, clk);
  dff _89291_ (\oc8051_gm_cxrom_1.cell1.data [3], _05166_, clk);
  dff _89292_ (\oc8051_gm_cxrom_1.cell1.data [4], _05170_, clk);
  dff _89293_ (\oc8051_gm_cxrom_1.cell1.data [5], _05174_, clk);
  dff _89294_ (\oc8051_gm_cxrom_1.cell1.data [6], _05178_, clk);
  dff _89295_ (\oc8051_gm_cxrom_1.cell1.data [7], _05148_, clk);
  dff _89296_ (\oc8051_gm_cxrom_1.cell1.valid , _05150_, clk);
  dff _89297_ (\oc8051_gm_cxrom_1.cell10.data [0], _05619_, clk);
  dff _89298_ (\oc8051_gm_cxrom_1.cell10.data [1], _05623_, clk);
  dff _89299_ (\oc8051_gm_cxrom_1.cell10.data [2], _05626_, clk);
  dff _89300_ (\oc8051_gm_cxrom_1.cell10.data [3], _05630_, clk);
  dff _89301_ (\oc8051_gm_cxrom_1.cell10.data [4], _05634_, clk);
  dff _89302_ (\oc8051_gm_cxrom_1.cell10.data [5], _05638_, clk);
  dff _89303_ (\oc8051_gm_cxrom_1.cell10.data [6], _05642_, clk);
  dff _89304_ (\oc8051_gm_cxrom_1.cell10.data [7], _05612_, clk);
  dff _89305_ (\oc8051_gm_cxrom_1.cell10.valid , _05615_, clk);
  dff _89306_ (\oc8051_gm_cxrom_1.cell11.data [0], _05670_, clk);
  dff _89307_ (\oc8051_gm_cxrom_1.cell11.data [1], _05674_, clk);
  dff _89308_ (\oc8051_gm_cxrom_1.cell11.data [2], _05678_, clk);
  dff _89309_ (\oc8051_gm_cxrom_1.cell11.data [3], _05682_, clk);
  dff _89310_ (\oc8051_gm_cxrom_1.cell11.data [4], _05686_, clk);
  dff _89311_ (\oc8051_gm_cxrom_1.cell11.data [5], _05690_, clk);
  dff _89312_ (\oc8051_gm_cxrom_1.cell11.data [6], _05694_, clk);
  dff _89313_ (\oc8051_gm_cxrom_1.cell11.data [7], _05663_, clk);
  dff _89314_ (\oc8051_gm_cxrom_1.cell11.valid , _05666_, clk);
  dff _89315_ (\oc8051_gm_cxrom_1.cell12.data [0], _05723_, clk);
  dff _89316_ (\oc8051_gm_cxrom_1.cell12.data [1], _05727_, clk);
  dff _89317_ (\oc8051_gm_cxrom_1.cell12.data [2], _05731_, clk);
  dff _89318_ (\oc8051_gm_cxrom_1.cell12.data [3], _05735_, clk);
  dff _89319_ (\oc8051_gm_cxrom_1.cell12.data [4], _05739_, clk);
  dff _89320_ (\oc8051_gm_cxrom_1.cell12.data [5], _05743_, clk);
  dff _89321_ (\oc8051_gm_cxrom_1.cell12.data [6], _05747_, clk);
  dff _89322_ (\oc8051_gm_cxrom_1.cell12.data [7], _05716_, clk);
  dff _89323_ (\oc8051_gm_cxrom_1.cell12.valid , _05719_, clk);
  dff _89324_ (\oc8051_gm_cxrom_1.cell13.data [0], _05776_, clk);
  dff _89325_ (\oc8051_gm_cxrom_1.cell13.data [1], _05780_, clk);
  dff _89326_ (\oc8051_gm_cxrom_1.cell13.data [2], _05784_, clk);
  dff _89327_ (\oc8051_gm_cxrom_1.cell13.data [3], _05788_, clk);
  dff _89328_ (\oc8051_gm_cxrom_1.cell13.data [4], _05792_, clk);
  dff _89329_ (\oc8051_gm_cxrom_1.cell13.data [5], _05796_, clk);
  dff _89330_ (\oc8051_gm_cxrom_1.cell13.data [6], _05800_, clk);
  dff _89331_ (\oc8051_gm_cxrom_1.cell13.data [7], _05769_, clk);
  dff _89332_ (\oc8051_gm_cxrom_1.cell13.valid , _05772_, clk);
  dff _89333_ (\oc8051_gm_cxrom_1.cell14.data [0], _05829_, clk);
  dff _89334_ (\oc8051_gm_cxrom_1.cell14.data [1], _05833_, clk);
  dff _89335_ (\oc8051_gm_cxrom_1.cell14.data [2], _05837_, clk);
  dff _89336_ (\oc8051_gm_cxrom_1.cell14.data [3], _05841_, clk);
  dff _89337_ (\oc8051_gm_cxrom_1.cell14.data [4], _05845_, clk);
  dff _89338_ (\oc8051_gm_cxrom_1.cell14.data [5], _05849_, clk);
  dff _89339_ (\oc8051_gm_cxrom_1.cell14.data [6], _05853_, clk);
  dff _89340_ (\oc8051_gm_cxrom_1.cell14.data [7], _05822_, clk);
  dff _89341_ (\oc8051_gm_cxrom_1.cell14.valid , _05825_, clk);
  dff _89342_ (\oc8051_gm_cxrom_1.cell15.data [0], _05882_, clk);
  dff _89343_ (\oc8051_gm_cxrom_1.cell15.data [1], _05886_, clk);
  dff _89344_ (\oc8051_gm_cxrom_1.cell15.data [2], _05890_, clk);
  dff _89345_ (\oc8051_gm_cxrom_1.cell15.data [3], _05894_, clk);
  dff _89346_ (\oc8051_gm_cxrom_1.cell15.data [4], _05898_, clk);
  dff _89347_ (\oc8051_gm_cxrom_1.cell15.data [5], _05902_, clk);
  dff _89348_ (\oc8051_gm_cxrom_1.cell15.data [6], _05906_, clk);
  dff _89349_ (\oc8051_gm_cxrom_1.cell15.data [7], _05875_, clk);
  dff _89350_ (\oc8051_gm_cxrom_1.cell15.valid , _05878_, clk);
  dff _89351_ (\oc8051_gm_cxrom_1.cell2.data [0], _05206_, clk);
  dff _89352_ (\oc8051_gm_cxrom_1.cell2.data [1], _05210_, clk);
  dff _89353_ (\oc8051_gm_cxrom_1.cell2.data [2], _05214_, clk);
  dff _89354_ (\oc8051_gm_cxrom_1.cell2.data [3], _05218_, clk);
  dff _89355_ (\oc8051_gm_cxrom_1.cell2.data [4], _05222_, clk);
  dff _89356_ (\oc8051_gm_cxrom_1.cell2.data [5], _05225_, clk);
  dff _89357_ (\oc8051_gm_cxrom_1.cell2.data [6], _05229_, clk);
  dff _89358_ (\oc8051_gm_cxrom_1.cell2.data [7], _05199_, clk);
  dff _89359_ (\oc8051_gm_cxrom_1.cell2.valid , _05202_, clk);
  dff _89360_ (\oc8051_gm_cxrom_1.cell3.data [0], _05258_, clk);
  dff _89361_ (\oc8051_gm_cxrom_1.cell3.data [1], _05261_, clk);
  dff _89362_ (\oc8051_gm_cxrom_1.cell3.data [2], _05265_, clk);
  dff _89363_ (\oc8051_gm_cxrom_1.cell3.data [3], _05269_, clk);
  dff _89364_ (\oc8051_gm_cxrom_1.cell3.data [4], _05273_, clk);
  dff _89365_ (\oc8051_gm_cxrom_1.cell3.data [5], _05277_, clk);
  dff _89366_ (\oc8051_gm_cxrom_1.cell3.data [6], _05281_, clk);
  dff _89367_ (\oc8051_gm_cxrom_1.cell3.data [7], _05251_, clk);
  dff _89368_ (\oc8051_gm_cxrom_1.cell3.valid , _05254_, clk);
  dff _89369_ (\oc8051_gm_cxrom_1.cell4.data [0], _05309_, clk);
  dff _89370_ (\oc8051_gm_cxrom_1.cell4.data [1], _05313_, clk);
  dff _89371_ (\oc8051_gm_cxrom_1.cell4.data [2], _05317_, clk);
  dff _89372_ (\oc8051_gm_cxrom_1.cell4.data [3], _05321_, clk);
  dff _89373_ (\oc8051_gm_cxrom_1.cell4.data [4], _05325_, clk);
  dff _89374_ (\oc8051_gm_cxrom_1.cell4.data [5], _05329_, clk);
  dff _89375_ (\oc8051_gm_cxrom_1.cell4.data [6], _05333_, clk);
  dff _89376_ (\oc8051_gm_cxrom_1.cell4.data [7], _05302_, clk);
  dff _89377_ (\oc8051_gm_cxrom_1.cell4.valid , _05305_, clk);
  dff _89378_ (\oc8051_gm_cxrom_1.cell5.data [0], _05361_, clk);
  dff _89379_ (\oc8051_gm_cxrom_1.cell5.data [1], _05365_, clk);
  dff _89380_ (\oc8051_gm_cxrom_1.cell5.data [2], _05369_, clk);
  dff _89381_ (\oc8051_gm_cxrom_1.cell5.data [3], _05372_, clk);
  dff _89382_ (\oc8051_gm_cxrom_1.cell5.data [4], _05376_, clk);
  dff _89383_ (\oc8051_gm_cxrom_1.cell5.data [5], _05380_, clk);
  dff _89384_ (\oc8051_gm_cxrom_1.cell5.data [6], _05384_, clk);
  dff _89385_ (\oc8051_gm_cxrom_1.cell5.data [7], _05354_, clk);
  dff _89386_ (\oc8051_gm_cxrom_1.cell5.valid , _05357_, clk);
  dff _89387_ (\oc8051_gm_cxrom_1.cell6.data [0], _05412_, clk);
  dff _89388_ (\oc8051_gm_cxrom_1.cell6.data [1], _05416_, clk);
  dff _89389_ (\oc8051_gm_cxrom_1.cell6.data [2], _05420_, clk);
  dff _89390_ (\oc8051_gm_cxrom_1.cell6.data [3], _05424_, clk);
  dff _89391_ (\oc8051_gm_cxrom_1.cell6.data [4], _05428_, clk);
  dff _89392_ (\oc8051_gm_cxrom_1.cell6.data [5], _05432_, clk);
  dff _89393_ (\oc8051_gm_cxrom_1.cell6.data [6], _05436_, clk);
  dff _89394_ (\oc8051_gm_cxrom_1.cell6.data [7], _05405_, clk);
  dff _89395_ (\oc8051_gm_cxrom_1.cell6.valid , _05408_, clk);
  dff _89396_ (\oc8051_gm_cxrom_1.cell7.data [0], _05464_, clk);
  dff _89397_ (\oc8051_gm_cxrom_1.cell7.data [1], _05468_, clk);
  dff _89398_ (\oc8051_gm_cxrom_1.cell7.data [2], _05472_, clk);
  dff _89399_ (\oc8051_gm_cxrom_1.cell7.data [3], _05476_, clk);
  dff _89400_ (\oc8051_gm_cxrom_1.cell7.data [4], _05479_, clk);
  dff _89401_ (\oc8051_gm_cxrom_1.cell7.data [5], _05483_, clk);
  dff _89402_ (\oc8051_gm_cxrom_1.cell7.data [6], _05487_, clk);
  dff _89403_ (\oc8051_gm_cxrom_1.cell7.data [7], _05457_, clk);
  dff _89404_ (\oc8051_gm_cxrom_1.cell7.valid , _05460_, clk);
  dff _89405_ (\oc8051_gm_cxrom_1.cell8.data [0], _05515_, clk);
  dff _89406_ (\oc8051_gm_cxrom_1.cell8.data [1], _05519_, clk);
  dff _89407_ (\oc8051_gm_cxrom_1.cell8.data [2], _05523_, clk);
  dff _89408_ (\oc8051_gm_cxrom_1.cell8.data [3], _05527_, clk);
  dff _89409_ (\oc8051_gm_cxrom_1.cell8.data [4], _05531_, clk);
  dff _89410_ (\oc8051_gm_cxrom_1.cell8.data [5], _05535_, clk);
  dff _89411_ (\oc8051_gm_cxrom_1.cell8.data [6], _05539_, clk);
  dff _89412_ (\oc8051_gm_cxrom_1.cell8.data [7], _05509_, clk);
  dff _89413_ (\oc8051_gm_cxrom_1.cell8.valid , _05512_, clk);
  dff _89414_ (\oc8051_gm_cxrom_1.cell9.data [0], _05567_, clk);
  dff _89415_ (\oc8051_gm_cxrom_1.cell9.data [1], _05571_, clk);
  dff _89416_ (\oc8051_gm_cxrom_1.cell9.data [2], _05575_, clk);
  dff _89417_ (\oc8051_gm_cxrom_1.cell9.data [3], _05579_, clk);
  dff _89418_ (\oc8051_gm_cxrom_1.cell9.data [4], _05583_, clk);
  dff _89419_ (\oc8051_gm_cxrom_1.cell9.data [5], _05587_, clk);
  dff _89420_ (\oc8051_gm_cxrom_1.cell9.data [6], _05590_, clk);
  dff _89421_ (\oc8051_gm_cxrom_1.cell9.data [7], _05560_, clk);
  dff _89422_ (\oc8051_gm_cxrom_1.cell9.valid , _05563_, clk);
  dff _89423_ (\oc8051_golden_model_1.IRAM[15] [0], _41724_, clk);
  dff _89424_ (\oc8051_golden_model_1.IRAM[15] [1], _41725_, clk);
  dff _89425_ (\oc8051_golden_model_1.IRAM[15] [2], _41726_, clk);
  dff _89426_ (\oc8051_golden_model_1.IRAM[15] [3], _41728_, clk);
  dff _89427_ (\oc8051_golden_model_1.IRAM[15] [4], _41729_, clk);
  dff _89428_ (\oc8051_golden_model_1.IRAM[15] [5], _41730_, clk);
  dff _89429_ (\oc8051_golden_model_1.IRAM[15] [6], _41731_, clk);
  dff _89430_ (\oc8051_golden_model_1.IRAM[15] [7], _41495_, clk);
  dff _89431_ (\oc8051_golden_model_1.IRAM[14] [0], _41712_, clk);
  dff _89432_ (\oc8051_golden_model_1.IRAM[14] [1], _41713_, clk);
  dff _89433_ (\oc8051_golden_model_1.IRAM[14] [2], _41714_, clk);
  dff _89434_ (\oc8051_golden_model_1.IRAM[14] [3], _41716_, clk);
  dff _89435_ (\oc8051_golden_model_1.IRAM[14] [4], _41717_, clk);
  dff _89436_ (\oc8051_golden_model_1.IRAM[14] [5], _41718_, clk);
  dff _89437_ (\oc8051_golden_model_1.IRAM[14] [6], _41719_, clk);
  dff _89438_ (\oc8051_golden_model_1.IRAM[14] [7], _41720_, clk);
  dff _89439_ (\oc8051_golden_model_1.IRAM[13] [0], _41700_, clk);
  dff _89440_ (\oc8051_golden_model_1.IRAM[13] [1], _41701_, clk);
  dff _89441_ (\oc8051_golden_model_1.IRAM[13] [2], _41702_, clk);
  dff _89442_ (\oc8051_golden_model_1.IRAM[13] [3], _41703_, clk);
  dff _89443_ (\oc8051_golden_model_1.IRAM[13] [4], _41705_, clk);
  dff _89444_ (\oc8051_golden_model_1.IRAM[13] [5], _41706_, clk);
  dff _89445_ (\oc8051_golden_model_1.IRAM[13] [6], _41707_, clk);
  dff _89446_ (\oc8051_golden_model_1.IRAM[13] [7], _41708_, clk);
  dff _89447_ (\oc8051_golden_model_1.IRAM[12] [0], _41689_, clk);
  dff _89448_ (\oc8051_golden_model_1.IRAM[12] [1], _41690_, clk);
  dff _89449_ (\oc8051_golden_model_1.IRAM[12] [2], _41691_, clk);
  dff _89450_ (\oc8051_golden_model_1.IRAM[12] [3], _41692_, clk);
  dff _89451_ (\oc8051_golden_model_1.IRAM[12] [4], _41694_, clk);
  dff _89452_ (\oc8051_golden_model_1.IRAM[12] [5], _41695_, clk);
  dff _89453_ (\oc8051_golden_model_1.IRAM[12] [6], _41696_, clk);
  dff _89454_ (\oc8051_golden_model_1.IRAM[12] [7], _41697_, clk);
  dff _89455_ (\oc8051_golden_model_1.IRAM[11] [0], _41677_, clk);
  dff _89456_ (\oc8051_golden_model_1.IRAM[11] [1], _41679_, clk);
  dff _89457_ (\oc8051_golden_model_1.IRAM[11] [2], _41680_, clk);
  dff _89458_ (\oc8051_golden_model_1.IRAM[11] [3], _41681_, clk);
  dff _89459_ (\oc8051_golden_model_1.IRAM[11] [4], _41682_, clk);
  dff _89460_ (\oc8051_golden_model_1.IRAM[11] [5], _41683_, clk);
  dff _89461_ (\oc8051_golden_model_1.IRAM[11] [6], _41684_, clk);
  dff _89462_ (\oc8051_golden_model_1.IRAM[11] [7], _41685_, clk);
  dff _89463_ (\oc8051_golden_model_1.IRAM[10] [0], _41665_, clk);
  dff _89464_ (\oc8051_golden_model_1.IRAM[10] [1], _41667_, clk);
  dff _89465_ (\oc8051_golden_model_1.IRAM[10] [2], _41668_, clk);
  dff _89466_ (\oc8051_golden_model_1.IRAM[10] [3], _41669_, clk);
  dff _89467_ (\oc8051_golden_model_1.IRAM[10] [4], _41670_, clk);
  dff _89468_ (\oc8051_golden_model_1.IRAM[10] [5], _41671_, clk);
  dff _89469_ (\oc8051_golden_model_1.IRAM[10] [6], _41673_, clk);
  dff _89470_ (\oc8051_golden_model_1.IRAM[10] [7], _41674_, clk);
  dff _89471_ (\oc8051_golden_model_1.IRAM[9] [0], _41652_, clk);
  dff _89472_ (\oc8051_golden_model_1.IRAM[9] [1], _41653_, clk);
  dff _89473_ (\oc8051_golden_model_1.IRAM[9] [2], _41656_, clk);
  dff _89474_ (\oc8051_golden_model_1.IRAM[9] [3], _41657_, clk);
  dff _89475_ (\oc8051_golden_model_1.IRAM[9] [4], _41658_, clk);
  dff _89476_ (\oc8051_golden_model_1.IRAM[9] [5], _41659_, clk);
  dff _89477_ (\oc8051_golden_model_1.IRAM[9] [6], _41660_, clk);
  dff _89478_ (\oc8051_golden_model_1.IRAM[9] [7], _41662_, clk);
  dff _89479_ (\oc8051_golden_model_1.IRAM[8] [0], _41641_, clk);
  dff _89480_ (\oc8051_golden_model_1.IRAM[8] [1], _41642_, clk);
  dff _89481_ (\oc8051_golden_model_1.IRAM[8] [2], _41644_, clk);
  dff _89482_ (\oc8051_golden_model_1.IRAM[8] [3], _41645_, clk);
  dff _89483_ (\oc8051_golden_model_1.IRAM[8] [4], _41646_, clk);
  dff _89484_ (\oc8051_golden_model_1.IRAM[8] [5], _41647_, clk);
  dff _89485_ (\oc8051_golden_model_1.IRAM[8] [6], _41648_, clk);
  dff _89486_ (\oc8051_golden_model_1.IRAM[8] [7], _41649_, clk);
  dff _89487_ (\oc8051_golden_model_1.IRAM[7] [0], _41628_, clk);
  dff _89488_ (\oc8051_golden_model_1.IRAM[7] [1], _41630_, clk);
  dff _89489_ (\oc8051_golden_model_1.IRAM[7] [2], _41631_, clk);
  dff _89490_ (\oc8051_golden_model_1.IRAM[7] [3], _41632_, clk);
  dff _89491_ (\oc8051_golden_model_1.IRAM[7] [4], _41633_, clk);
  dff _89492_ (\oc8051_golden_model_1.IRAM[7] [5], _41634_, clk);
  dff _89493_ (\oc8051_golden_model_1.IRAM[7] [6], _41636_, clk);
  dff _89494_ (\oc8051_golden_model_1.IRAM[7] [7], _41637_, clk);
  dff _89495_ (\oc8051_golden_model_1.IRAM[6] [0], _41616_, clk);
  dff _89496_ (\oc8051_golden_model_1.IRAM[6] [1], _41618_, clk);
  dff _89497_ (\oc8051_golden_model_1.IRAM[6] [2], _41619_, clk);
  dff _89498_ (\oc8051_golden_model_1.IRAM[6] [3], _41620_, clk);
  dff _89499_ (\oc8051_golden_model_1.IRAM[6] [4], _41621_, clk);
  dff _89500_ (\oc8051_golden_model_1.IRAM[6] [5], _41622_, clk);
  dff _89501_ (\oc8051_golden_model_1.IRAM[6] [6], _41624_, clk);
  dff _89502_ (\oc8051_golden_model_1.IRAM[6] [7], _41625_, clk);
  dff _89503_ (\oc8051_golden_model_1.IRAM[5] [0], _41604_, clk);
  dff _89504_ (\oc8051_golden_model_1.IRAM[5] [1], _41605_, clk);
  dff _89505_ (\oc8051_golden_model_1.IRAM[5] [2], _41607_, clk);
  dff _89506_ (\oc8051_golden_model_1.IRAM[5] [3], _41608_, clk);
  dff _89507_ (\oc8051_golden_model_1.IRAM[5] [4], _41609_, clk);
  dff _89508_ (\oc8051_golden_model_1.IRAM[5] [5], _41610_, clk);
  dff _89509_ (\oc8051_golden_model_1.IRAM[5] [6], _41611_, clk);
  dff _89510_ (\oc8051_golden_model_1.IRAM[5] [7], _41613_, clk);
  dff _89511_ (\oc8051_golden_model_1.IRAM[4] [0], _41592_, clk);
  dff _89512_ (\oc8051_golden_model_1.IRAM[4] [1], _41593_, clk);
  dff _89513_ (\oc8051_golden_model_1.IRAM[4] [2], _41594_, clk);
  dff _89514_ (\oc8051_golden_model_1.IRAM[4] [3], _41595_, clk);
  dff _89515_ (\oc8051_golden_model_1.IRAM[4] [4], _41596_, clk);
  dff _89516_ (\oc8051_golden_model_1.IRAM[4] [5], _41597_, clk);
  dff _89517_ (\oc8051_golden_model_1.IRAM[4] [6], _41598_, clk);
  dff _89518_ (\oc8051_golden_model_1.IRAM[4] [7], _41601_, clk);
  dff _89519_ (\oc8051_golden_model_1.IRAM[3] [0], _41579_, clk);
  dff _89520_ (\oc8051_golden_model_1.IRAM[3] [1], _41581_, clk);
  dff _89521_ (\oc8051_golden_model_1.IRAM[3] [2], _41582_, clk);
  dff _89522_ (\oc8051_golden_model_1.IRAM[3] [3], _41583_, clk);
  dff _89523_ (\oc8051_golden_model_1.IRAM[3] [4], _41584_, clk);
  dff _89524_ (\oc8051_golden_model_1.IRAM[3] [5], _41585_, clk);
  dff _89525_ (\oc8051_golden_model_1.IRAM[3] [6], _41587_, clk);
  dff _89526_ (\oc8051_golden_model_1.IRAM[3] [7], _41588_, clk);
  dff _89527_ (\oc8051_golden_model_1.IRAM[2] [0], _41567_, clk);
  dff _89528_ (\oc8051_golden_model_1.IRAM[2] [1], _41568_, clk);
  dff _89529_ (\oc8051_golden_model_1.IRAM[2] [2], _41570_, clk);
  dff _89530_ (\oc8051_golden_model_1.IRAM[2] [3], _41571_, clk);
  dff _89531_ (\oc8051_golden_model_1.IRAM[2] [4], _41572_, clk);
  dff _89532_ (\oc8051_golden_model_1.IRAM[2] [5], _41573_, clk);
  dff _89533_ (\oc8051_golden_model_1.IRAM[2] [6], _41574_, clk);
  dff _89534_ (\oc8051_golden_model_1.IRAM[2] [7], _41576_, clk);
  dff _89535_ (\oc8051_golden_model_1.IRAM[1] [0], _41554_, clk);
  dff _89536_ (\oc8051_golden_model_1.IRAM[1] [1], _41556_, clk);
  dff _89537_ (\oc8051_golden_model_1.IRAM[1] [2], _41557_, clk);
  dff _89538_ (\oc8051_golden_model_1.IRAM[1] [3], _41558_, clk);
  dff _89539_ (\oc8051_golden_model_1.IRAM[1] [4], _41559_, clk);
  dff _89540_ (\oc8051_golden_model_1.IRAM[1] [5], _41560_, clk);
  dff _89541_ (\oc8051_golden_model_1.IRAM[1] [6], _41562_, clk);
  dff _89542_ (\oc8051_golden_model_1.IRAM[1] [7], _41563_, clk);
  dff _89543_ (\oc8051_golden_model_1.IRAM[0] [0], _41541_, clk);
  dff _89544_ (\oc8051_golden_model_1.IRAM[0] [1], _41542_, clk);
  dff _89545_ (\oc8051_golden_model_1.IRAM[0] [2], _41543_, clk);
  dff _89546_ (\oc8051_golden_model_1.IRAM[0] [3], _41545_, clk);
  dff _89547_ (\oc8051_golden_model_1.IRAM[0] [4], _41546_, clk);
  dff _89548_ (\oc8051_golden_model_1.IRAM[0] [5], _41548_, clk);
  dff _89549_ (\oc8051_golden_model_1.IRAM[0] [6], _41549_, clk);
  dff _89550_ (\oc8051_golden_model_1.IRAM[0] [7], _41550_, clk);
  dff _89551_ (\oc8051_golden_model_1.B [0], _44115_, clk);
  dff _89552_ (\oc8051_golden_model_1.B [1], _44116_, clk);
  dff _89553_ (\oc8051_golden_model_1.B [2], _44117_, clk);
  dff _89554_ (\oc8051_golden_model_1.B [3], _44118_, clk);
  dff _89555_ (\oc8051_golden_model_1.B [4], _44119_, clk);
  dff _89556_ (\oc8051_golden_model_1.B [5], _44121_, clk);
  dff _89557_ (\oc8051_golden_model_1.B [6], _44122_, clk);
  dff _89558_ (\oc8051_golden_model_1.B [7], _41496_, clk);
  dff _89559_ (\oc8051_golden_model_1.ACC [0], _44123_, clk);
  dff _89560_ (\oc8051_golden_model_1.ACC [1], _44125_, clk);
  dff _89561_ (\oc8051_golden_model_1.ACC [2], _44126_, clk);
  dff _89562_ (\oc8051_golden_model_1.ACC [3], _44127_, clk);
  dff _89563_ (\oc8051_golden_model_1.ACC [4], _44128_, clk);
  dff _89564_ (\oc8051_golden_model_1.ACC [5], _44129_, clk);
  dff _89565_ (\oc8051_golden_model_1.ACC [6], _44130_, clk);
  dff _89566_ (\oc8051_golden_model_1.ACC [7], _41497_, clk);
  dff _89567_ (\oc8051_golden_model_1.PCON [0], _44132_, clk);
  dff _89568_ (\oc8051_golden_model_1.PCON [1], _44133_, clk);
  dff _89569_ (\oc8051_golden_model_1.PCON [2], _44134_, clk);
  dff _89570_ (\oc8051_golden_model_1.PCON [3], _44135_, clk);
  dff _89571_ (\oc8051_golden_model_1.PCON [4], _44136_, clk);
  dff _89572_ (\oc8051_golden_model_1.PCON [5], _44137_, clk);
  dff _89573_ (\oc8051_golden_model_1.PCON [6], _44138_, clk);
  dff _89574_ (\oc8051_golden_model_1.PCON [7], _41498_, clk);
  dff _89575_ (\oc8051_golden_model_1.TMOD [0], _44140_, clk);
  dff _89576_ (\oc8051_golden_model_1.TMOD [1], _44141_, clk);
  dff _89577_ (\oc8051_golden_model_1.TMOD [2], _44142_, clk);
  dff _89578_ (\oc8051_golden_model_1.TMOD [3], _44144_, clk);
  dff _89579_ (\oc8051_golden_model_1.TMOD [4], _44145_, clk);
  dff _89580_ (\oc8051_golden_model_1.TMOD [5], _44146_, clk);
  dff _89581_ (\oc8051_golden_model_1.TMOD [6], _44147_, clk);
  dff _89582_ (\oc8051_golden_model_1.TMOD [7], _41499_, clk);
  dff _89583_ (\oc8051_golden_model_1.DPL [0], _44149_, clk);
  dff _89584_ (\oc8051_golden_model_1.DPL [1], _44150_, clk);
  dff _89585_ (\oc8051_golden_model_1.DPL [2], _44151_, clk);
  dff _89586_ (\oc8051_golden_model_1.DPL [3], _44152_, clk);
  dff _89587_ (\oc8051_golden_model_1.DPL [4], _44153_, clk);
  dff _89588_ (\oc8051_golden_model_1.DPL [5], _44154_, clk);
  dff _89589_ (\oc8051_golden_model_1.DPL [6], _44155_, clk);
  dff _89590_ (\oc8051_golden_model_1.DPL [7], _41501_, clk);
  dff _89591_ (\oc8051_golden_model_1.DPH [0], _44157_, clk);
  dff _89592_ (\oc8051_golden_model_1.DPH [1], _44158_, clk);
  dff _89593_ (\oc8051_golden_model_1.DPH [2], _44159_, clk);
  dff _89594_ (\oc8051_golden_model_1.DPH [3], _44160_, clk);
  dff _89595_ (\oc8051_golden_model_1.DPH [4], _44161_, clk);
  dff _89596_ (\oc8051_golden_model_1.DPH [5], _44162_, clk);
  dff _89597_ (\oc8051_golden_model_1.DPH [6], _44163_, clk);
  dff _89598_ (\oc8051_golden_model_1.DPH [7], _41502_, clk);
  dff _89599_ (\oc8051_golden_model_1.TL1 [0], _44164_, clk);
  dff _89600_ (\oc8051_golden_model_1.TL1 [1], _44166_, clk);
  dff _89601_ (\oc8051_golden_model_1.TL1 [2], _44167_, clk);
  dff _89602_ (\oc8051_golden_model_1.TL1 [3], _44168_, clk);
  dff _89603_ (\oc8051_golden_model_1.TL1 [4], _44169_, clk);
  dff _89604_ (\oc8051_golden_model_1.TL1 [5], _44170_, clk);
  dff _89605_ (\oc8051_golden_model_1.TL1 [6], _44171_, clk);
  dff _89606_ (\oc8051_golden_model_1.TL1 [7], _41503_, clk);
  dff _89607_ (\oc8051_golden_model_1.TL0 [0], _44172_, clk);
  dff _89608_ (\oc8051_golden_model_1.TL0 [1], _44173_, clk);
  dff _89609_ (\oc8051_golden_model_1.TL0 [2], _44174_, clk);
  dff _89610_ (\oc8051_golden_model_1.TL0 [3], _44175_, clk);
  dff _89611_ (\oc8051_golden_model_1.TL0 [4], _44176_, clk);
  dff _89612_ (\oc8051_golden_model_1.TL0 [5], _44177_, clk);
  dff _89613_ (\oc8051_golden_model_1.TL0 [6], _44178_, clk);
  dff _89614_ (\oc8051_golden_model_1.TL0 [7], _41504_, clk);
  dff _89615_ (\oc8051_golden_model_1.TCON [0], _44180_, clk);
  dff _89616_ (\oc8051_golden_model_1.TCON [1], _44181_, clk);
  dff _89617_ (\oc8051_golden_model_1.TCON [2], _44182_, clk);
  dff _89618_ (\oc8051_golden_model_1.TCON [3], _44184_, clk);
  dff _89619_ (\oc8051_golden_model_1.TCON [4], _44185_, clk);
  dff _89620_ (\oc8051_golden_model_1.TCON [5], _44186_, clk);
  dff _89621_ (\oc8051_golden_model_1.TCON [6], _44187_, clk);
  dff _89622_ (\oc8051_golden_model_1.TCON [7], _41505_, clk);
  dff _89623_ (\oc8051_golden_model_1.TH1 [0], _44189_, clk);
  dff _89624_ (\oc8051_golden_model_1.TH1 [1], _44190_, clk);
  dff _89625_ (\oc8051_golden_model_1.TH1 [2], _44191_, clk);
  dff _89626_ (\oc8051_golden_model_1.TH1 [3], _44192_, clk);
  dff _89627_ (\oc8051_golden_model_1.TH1 [4], _44193_, clk);
  dff _89628_ (\oc8051_golden_model_1.TH1 [5], _44194_, clk);
  dff _89629_ (\oc8051_golden_model_1.TH1 [6], _44195_, clk);
  dff _89630_ (\oc8051_golden_model_1.TH1 [7], _41507_, clk);
  dff _89631_ (\oc8051_golden_model_1.TH0 [0], _44197_, clk);
  dff _89632_ (\oc8051_golden_model_1.TH0 [1], _44198_, clk);
  dff _89633_ (\oc8051_golden_model_1.TH0 [2], _44199_, clk);
  dff _89634_ (\oc8051_golden_model_1.TH0 [3], _44200_, clk);
  dff _89635_ (\oc8051_golden_model_1.TH0 [4], _44201_, clk);
  dff _89636_ (\oc8051_golden_model_1.TH0 [5], _44203_, clk);
  dff _89637_ (\oc8051_golden_model_1.TH0 [6], _44204_, clk);
  dff _89638_ (\oc8051_golden_model_1.TH0 [7], _41508_, clk);
  dff _89639_ (\oc8051_golden_model_1.PC [0], _44206_, clk);
  dff _89640_ (\oc8051_golden_model_1.PC [1], _44207_, clk);
  dff _89641_ (\oc8051_golden_model_1.PC [2], _44208_, clk);
  dff _89642_ (\oc8051_golden_model_1.PC [3], _44210_, clk);
  dff _89643_ (\oc8051_golden_model_1.PC [4], _44211_, clk);
  dff _89644_ (\oc8051_golden_model_1.PC [5], _44212_, clk);
  dff _89645_ (\oc8051_golden_model_1.PC [6], _44213_, clk);
  dff _89646_ (\oc8051_golden_model_1.PC [7], _44214_, clk);
  dff _89647_ (\oc8051_golden_model_1.PC [8], _44215_, clk);
  dff _89648_ (\oc8051_golden_model_1.PC [9], _44216_, clk);
  dff _89649_ (\oc8051_golden_model_1.PC [10], _44217_, clk);
  dff _89650_ (\oc8051_golden_model_1.PC [11], _44218_, clk);
  dff _89651_ (\oc8051_golden_model_1.PC [12], _44219_, clk);
  dff _89652_ (\oc8051_golden_model_1.PC [13], _44221_, clk);
  dff _89653_ (\oc8051_golden_model_1.PC [14], _44222_, clk);
  dff _89654_ (\oc8051_golden_model_1.PC [15], _41509_, clk);
  dff _89655_ (\oc8051_golden_model_1.P2 [0], _44223_, clk);
  dff _89656_ (\oc8051_golden_model_1.P2 [1], _44225_, clk);
  dff _89657_ (\oc8051_golden_model_1.P2 [2], _44226_, clk);
  dff _89658_ (\oc8051_golden_model_1.P2 [3], _44227_, clk);
  dff _89659_ (\oc8051_golden_model_1.P2 [4], _44228_, clk);
  dff _89660_ (\oc8051_golden_model_1.P2 [5], _44229_, clk);
  dff _89661_ (\oc8051_golden_model_1.P2 [6], _44230_, clk);
  dff _89662_ (\oc8051_golden_model_1.P2 [7], _41510_, clk);
  dff _89663_ (\oc8051_golden_model_1.P3 [0], _44232_, clk);
  dff _89664_ (\oc8051_golden_model_1.P3 [1], _44233_, clk);
  dff _89665_ (\oc8051_golden_model_1.P3 [2], _44234_, clk);
  dff _89666_ (\oc8051_golden_model_1.P3 [3], _44235_, clk);
  dff _89667_ (\oc8051_golden_model_1.P3 [4], _44236_, clk);
  dff _89668_ (\oc8051_golden_model_1.P3 [5], _44237_, clk);
  dff _89669_ (\oc8051_golden_model_1.P3 [6], _44238_, clk);
  dff _89670_ (\oc8051_golden_model_1.P3 [7], _41511_, clk);
  dff _89671_ (\oc8051_golden_model_1.P0 [0], _44240_, clk);
  dff _89672_ (\oc8051_golden_model_1.P0 [1], _44241_, clk);
  dff _89673_ (\oc8051_golden_model_1.P0 [2], _44242_, clk);
  dff _89674_ (\oc8051_golden_model_1.P0 [3], _44244_, clk);
  dff _89675_ (\oc8051_golden_model_1.P0 [4], _44245_, clk);
  dff _89676_ (\oc8051_golden_model_1.P0 [5], _44246_, clk);
  dff _89677_ (\oc8051_golden_model_1.P0 [6], _44247_, clk);
  dff _89678_ (\oc8051_golden_model_1.P0 [7], _41513_, clk);
  dff _89679_ (\oc8051_golden_model_1.P1 [0], _44249_, clk);
  dff _89680_ (\oc8051_golden_model_1.P1 [1], _44250_, clk);
  dff _89681_ (\oc8051_golden_model_1.P1 [2], _44251_, clk);
  dff _89682_ (\oc8051_golden_model_1.P1 [3], _44252_, clk);
  dff _89683_ (\oc8051_golden_model_1.P1 [4], _44253_, clk);
  dff _89684_ (\oc8051_golden_model_1.P1 [5], _44254_, clk);
  dff _89685_ (\oc8051_golden_model_1.P1 [6], _44255_, clk);
  dff _89686_ (\oc8051_golden_model_1.P1 [7], _41514_, clk);
  dff _89687_ (\oc8051_golden_model_1.IP [0], _44257_, clk);
  dff _89688_ (\oc8051_golden_model_1.IP [1], _44258_, clk);
  dff _89689_ (\oc8051_golden_model_1.IP [2], _44259_, clk);
  dff _89690_ (\oc8051_golden_model_1.IP [3], _44260_, clk);
  dff _89691_ (\oc8051_golden_model_1.IP [4], _44261_, clk);
  dff _89692_ (\oc8051_golden_model_1.IP [5], _44263_, clk);
  dff _89693_ (\oc8051_golden_model_1.IP [6], _44264_, clk);
  dff _89694_ (\oc8051_golden_model_1.IP [7], _41515_, clk);
  dff _89695_ (\oc8051_golden_model_1.IE [0], _44265_, clk);
  dff _89696_ (\oc8051_golden_model_1.IE [1], _44267_, clk);
  dff _89697_ (\oc8051_golden_model_1.IE [2], _44268_, clk);
  dff _89698_ (\oc8051_golden_model_1.IE [3], _44269_, clk);
  dff _89699_ (\oc8051_golden_model_1.IE [4], _44270_, clk);
  dff _89700_ (\oc8051_golden_model_1.IE [5], _44271_, clk);
  dff _89701_ (\oc8051_golden_model_1.IE [6], _44272_, clk);
  dff _89702_ (\oc8051_golden_model_1.IE [7], _41516_, clk);
  dff _89703_ (\oc8051_golden_model_1.SCON [0], _44274_, clk);
  dff _89704_ (\oc8051_golden_model_1.SCON [1], _44275_, clk);
  dff _89705_ (\oc8051_golden_model_1.SCON [2], _44276_, clk);
  dff _89706_ (\oc8051_golden_model_1.SCON [3], _44277_, clk);
  dff _89707_ (\oc8051_golden_model_1.SCON [4], _44278_, clk);
  dff _89708_ (\oc8051_golden_model_1.SCON [5], _44279_, clk);
  dff _89709_ (\oc8051_golden_model_1.SCON [6], _44280_, clk);
  dff _89710_ (\oc8051_golden_model_1.SCON [7], _41517_, clk);
  dff _89711_ (\oc8051_golden_model_1.SP [0], _44282_, clk);
  dff _89712_ (\oc8051_golden_model_1.SP [1], _44283_, clk);
  dff _89713_ (\oc8051_golden_model_1.SP [2], _44284_, clk);
  dff _89714_ (\oc8051_golden_model_1.SP [3], _44286_, clk);
  dff _89715_ (\oc8051_golden_model_1.SP [4], _44287_, clk);
  dff _89716_ (\oc8051_golden_model_1.SP [5], _44288_, clk);
  dff _89717_ (\oc8051_golden_model_1.SP [6], _44289_, clk);
  dff _89718_ (\oc8051_golden_model_1.SP [7], _41519_, clk);
  dff _89719_ (\oc8051_golden_model_1.SBUF [0], _44291_, clk);
  dff _89720_ (\oc8051_golden_model_1.SBUF [1], _44292_, clk);
  dff _89721_ (\oc8051_golden_model_1.SBUF [2], _44293_, clk);
  dff _89722_ (\oc8051_golden_model_1.SBUF [3], _44294_, clk);
  dff _89723_ (\oc8051_golden_model_1.SBUF [4], _44295_, clk);
  dff _89724_ (\oc8051_golden_model_1.SBUF [5], _44296_, clk);
  dff _89725_ (\oc8051_golden_model_1.SBUF [6], _44297_, clk);
  dff _89726_ (\oc8051_golden_model_1.SBUF [7], _41520_, clk);
  dff _89727_ (\oc8051_golden_model_1.PSW [0], _44299_, clk);
  dff _89728_ (\oc8051_golden_model_1.PSW [1], _44300_, clk);
  dff _89729_ (\oc8051_golden_model_1.PSW [2], _44301_, clk);
  dff _89730_ (\oc8051_golden_model_1.PSW [3], _44302_, clk);
  dff _89731_ (\oc8051_golden_model_1.PSW [4], _44303_, clk);
  dff _89732_ (\oc8051_golden_model_1.PSW [5], _44305_, clk);
  dff _89733_ (\oc8051_golden_model_1.PSW [6], _44306_, clk);
  dff _89734_ (\oc8051_golden_model_1.PSW [7], _41521_, clk);
  dff _89735_ (\oc8051_golden_model_1.P0INREG [0], _44307_, clk);
  dff _89736_ (\oc8051_golden_model_1.P0INREG [1], _44309_, clk);
  dff _89737_ (\oc8051_golden_model_1.P0INREG [2], _44310_, clk);
  dff _89738_ (\oc8051_golden_model_1.P0INREG [3], _44311_, clk);
  dff _89739_ (\oc8051_golden_model_1.P0INREG [4], _44312_, clk);
  dff _89740_ (\oc8051_golden_model_1.P0INREG [5], _44313_, clk);
  dff _89741_ (\oc8051_golden_model_1.P0INREG [6], _44314_, clk);
  dff _89742_ (\oc8051_golden_model_1.P0INREG [7], _41522_, clk);
  dff _89743_ (\oc8051_golden_model_1.P1INREG [0], _44316_, clk);
  dff _89744_ (\oc8051_golden_model_1.P1INREG [1], _44317_, clk);
  dff _89745_ (\oc8051_golden_model_1.P1INREG [2], _44318_, clk);
  dff _89746_ (\oc8051_golden_model_1.P1INREG [3], _44319_, clk);
  dff _89747_ (\oc8051_golden_model_1.P1INREG [4], _44320_, clk);
  dff _89748_ (\oc8051_golden_model_1.P1INREG [5], _44321_, clk);
  dff _89749_ (\oc8051_golden_model_1.P1INREG [6], _44322_, clk);
  dff _89750_ (\oc8051_golden_model_1.P1INREG [7], _41523_, clk);
  dff _89751_ (\oc8051_golden_model_1.P2INREG [0], _44324_, clk);
  dff _89752_ (\oc8051_golden_model_1.P2INREG [1], _44325_, clk);
  dff _89753_ (\oc8051_golden_model_1.P2INREG [2], _44326_, clk);
  dff _89754_ (\oc8051_golden_model_1.P2INREG [3], _44328_, clk);
  dff _89755_ (\oc8051_golden_model_1.P2INREG [4], _44329_, clk);
  dff _89756_ (\oc8051_golden_model_1.P2INREG [5], _44330_, clk);
  dff _89757_ (\oc8051_golden_model_1.P2INREG [6], _44331_, clk);
  dff _89758_ (\oc8051_golden_model_1.P2INREG [7], _41525_, clk);
  dff _89759_ (\oc8051_golden_model_1.P3INREG [0], _44333_, clk);
  dff _89760_ (\oc8051_golden_model_1.P3INREG [1], _44334_, clk);
  dff _89761_ (\oc8051_golden_model_1.P3INREG [2], _44335_, clk);
  dff _89762_ (\oc8051_golden_model_1.P3INREG [3], _44336_, clk);
  dff _89763_ (\oc8051_golden_model_1.P3INREG [4], _44337_, clk);
  dff _89764_ (\oc8051_golden_model_1.P3INREG [5], _44338_, clk);
  dff _89765_ (\oc8051_golden_model_1.P3INREG [6], _44339_, clk);
  dff _89766_ (\oc8051_golden_model_1.P3INREG [7], _41526_, clk);
  dff _89767_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02847_, clk);
  dff _89768_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02859_, clk);
  dff _89769_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02881_, clk);
  dff _89770_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02906_, clk);
  dff _89771_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02931_, clk);
  dff _89772_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00956_, clk);
  dff _89773_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02942_, clk);
  dff _89774_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00926_, clk);
  dff _89775_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02955_, clk);
  dff _89776_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02968_, clk);
  dff _89777_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02980_, clk);
  dff _89778_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02992_, clk);
  dff _89779_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03005_, clk);
  dff _89780_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03016_, clk);
  dff _89781_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03029_, clk);
  dff _89782_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00976_, clk);
  dff _89783_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02349_, clk);
  dff _89784_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22076_, clk);
  dff _89785_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02541_, clk);
  dff _89786_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02720_, clk);
  dff _89787_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02893_, clk);
  dff _89788_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03129_, clk);
  dff _89789_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03347_, clk);
  dff _89790_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03548_, clk);
  dff _89791_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03749_, clk);
  dff _89792_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03948_, clk);
  dff _89793_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04045_, clk);
  dff _89794_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04144_, clk);
  dff _89795_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04243_, clk);
  dff _89796_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04343_, clk);
  dff _89797_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04436_, clk);
  dff _89798_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04536_, clk);
  dff _89799_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04634_, clk);
  dff _89800_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24254_, clk);
  dff _89801_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _39706_, clk);
  dff _89802_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _39708_, clk);
  dff _89803_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _39709_, clk);
  dff _89804_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _39710_, clk);
  dff _89805_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _39711_, clk);
  dff _89806_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _39712_, clk);
  dff _89807_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _39713_, clk);
  dff _89808_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _39695_, clk);
  dff _89809_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _39714_, clk);
  dff _89810_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _39715_, clk);
  dff _89811_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _39717_, clk);
  dff _89812_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _39718_, clk);
  dff _89813_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _39719_, clk);
  dff _89814_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _39720_, clk);
  dff _89815_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _39721_, clk);
  dff _89816_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _39696_, clk);
  dff _89817_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _39722_, clk);
  dff _89818_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _39723_, clk);
  dff _89819_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _39724_, clk);
  dff _89820_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _39725_, clk);
  dff _89821_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _39726_, clk);
  dff _89822_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _39728_, clk);
  dff _89823_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _39729_, clk);
  dff _89824_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _39698_, clk);
  dff _89825_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34139_, clk);
  dff _89826_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34142_, clk);
  dff _89827_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09702_, clk);
  dff _89828_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34144_, clk);
  dff _89829_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34146_, clk);
  dff _89830_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09705_, clk);
  dff _89831_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34148_, clk);
  dff _89832_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09708_, clk);
  dff _89833_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34150_, clk);
  dff _89834_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34152_, clk);
  dff _89835_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34154_, clk);
  dff _89836_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09711_, clk);
  dff _89837_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34156_, clk);
  dff _89838_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09714_, clk);
  dff _89839_ (\oc8051_top_1.oc8051_decoder1.wr , _09717_, clk);
  dff _89840_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09776_, clk);
  dff _89841_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09778_, clk);
  dff _89842_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09681_, clk);
  dff _89843_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09781_, clk);
  dff _89844_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09784_, clk);
  dff _89845_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09684_, clk);
  dff _89846_ (\oc8051_top_1.oc8051_decoder1.state [0], _09787_, clk);
  dff _89847_ (\oc8051_top_1.oc8051_decoder1.state [1], _09687_, clk);
  dff _89848_ (\oc8051_top_1.oc8051_decoder1.op [0], _09790_, clk);
  dff _89849_ (\oc8051_top_1.oc8051_decoder1.op [1], _09793_, clk);
  dff _89850_ (\oc8051_top_1.oc8051_decoder1.op [2], _09796_, clk);
  dff _89851_ (\oc8051_top_1.oc8051_decoder1.op [3], _09799_, clk);
  dff _89852_ (\oc8051_top_1.oc8051_decoder1.op [4], _09802_, clk);
  dff _89853_ (\oc8051_top_1.oc8051_decoder1.op [5], _09805_, clk);
  dff _89854_ (\oc8051_top_1.oc8051_decoder1.op [6], _09808_, clk);
  dff _89855_ (\oc8051_top_1.oc8051_decoder1.op [7], _09690_, clk);
  dff _89856_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09693_, clk);
  dff _89857_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34137_, clk);
  dff _89858_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09699_, clk);
  dff _89859_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09811_, clk);
  dff _89860_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09696_, clk);
  dff _89861_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _40499_, clk);
  dff _89862_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _40531_, clk);
  dff _89863_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _40532_, clk);
  dff _89864_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _40533_, clk);
  dff _89865_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _40534_, clk);
  dff _89866_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _40535_, clk);
  dff _89867_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _40536_, clk);
  dff _89868_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _40537_, clk);
  dff _89869_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _40500_, clk);
  dff _89870_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _40539_, clk);
  dff _89871_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _40540_, clk);
  dff _89872_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _40541_, clk);
  dff _89873_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _40542_, clk);
  dff _89874_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _40543_, clk);
  dff _89875_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _40544_, clk);
  dff _89876_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _40545_, clk);
  dff _89877_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _40501_, clk);
  dff _89878_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _40546_, clk);
  dff _89879_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _40547_, clk);
  dff _89880_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _40548_, clk);
  dff _89881_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _40550_, clk);
  dff _89882_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _40551_, clk);
  dff _89883_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _40552_, clk);
  dff _89884_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _40553_, clk);
  dff _89885_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _40502_, clk);
  dff _89886_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _40554_, clk);
  dff _89887_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _40555_, clk);
  dff _89888_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _40556_, clk);
  dff _89889_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _40557_, clk);
  dff _89890_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _40558_, clk);
  dff _89891_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _40559_, clk);
  dff _89892_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _40561_, clk);
  dff _89893_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _40504_, clk);
  dff _89894_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _40076_, clk);
  dff _89895_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _40077_, clk);
  dff _89896_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _40078_, clk);
  dff _89897_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _40079_, clk);
  dff _89898_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39791_, clk);
  dff _89899_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39863_, clk);
  dff _89900_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39864_, clk);
  dff _89901_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39865_, clk);
  dff _89902_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39866_, clk);
  dff _89903_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39867_, clk);
  dff _89904_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39869_, clk);
  dff _89905_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39870_, clk);
  dff _89906_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39871_, clk);
  dff _89907_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39872_, clk);
  dff _89908_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39873_, clk);
  dff _89909_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39874_, clk);
  dff _89910_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39875_, clk);
  dff _89911_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39876_, clk);
  dff _89912_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39877_, clk);
  dff _89913_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39878_, clk);
  dff _89914_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39751_, clk);
  dff _89915_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39883_, clk);
  dff _89916_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39884_, clk);
  dff _89917_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39885_, clk);
  dff _89918_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39886_, clk);
  dff _89919_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39887_, clk);
  dff _89920_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39888_, clk);
  dff _89921_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39889_, clk);
  dff _89922_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39890_, clk);
  dff _89923_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39891_, clk);
  dff _89924_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39892_, clk);
  dff _89925_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39894_, clk);
  dff _89926_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39895_, clk);
  dff _89927_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39896_, clk);
  dff _89928_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39897_, clk);
  dff _89929_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39898_, clk);
  dff _89930_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39752_, clk);
  dff _89931_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _40080_, clk);
  dff _89932_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _40081_, clk);
  dff _89933_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _40082_, clk);
  dff _89934_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _40083_, clk);
  dff _89935_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _40084_, clk);
  dff _89936_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _40085_, clk);
  dff _89937_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _40086_, clk);
  dff _89938_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _40087_, clk);
  dff _89939_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _40088_, clk);
  dff _89940_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _40089_, clk);
  dff _89941_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _40090_, clk);
  dff _89942_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _40091_, clk);
  dff _89943_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _40092_, clk);
  dff _89944_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _40093_, clk);
  dff _89945_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _40095_, clk);
  dff _89946_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _40096_, clk);
  dff _89947_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _40097_, clk);
  dff _89948_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _40098_, clk);
  dff _89949_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _40099_, clk);
  dff _89950_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _40100_, clk);
  dff _89951_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _40101_, clk);
  dff _89952_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _40102_, clk);
  dff _89953_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _40103_, clk);
  dff _89954_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _40104_, clk);
  dff _89955_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _40106_, clk);
  dff _89956_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _40107_, clk);
  dff _89957_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _40108_, clk);
  dff _89958_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _40109_, clk);
  dff _89959_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _40110_, clk);
  dff _89960_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _40111_, clk);
  dff _89961_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _40112_, clk);
  dff _89962_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39816_, clk);
  dff _89963_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39789_, clk);
  dff _89964_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _89965_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _40113_, clk);
  dff _89966_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _40115_, clk);
  dff _89967_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _40116_, clk);
  dff _89968_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _40117_, clk);
  dff _89969_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _40118_, clk);
  dff _89970_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _40119_, clk);
  dff _89971_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _40121_, clk);
  dff _89972_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39792_, clk);
  dff _89973_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _40122_, clk);
  dff _89974_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _40123_, clk);
  dff _89975_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _40124_, clk);
  dff _89976_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _40125_, clk);
  dff _89977_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _40126_, clk);
  dff _89978_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _40127_, clk);
  dff _89979_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _40128_, clk);
  dff _89980_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39793_, clk);
  dff _89981_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _40129_, clk);
  dff _89982_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _40130_, clk);
  dff _89983_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _40132_, clk);
  dff _89984_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _40133_, clk);
  dff _89985_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _40134_, clk);
  dff _89986_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _40135_, clk);
  dff _89987_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _40136_, clk);
  dff _89988_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39795_, clk);
  dff _89989_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39796_, clk);
  dff _89990_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39797_, clk);
  dff _89991_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _40137_, clk);
  dff _89992_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _40138_, clk);
  dff _89993_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _40139_, clk);
  dff _89994_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _40140_, clk);
  dff _89995_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _40141_, clk);
  dff _89996_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _40143_, clk);
  dff _89997_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _40144_, clk);
  dff _89998_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39798_, clk);
  dff _89999_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _40145_, clk);
  dff _90000_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _40146_, clk);
  dff _90001_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _40147_, clk);
  dff _90002_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _40148_, clk);
  dff _90003_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _40149_, clk);
  dff _90004_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _40150_, clk);
  dff _90005_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _40151_, clk);
  dff _90006_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _40152_, clk);
  dff _90007_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _40154_, clk);
  dff _90008_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _40155_, clk);
  dff _90009_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _40156_, clk);
  dff _90010_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _40157_, clk);
  dff _90011_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _40158_, clk);
  dff _90012_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _40159_, clk);
  dff _90013_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _40160_, clk);
  dff _90014_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39799_, clk);
  dff _90015_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _40161_, clk);
  dff _90016_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _40162_, clk);
  dff _90017_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _40163_, clk);
  dff _90018_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _40165_, clk);
  dff _90019_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _40166_, clk);
  dff _90020_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _40167_, clk);
  dff _90021_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _40168_, clk);
  dff _90022_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _40169_, clk);
  dff _90023_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _40170_, clk);
  dff _90024_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _40171_, clk);
  dff _90025_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _40172_, clk);
  dff _90026_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _40173_, clk);
  dff _90027_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _40174_, clk);
  dff _90028_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _40176_, clk);
  dff _90029_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _40177_, clk);
  dff _90030_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39801_, clk);
  dff _90031_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39802_, clk);
  dff _90032_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39804_, clk);
  dff _90033_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39803_, clk);
  dff _90034_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _40178_, clk);
  dff _90035_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _40179_, clk);
  dff _90036_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _40180_, clk);
  dff _90037_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _40181_, clk);
  dff _90038_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _40182_, clk);
  dff _90039_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _40183_, clk);
  dff _90040_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _40184_, clk);
  dff _90041_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39806_, clk);
  dff _90042_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _40185_, clk);
  dff _90043_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _40187_, clk);
  dff _90044_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39807_, clk);
  dff _90045_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _40188_, clk);
  dff _90046_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _40189_, clk);
  dff _90047_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _40190_, clk);
  dff _90048_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _40191_, clk);
  dff _90049_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _40192_, clk);
  dff _90050_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _40193_, clk);
  dff _90051_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _40194_, clk);
  dff _90052_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39808_, clk);
  dff _90053_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _40195_, clk);
  dff _90054_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _40196_, clk);
  dff _90055_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _40198_, clk);
  dff _90056_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _40199_, clk);
  dff _90057_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _40200_, clk);
  dff _90058_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _40201_, clk);
  dff _90059_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _40202_, clk);
  dff _90060_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39809_, clk);
  dff _90061_ (\oc8051_top_1.oc8051_memory_interface1.reti , _39810_, clk);
  dff _90062_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _40203_, clk);
  dff _90063_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _40204_, clk);
  dff _90064_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _40205_, clk);
  dff _90065_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _40206_, clk);
  dff _90066_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _40207_, clk);
  dff _90067_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _40209_, clk);
  dff _90068_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _40210_, clk);
  dff _90069_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39811_, clk);
  dff _90070_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _39813_, clk);
  dff _90071_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39814_, clk);
  dff _90072_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _40211_, clk);
  dff _90073_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _40212_, clk);
  dff _90074_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _40213_, clk);
  dff _90075_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39815_, clk);
  dff _90076_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _40214_, clk);
  dff _90077_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _40215_, clk);
  dff _90078_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _40216_, clk);
  dff _90079_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _40217_, clk);
  dff _90080_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _40218_, clk);
  dff _90081_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _40220_, clk);
  dff _90082_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _40221_, clk);
  dff _90083_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _40222_, clk);
  dff _90084_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _40223_, clk);
  dff _90085_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _40224_, clk);
  dff _90086_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _40225_, clk);
  dff _90087_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _40226_, clk);
  dff _90088_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _40227_, clk);
  dff _90089_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _40228_, clk);
  dff _90090_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _40229_, clk);
  dff _90091_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _40231_, clk);
  dff _90092_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _40232_, clk);
  dff _90093_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _40233_, clk);
  dff _90094_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _40234_, clk);
  dff _90095_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _40235_, clk);
  dff _90096_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _40236_, clk);
  dff _90097_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _40237_, clk);
  dff _90098_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _40238_, clk);
  dff _90099_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _40239_, clk);
  dff _90100_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _40240_, clk);
  dff _90101_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _40242_, clk);
  dff _90102_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _40243_, clk);
  dff _90103_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _40244_, clk);
  dff _90104_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _40245_, clk);
  dff _90105_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _40246_, clk);
  dff _90106_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _40247_, clk);
  dff _90107_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39817_, clk);
  dff _90108_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _40248_, clk);
  dff _90109_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _40249_, clk);
  dff _90110_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _40250_, clk);
  dff _90111_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _40251_, clk);
  dff _90112_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _40253_, clk);
  dff _90113_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _40254_, clk);
  dff _90114_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _40255_, clk);
  dff _90115_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39818_, clk);
  dff _90116_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39819_, clk);
  dff _90117_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39821_, clk);
  dff _90118_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _40256_, clk);
  dff _90119_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _40257_, clk);
  dff _90120_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _40258_, clk);
  dff _90121_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _40259_, clk);
  dff _90122_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _40260_, clk);
  dff _90123_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _40261_, clk);
  dff _90124_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _40262_, clk);
  dff _90125_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _40264_, clk);
  dff _90126_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _40265_, clk);
  dff _90127_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _40266_, clk);
  dff _90128_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _40267_, clk);
  dff _90129_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _40268_, clk);
  dff _90130_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _40269_, clk);
  dff _90131_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _40270_, clk);
  dff _90132_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _40271_, clk);
  dff _90133_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39822_, clk);
  dff _90134_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39823_, clk);
  dff _90135_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39824_, clk);
  dff _90136_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39825_, clk);
  dff _90137_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _40272_, clk);
  dff _90138_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _40273_, clk);
  dff _90139_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _40274_, clk);
  dff _90140_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _40275_, clk);
  dff _90141_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _40276_, clk);
  dff _90142_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _40277_, clk);
  dff _90143_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _40278_, clk);
  dff _90144_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _40279_, clk);
  dff _90145_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _40280_, clk);
  dff _90146_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _40281_, clk);
  dff _90147_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _40282_, clk);
  dff _90148_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _40283_, clk);
  dff _90149_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _40285_, clk);
  dff _90150_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _40286_, clk);
  dff _90151_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _40287_, clk);
  dff _90152_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39826_, clk);
  dff _90153_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39827_, clk);
  dff _90154_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40750_, clk);
  dff _90155_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40772_, clk);
  dff _90156_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40773_, clk);
  dff _90157_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40774_, clk);
  dff _90158_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40775_, clk);
  dff _90159_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40776_, clk);
  dff _90160_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40777_, clk);
  dff _90161_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40778_, clk);
  dff _90162_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40752_, clk);
  dff _90163_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40753_, clk);
  dff _90164_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40779_, clk);
  dff _90165_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40780_, clk);
  dff _90166_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40754_, clk);
  dff _90167_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03258_, clk);
  dff _90168_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03262_, clk);
  dff _90169_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03265_, clk);
  dff _90170_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03269_, clk);
  dff _90171_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03273_, clk);
  dff _90172_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03276_, clk);
  dff _90173_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03279_, clk);
  dff _90174_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02576_, clk);
  dff _90175_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03230_, clk);
  dff _90176_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03233_, clk);
  dff _90177_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03237_, clk);
  dff _90178_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03240_, clk);
  dff _90179_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03244_, clk);
  dff _90180_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03247_, clk);
  dff _90181_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03251_, clk);
  dff _90182_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03254_, clk);
  dff _90183_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03201_, clk);
  dff _90184_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03205_, clk);
  dff _90185_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03208_, clk);
  dff _90186_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03212_, clk);
  dff _90187_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03215_, clk);
  dff _90188_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03219_, clk);
  dff _90189_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03222_, clk);
  dff _90190_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03225_, clk);
  dff _90191_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02812_, clk);
  dff _90192_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02816_, clk);
  dff _90193_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02821_, clk);
  dff _90194_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02826_, clk);
  dff _90195_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02831_, clk);
  dff _90196_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02835_, clk);
  dff _90197_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02840_, clk);
  dff _90198_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02843_, clk);
  dff _90199_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02850_, clk);
  dff _90200_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02853_, clk);
  dff _90201_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02856_, clk);
  dff _90202_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02861_, clk);
  dff _90203_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02864_, clk);
  dff _90204_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02867_, clk);
  dff _90205_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02870_, clk);
  dff _90206_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02873_, clk);
  dff _90207_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02879_, clk);
  dff _90208_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02883_, clk);
  dff _90209_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02887_, clk);
  dff _90210_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02890_, clk);
  dff _90211_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02895_, clk);
  dff _90212_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02898_, clk);
  dff _90213_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02902_, clk);
  dff _90214_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02905_, clk);
  dff _90215_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02944_, clk);
  dff _90216_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02948_, clk);
  dff _90217_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02951_, clk);
  dff _90218_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02956_, clk);
  dff _90219_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02959_, clk);
  dff _90220_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02963_, clk);
  dff _90221_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02966_, clk);
  dff _90222_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02970_, clk);
  dff _90223_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02911_, clk);
  dff _90224_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02914_, clk);
  dff _90225_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02918_, clk);
  dff _90226_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02922_, clk);
  dff _90227_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02925_, clk);
  dff _90228_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02929_, clk);
  dff _90229_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02933_, clk);
  dff _90230_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02936_, clk);
  dff _90231_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03087_, clk);
  dff _90232_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03091_, clk);
  dff _90233_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03095_, clk);
  dff _90234_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03099_, clk);
  dff _90235_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03102_, clk);
  dff _90236_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03106_, clk);
  dff _90237_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03109_, clk);
  dff _90238_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03112_, clk);
  dff _90239_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03060_, clk);
  dff _90240_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03063_, clk);
  dff _90241_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03067_, clk);
  dff _90242_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03069_, clk);
  dff _90243_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03073_, clk);
  dff _90244_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03076_, clk);
  dff _90245_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03080_, clk);
  dff _90246_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03083_, clk);
  dff _90247_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03032_, clk);
  dff _90248_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03035_, clk);
  dff _90249_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03038_, clk);
  dff _90250_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03042_, clk);
  dff _90251_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03045_, clk);
  dff _90252_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03048_, clk);
  dff _90253_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03051_, clk);
  dff _90254_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03054_, clk);
  dff _90255_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _03003_, clk);
  dff _90256_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _03007_, clk);
  dff _90257_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _03010_, clk);
  dff _90258_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _03014_, clk);
  dff _90259_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _03018_, clk);
  dff _90260_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03021_, clk);
  dff _90261_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03024_, clk);
  dff _90262_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03027_, clk);
  dff _90263_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02974_, clk);
  dff _90264_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02977_, clk);
  dff _90265_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02982_, clk);
  dff _90266_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02985_, clk);
  dff _90267_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02988_, clk);
  dff _90268_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02993_, clk);
  dff _90269_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02996_, clk);
  dff _90270_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02999_, clk);
  dff _90271_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03116_, clk);
  dff _90272_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03119_, clk);
  dff _90273_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03122_, clk);
  dff _90274_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03125_, clk);
  dff _90275_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03130_, clk);
  dff _90276_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03133_, clk);
  dff _90277_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03136_, clk);
  dff _90278_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03139_, clk);
  dff _90279_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03172_, clk);
  dff _90280_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03176_, clk);
  dff _90281_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03180_, clk);
  dff _90282_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03183_, clk);
  dff _90283_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03187_, clk);
  dff _90284_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03190_, clk);
  dff _90285_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03194_, clk);
  dff _90286_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03197_, clk);
  dff _90287_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03143_, clk);
  dff _90288_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03147_, clk);
  dff _90289_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03150_, clk);
  dff _90290_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03154_, clk);
  dff _90291_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03157_, clk);
  dff _90292_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03161_, clk);
  dff _90293_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03164_, clk);
  dff _90294_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03167_, clk);
  dff _90295_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05076_, clk);
  dff _90296_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05078_, clk);
  dff _90297_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05080_, clk);
  dff _90298_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05082_, clk);
  dff _90299_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05084_, clk);
  dff _90300_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05086_, clk);
  dff _90301_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05088_, clk);
  dff _90302_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02564_, clk);
  dff _90303_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _90304_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _90305_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _90306_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _90307_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _90308_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _90309_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _90310_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _90311_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _90312_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _90313_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _90314_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _90315_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _90316_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _90317_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _90318_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _90319_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _90320_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _90321_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _90322_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _90323_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _90324_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _90325_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _90326_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _90327_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _90328_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _90329_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _90330_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _90331_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _90332_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _90333_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _90334_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _90335_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _90336_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _40590_, clk);
  dff _90337_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _40672_, clk);
  dff _90338_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _40673_, clk);
  dff _90339_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _40674_, clk);
  dff _90340_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _40592_, clk);
  dff _90341_ (\oc8051_top_1.oc8051_sfr1.bit_out , _40593_, clk);
  dff _90342_ (\oc8051_top_1.oc8051_sfr1.wait_data , _40594_, clk);
  dff _90343_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _40675_, clk);
  dff _90344_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _40677_, clk);
  dff _90345_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _40678_, clk);
  dff _90346_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _40679_, clk);
  dff _90347_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _40680_, clk);
  dff _90348_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _40681_, clk);
  dff _90349_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _40682_, clk);
  dff _90350_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _40595_, clk);
  dff _90351_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _40596_, clk);
  dff _90352_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19709_, clk);
  dff _90353_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19721_, clk);
  dff _90354_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19733_, clk);
  dff _90355_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19744_, clk);
  dff _90356_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19756_, clk);
  dff _90357_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19768_, clk);
  dff _90358_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19780_, clk);
  dff _90359_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17982_, clk);
  dff _90360_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08889_, clk);
  dff _90361_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08900_, clk);
  dff _90362_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08911_, clk);
  dff _90363_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08922_, clk);
  dff _90364_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08933_, clk);
  dff _90365_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08944_, clk);
  dff _90366_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08955_, clk);
  dff _90367_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06648_, clk);
  dff _90368_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13637_, clk);
  dff _90369_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13648_, clk);
  dff _90370_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13659_, clk);
  dff _90371_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13670_, clk);
  dff _90372_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13681_, clk);
  dff _90373_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13691_, clk);
  dff _90374_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13702_, clk);
  dff _90375_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12699_, clk);
  dff _90376_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13713_, clk);
  dff _90377_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13724_, clk);
  dff _90378_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13735_, clk);
  dff _90379_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13746_, clk);
  dff _90380_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13757_, clk);
  dff _90381_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13768_, clk);
  dff _90382_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13779_, clk);
  dff _90383_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12720_, clk);
  dff _90384_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _43638_, clk);
  dff _90385_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _43637_, clk);
  dff _90386_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _90387_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _43634_, clk);
  dff _90388_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00137_, clk);
  dff _90389_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00139_, clk);
  dff _90390_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00141_, clk);
  dff _90391_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00143_, clk);
  dff _90392_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00145_, clk);
  dff _90393_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00146_, clk);
  dff _90394_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00148_, clk);
  dff _90395_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _43632_, clk);
  dff _90396_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00150_, clk);
  dff _90397_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _43630_, clk);
  dff _90398_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _43628_, clk);
  dff _90399_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00152_, clk);
  dff _90400_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00154_, clk);
  dff _90401_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _43626_, clk);
  dff _90402_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00156_, clk);
  dff _90403_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00157_, clk);
  dff _90404_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _43624_, clk);
  dff _90405_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00159_, clk);
  dff _90406_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _43622_, clk);
  dff _90407_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00161_, clk);
  dff _90408_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _43620_, clk);
  dff _90409_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _43585_, clk);
  dff _90410_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _43584_, clk);
  dff _90411_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _43582_, clk);
  dff _90412_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _43580_, clk);
  dff _90413_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00163_, clk);
  dff _90414_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00165_, clk);
  dff _90415_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00167_, clk);
  dff _90416_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _43577_, clk);
  dff _90417_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00168_, clk);
  dff _90418_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00170_, clk);
  dff _90419_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00172_, clk);
  dff _90420_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00174_, clk);
  dff _90421_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00176_, clk);
  dff _90422_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00178_, clk);
  dff _90423_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00180_, clk);
  dff _90424_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _43575_, clk);
  dff _90425_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00181_, clk);
  dff _90426_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00183_, clk);
  dff _90427_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00185_, clk);
  dff _90428_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00187_, clk);
  dff _90429_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00189_, clk);
  dff _90430_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00191_, clk);
  dff _90431_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00192_, clk);
  dff _90432_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _43572_, clk);
  dff _90433_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41329_, clk);
  dff _90434_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41331_, clk);
  dff _90435_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41333_, clk);
  dff _90436_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41335_, clk);
  dff _90437_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41337_, clk);
  dff _90438_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41339_, clk);
  dff _90439_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41341_, clk);
  dff _90440_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _30987_, clk);
  dff _90441_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41343_, clk);
  dff _90442_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41345_, clk);
  dff _90443_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41347_, clk);
  dff _90444_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41348_, clk);
  dff _90445_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41350_, clk);
  dff _90446_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41352_, clk);
  dff _90447_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41354_, clk);
  dff _90448_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31010_, clk);
  dff _90449_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41356_, clk);
  dff _90450_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41358_, clk);
  dff _90451_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41360_, clk);
  dff _90452_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41362_, clk);
  dff _90453_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41363_, clk);
  dff _90454_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41365_, clk);
  dff _90455_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41367_, clk);
  dff _90456_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31033_, clk);
  dff _90457_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41369_, clk);
  dff _90458_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41370_, clk);
  dff _90459_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41372_, clk);
  dff _90460_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41374_, clk);
  dff _90461_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41376_, clk);
  dff _90462_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41377_, clk);
  dff _90463_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41379_, clk);
  dff _90464_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31056_, clk);
  dff _90465_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17358_, clk);
  dff _90466_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17369_, clk);
  dff _90467_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17380_, clk);
  dff _90468_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17391_, clk);
  dff _90469_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17402_, clk);
  dff _90470_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17413_, clk);
  dff _90471_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15177_, clk);
  dff _90472_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09506_, clk);
  dff _90473_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10682_, clk);
  dff _90474_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10693_, clk);
  dff _90475_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10704_, clk);
  dff _90476_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10715_, clk);
  dff _90477_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10726_, clk);
  dff _90478_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10737_, clk);
  dff _90479_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10748_, clk);
  dff _90480_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09527_, clk);
  dff _90481_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41828_, clk);
  dff _90482_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41831_, clk);
  dff _90483_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _42352_, clk);
  dff _90484_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _42354_, clk);
  dff _90485_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _42355_, clk);
  dff _90486_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _42357_, clk);
  dff _90487_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _42359_, clk);
  dff _90488_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _42361_, clk);
  dff _90489_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _42363_, clk);
  dff _90490_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41834_, clk);
  dff _90491_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _42364_, clk);
  dff _90492_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _42366_, clk);
  dff _90493_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _42368_, clk);
  dff _90494_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _42370_, clk);
  dff _90495_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _42371_, clk);
  dff _90496_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _42373_, clk);
  dff _90497_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _42375_, clk);
  dff _90498_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41837_, clk);
  dff _90499_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41840_, clk);
  dff _90500_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41843_, clk);
  dff _90501_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _42377_, clk);
  dff _90502_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _42378_, clk);
  dff _90503_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _42380_, clk);
  dff _90504_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _42382_, clk);
  dff _90505_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _42384_, clk);
  dff _90506_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _42385_, clk);
  dff _90507_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _42387_, clk);
  dff _90508_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41846_, clk);
  dff _90509_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _42389_, clk);
  dff _90510_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _42391_, clk);
  dff _90511_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _42392_, clk);
  dff _90512_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _42394_, clk);
  dff _90513_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _42396_, clk);
  dff _90514_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _42398_, clk);
  dff _90515_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _42399_, clk);
  dff _90516_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41849_, clk);
  dff _90517_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41852_, clk);
  dff _90518_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _42401_, clk);
  dff _90519_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _42402_, clk);
  dff _90520_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _42404_, clk);
  dff _90521_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _42406_, clk);
  dff _90522_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _42407_, clk);
  dff _90523_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _42409_, clk);
  dff _90524_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _42411_, clk);
  dff _90525_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41855_, clk);
  dff _90526_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01615_, clk);
  dff _90527_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01618_, clk);
  dff _90528_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01621_, clk);
  dff _90529_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01624_, clk);
  dff _90530_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02131_, clk);
  dff _90531_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02133_, clk);
  dff _90532_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02135_, clk);
  dff _90533_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02136_, clk);
  dff _90534_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02138_, clk);
  dff _90535_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02140_, clk);
  dff _90536_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02142_, clk);
  dff _90537_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01627_, clk);
  dff _90538_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02143_, clk);
  dff _90539_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02145_, clk);
  dff _90540_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02147_, clk);
  dff _90541_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02149_, clk);
  dff _90542_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02150_, clk);
  dff _90543_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02152_, clk);
  dff _90544_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02154_, clk);
  dff _90545_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01630_, clk);
  dff _90546_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01633_, clk);
  dff _90547_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02156_, clk);
  dff _90548_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02157_, clk);
  dff _90549_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02159_, clk);
  dff _90550_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02161_, clk);
  dff _90551_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02163_, clk);
  dff _90552_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02164_, clk);
  dff _90553_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02166_, clk);
  dff _90554_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01636_, clk);
  dff _90555_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02168_, clk);
  dff _90556_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02170_, clk);
  dff _90557_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02171_, clk);
  dff _90558_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02173_, clk);
  dff _90559_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02175_, clk);
  dff _90560_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02177_, clk);
  dff _90561_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02178_, clk);
  dff _90562_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01639_, clk);
  dff _90563_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01642_, clk);
  dff _90564_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02180_, clk);
  dff _90565_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02182_, clk);
  dff _90566_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02184_, clk);
  dff _90567_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02185_, clk);
  dff _90568_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02186_, clk);
  dff _90569_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02187_, clk);
  dff _90570_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02188_, clk);
  dff _90571_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01645_, clk);
  dff _90572_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01218_, clk);
  dff _90573_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01220_, clk);
  dff _90574_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01222_, clk);
  dff _90575_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01224_, clk);
  dff _90576_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01226_, clk);
  dff _90577_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01228_, clk);
  dff _90578_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01230_, clk);
  dff _90579_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01232_, clk);
  dff _90580_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01234_, clk);
  dff _90581_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01236_, clk);
  dff _90582_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01238_, clk);
  dff _90583_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00574_, clk);
  dff _90584_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00550_, clk);
  dff _90585_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00552_, clk);
  dff _90586_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00555_, clk);
  dff _90587_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00558_, clk);
  dff _90588_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00561_, clk);
  dff _90589_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00563_, clk);
  dff _90590_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01240_, clk);
  dff _90591_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00566_, clk);
  dff _90592_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01242_, clk);
  dff _90593_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01244_, clk);
  dff _90594_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01245_, clk);
  dff _90595_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00569_, clk);
  dff _90596_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01247_, clk);
  dff _90597_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01249_, clk);
  dff _90598_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01251_, clk);
  dff _90599_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01253_, clk);
  dff _90600_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01255_, clk);
  dff _90601_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01257_, clk);
  dff _90602_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01259_, clk);
  dff _90603_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00571_, clk);
  dff _90604_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00577_, clk);
  dff _90605_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00579_, clk);
  dff _90606_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00582_, clk);
  dff _90607_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00585_, clk);
  dff _90608_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00587_, clk);
  dff _90609_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01261_, clk);
  dff _90610_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01263_, clk);
  dff _90611_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01265_, clk);
  dff _90612_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00590_, clk);
  dff _90613_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01267_, clk);
  dff _90614_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01269_, clk);
  dff _90615_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01271_, clk);
  dff _90616_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01273_, clk);
  dff _90617_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01275_, clk);
  dff _90618_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01276_, clk);
  dff _90619_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01278_, clk);
  dff _90620_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01280_, clk);
  dff _90621_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01282_, clk);
  dff _90622_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01284_, clk);
  dff _90623_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00593_, clk);
  dff _90624_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01286_, clk);
  dff _90625_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01288_, clk);
  dff _90626_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01290_, clk);
  dff _90627_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01292_, clk);
  dff _90628_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01294_, clk);
  dff _90629_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01296_, clk);
  dff _90630_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01298_, clk);
  dff _90631_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00595_, clk);
  dff _90632_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01299_, clk);
  dff _90633_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01300_, clk);
  dff _90634_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01301_, clk);
  dff _90635_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01303_, clk);
  dff _90636_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01305_, clk);
  dff _90637_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01307_, clk);
  dff _90638_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01309_, clk);
  dff _90639_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00598_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1090 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1090 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1090 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1090 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1092 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1092 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1094 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1094 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1094 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1095 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1095 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1095 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1096 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1096 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1096 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1097 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1097 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1097 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1098 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1098 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1098 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1099 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1099 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1100 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1175 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1176 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1176 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1176 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1176 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1176 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1176 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1176 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1176 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1177 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1177 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1177 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1177 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1177 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1177 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1177 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1177 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1178 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1178 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1178 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1178 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1178 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1178 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1178 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1178 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1179 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1180 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1182 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1184 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1184 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1184 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1184 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1184 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1184 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1184 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1211 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1211 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1211 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1211 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1211 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1211 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1211 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1211 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1211 [9], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1211 [10], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1211 [11], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1211 [12], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1211 [13], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1211 [14], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1211 [15], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1213 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1213 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1213 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1213 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1213 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1213 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1213 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1213 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1215 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1215 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1215 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1215 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1215 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1215 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1215 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1215 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1219 [8], \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1220 , \oc8051_golden_model_1.n1237 [7]);
  buf(\oc8051_golden_model_1.n1221 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1221 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1221 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1221 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1222 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1222 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1222 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1222 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1226 [4], \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1227 , \oc8051_golden_model_1.n1237 [6]);
  buf(\oc8051_golden_model_1.n1228 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1228 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1228 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1228 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1228 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1228 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1228 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1228 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1228 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1236 , \oc8051_golden_model_1.n1237 [2]);
  buf(\oc8051_golden_model_1.n1237 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1237 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1237 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1237 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1237 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1242 , \oc8051_golden_model_1.n1257 [7]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.n1257 [6]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.n1257 [2]);
  buf(\oc8051_golden_model_1.n1257 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1257 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1257 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1257 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1257 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1259 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1259 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1259 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1259 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1259 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1259 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1259 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1259 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1259 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1262 , \oc8051_golden_model_1.n1276 [7]);
  buf(\oc8051_golden_model_1.n1263 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1263 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1263 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1263 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.n1913 [0]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.n1913 [1]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.n1913 [2]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.n1913 [3]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1268 [8], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1276 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1288 [6]);
  buf(\oc8051_golden_model_1.n1279 [8], \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1288 [7]);
  buf(\oc8051_golden_model_1.n1287 , \oc8051_golden_model_1.n1288 [2]);
  buf(\oc8051_golden_model_1.n1288 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1288 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1288 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1288 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1288 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1290 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1290 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1290 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1290 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1290 [4], \oc8051_golden_model_1.n1298 [4]);
  buf(\oc8051_golden_model_1.n1290 [5], \oc8051_golden_model_1.n1298 [5]);
  buf(\oc8051_golden_model_1.n1290 [6], \oc8051_golden_model_1.n1298 [6]);
  buf(\oc8051_golden_model_1.n1290 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1290 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1292 [8], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1293 , \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1294 [0], \oc8051_golden_model_1.n1298 [0]);
  buf(\oc8051_golden_model_1.n1294 [1], \oc8051_golden_model_1.n1298 [1]);
  buf(\oc8051_golden_model_1.n1294 [2], \oc8051_golden_model_1.n1298 [2]);
  buf(\oc8051_golden_model_1.n1294 [3], \oc8051_golden_model_1.n1298 [3]);
  buf(\oc8051_golden_model_1.n1294 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1297 , \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1298 [7], \oc8051_golden_model_1.n1298 [8]);
  buf(\oc8051_golden_model_1.n1305 , \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1306 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1306 [2], \oc8051_golden_model_1.n1310 [2]);
  buf(\oc8051_golden_model_1.n1306 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1306 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1306 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1306 [6], \oc8051_golden_model_1.n1322 [6]);
  buf(\oc8051_golden_model_1.n1306 [7], \oc8051_golden_model_1.n1310 [7]);
  buf(\oc8051_golden_model_1.n1308 [4], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1309 , \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1310 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1310 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1310 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1310 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1310 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1310 [6], \oc8051_golden_model_1.n1321 [6]);
  buf(\oc8051_golden_model_1.n1312 [8], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1313 , \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1321 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1321 [2], \oc8051_golden_model_1.n1322 [2]);
  buf(\oc8051_golden_model_1.n1321 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1321 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1321 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1321 [7], \oc8051_golden_model_1.n1322 [7]);
  buf(\oc8051_golden_model_1.n1322 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1322 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1322 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1322 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1322 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1326 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1326 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1326 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1326 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1326 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1326 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1326 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1327 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1327 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1327 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1327 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1327 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1327 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1327 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1327 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1329 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1329 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1329 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1329 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1329 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1329 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1329 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1329 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1330 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1330 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1330 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1333 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1333 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1335 [8], \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1336 , \oc8051_golden_model_1.n1348 [7]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1337 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1337 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1339 [4], \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1348 [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.n1348 [2]);
  buf(\oc8051_golden_model_1.n1348 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1348 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1348 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1348 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1348 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1352 [8], \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.n1364 [7]);
  buf(\oc8051_golden_model_1.n1355 [4], \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1356 , \oc8051_golden_model_1.n1364 [6]);
  buf(\oc8051_golden_model_1.n1363 , \oc8051_golden_model_1.n1364 [2]);
  buf(\oc8051_golden_model_1.n1364 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1364 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1364 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1364 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1364 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1368 [8], \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1369 , \oc8051_golden_model_1.n1380 [7]);
  buf(\oc8051_golden_model_1.n1371 [4], \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1372 , \oc8051_golden_model_1.n1380 [6]);
  buf(\oc8051_golden_model_1.n1379 , \oc8051_golden_model_1.n1380 [2]);
  buf(\oc8051_golden_model_1.n1380 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1380 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1380 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1380 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1380 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1384 [8], \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1385 , \oc8051_golden_model_1.n1396 [7]);
  buf(\oc8051_golden_model_1.n1387 [4], \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1388 , \oc8051_golden_model_1.n1396 [6]);
  buf(\oc8051_golden_model_1.n1395 , \oc8051_golden_model_1.n1396 [2]);
  buf(\oc8051_golden_model_1.n1396 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1396 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1396 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1396 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1396 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.n1558 [7]);
  buf(\oc8051_golden_model_1.n1557 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1557 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1557 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1557 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1557 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1557 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1557 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1558 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1558 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1558 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1558 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1558 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1558 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1558 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1581 , \oc8051_golden_model_1.n1582 [7]);
  buf(\oc8051_golden_model_1.n1582 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1589 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1589 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1589 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1589 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1590 , \oc8051_golden_model_1.n1591 [2]);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1591 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1591 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1591 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1591 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1591 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1735 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1738 , \oc8051_golden_model_1.n1747 [7]);
  buf(\oc8051_golden_model_1.n1740 , \oc8051_golden_model_1.n1747 [6]);
  buf(\oc8051_golden_model_1.n1746 , \oc8051_golden_model_1.n1747 [2]);
  buf(\oc8051_golden_model_1.n1747 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1751 , \oc8051_golden_model_1.n1760 [7]);
  buf(\oc8051_golden_model_1.n1753 , \oc8051_golden_model_1.n1760 [6]);
  buf(\oc8051_golden_model_1.n1759 , \oc8051_golden_model_1.n1760 [2]);
  buf(\oc8051_golden_model_1.n1760 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1760 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1760 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1760 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1760 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1764 , \oc8051_golden_model_1.n1773 [7]);
  buf(\oc8051_golden_model_1.n1766 , \oc8051_golden_model_1.n1773 [6]);
  buf(\oc8051_golden_model_1.n1772 , \oc8051_golden_model_1.n1773 [2]);
  buf(\oc8051_golden_model_1.n1773 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1773 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1773 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1773 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1773 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1786 [7]);
  buf(\oc8051_golden_model_1.n1779 , \oc8051_golden_model_1.n1786 [6]);
  buf(\oc8051_golden_model_1.n1785 , \oc8051_golden_model_1.n1786 [2]);
  buf(\oc8051_golden_model_1.n1786 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1786 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1786 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1786 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1786 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1788 , \oc8051_golden_model_1.n1789 [7]);
  buf(\oc8051_golden_model_1.n1789 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1789 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1789 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1789 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1789 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1789 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1789 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1794 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1794 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1794 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1794 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1794 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1794 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1794 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1794 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1794 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1794 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1800 , \oc8051_golden_model_1.n1801 [2]);
  buf(\oc8051_golden_model_1.n1801 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1801 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1801 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1801 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1801 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1801 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1801 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [7]);
  buf(\oc8051_golden_model_1.n1805 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1825 , \oc8051_golden_model_1.n1826 [7]);
  buf(\oc8051_golden_model_1.n1826 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1826 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1826 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1826 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1826 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1826 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1826 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1831 , \oc8051_golden_model_1.n1832 [7]);
  buf(\oc8051_golden_model_1.n1832 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1832 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1832 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1832 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1832 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1832 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1832 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1837 , \oc8051_golden_model_1.n1838 [7]);
  buf(\oc8051_golden_model_1.n1838 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1838 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1838 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1838 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1838 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1838 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1838 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1843 , \oc8051_golden_model_1.n1844 [7]);
  buf(\oc8051_golden_model_1.n1844 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1844 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1844 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1844 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1844 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1844 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1844 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1849 , \oc8051_golden_model_1.n1850 [7]);
  buf(\oc8051_golden_model_1.n1850 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1850 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1850 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1850 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1850 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1850 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1850 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1851 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1851 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1851 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1851 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1851 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1851 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1851 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1852 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1853 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1853 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1853 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1889 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1889 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1889 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1889 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1889 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1889 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1889 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1889 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1908 , \oc8051_golden_model_1.n1909 [7]);
  buf(\oc8051_golden_model_1.n1909 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1909 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1909 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1909 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1909 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1909 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1909 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1913 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1913 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1913 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1913 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1914 [0], \oc8051_golden_model_1.n1915 [4]);
  buf(\oc8051_golden_model_1.n1914 [1], \oc8051_golden_model_1.n1915 [5]);
  buf(\oc8051_golden_model_1.n1914 [2], \oc8051_golden_model_1.n1915 [6]);
  buf(\oc8051_golden_model_1.n1914 [3], \oc8051_golden_model_1.n1915 [7]);
  buf(\oc8051_golden_model_1.n1915 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1915 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1915 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1915 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
