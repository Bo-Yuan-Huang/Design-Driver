
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jnc, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jnc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _14054_ (_05685_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not _14055_ (_05686_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _14056_ (_05687_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor _14057_ (_05688_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _14058_ (_05689_, _05688_, _05687_);
  and _14059_ (_05690_, _05689_, _05686_);
  and _14060_ (_05691_, _05690_, _05685_);
  nor _14061_ (_05692_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14062_ (_05693_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not _14063_ (_05694_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _14064_ (_05695_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14065_ (_05696_, _05695_, _05694_);
  or _14066_ (_05697_, _05696_, _05693_);
  not _14067_ (_05698_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _14068_ (_05699_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05698_);
  nand _14069_ (_05700_, _05699_, _05694_);
  not _14070_ (_05701_, _05700_);
  nand _14071_ (_05702_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _14072_ (_05703_, _05702_, _05697_);
  nand _14073_ (_05704_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14074_ (_05705_, _05704_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _14075_ (_05706_, _05705_);
  nand _14076_ (_05707_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not _14077_ (_05708_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  not _14078_ (_05709_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _14079_ (_05710_, _05694_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nand _14080_ (_05711_, _05710_, _05709_);
  or _14081_ (_05712_, _05711_, _05708_);
  and _14082_ (_05713_, _05712_, _05707_);
  and _14083_ (_05714_, _05695_, _05694_);
  nand _14084_ (_05715_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _14085_ (_05716_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _14086_ (_05717_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or _14087_ (_05718_, _05717_, _05694_);
  or _14088_ (_05719_, _05718_, _05716_);
  and _14089_ (_05720_, _05719_, _05715_);
  and _14090_ (_05721_, _05720_, _05713_);
  nand _14091_ (_05722_, _05721_, _05703_);
  nand _14092_ (_05723_, _05722_, _05692_);
  and _14093_ (_05724_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14094_ (_05725_, _05724_);
  nand _14095_ (_05726_, _05725_, _05723_);
  not _14096_ (_05727_, _05726_);
  or _14097_ (_05728_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand _14098_ (_05729_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _14099_ (_05730_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _14100_ (_05731_, _05730_, _05729_);
  not _14101_ (_05732_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _14102_ (_05733_, _05711_, _05732_);
  not _14103_ (_05734_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _14104_ (_05735_, _05700_, _05734_);
  and _14105_ (_05736_, _05735_, _05733_);
  not _14106_ (_05737_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _14107_ (_05738_, _05696_, _05737_);
  not _14108_ (_05739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or _14109_ (_05740_, _05718_, _05739_);
  and _14110_ (_05741_, _05740_, _05738_);
  and _14111_ (_05742_, _05741_, _05736_);
  and _14112_ (_05743_, _05742_, _05731_);
  or _14113_ (_05744_, _05743_, _05728_);
  and _14114_ (_05745_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14115_ (_05746_, _05745_);
  nand _14116_ (_05747_, _05746_, _05744_);
  not _14117_ (_05748_, _05747_);
  not _14118_ (_05749_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _14119_ (_05751_, _05696_, _05749_);
  nand _14120_ (_05752_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _14121_ (_05753_, _05752_, _05751_);
  not _14122_ (_05754_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _14123_ (_05755_, _05705_, _05754_);
  not _14124_ (_05756_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _14125_ (_05757_, _05711_, _05756_);
  and _14126_ (_05758_, _05757_, _05755_);
  nand _14127_ (_05759_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not _14128_ (_05760_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or _14129_ (_05761_, _05718_, _05760_);
  and _14130_ (_05762_, _05761_, _05759_);
  and _14131_ (_05763_, _05762_, _05758_);
  and _14132_ (_05764_, _05763_, _05753_);
  or _14133_ (_05765_, _05764_, _05728_);
  and _14134_ (_05766_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14135_ (_05767_, _05766_);
  nand _14136_ (_05768_, _05767_, _05765_);
  and _14137_ (_05769_, _05768_, _05748_);
  and _14138_ (_05770_, _05769_, _05727_);
  and _14139_ (_05771_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14140_ (_05772_, _05771_);
  not _14141_ (_05773_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or _14142_ (_05774_, _05718_, _05773_);
  nand _14143_ (_05775_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _14144_ (_05776_, _05775_, _05774_);
  nand _14145_ (_05777_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _14146_ (_05778_, _05711_);
  nand _14147_ (_05779_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _14148_ (_05780_, _05779_, _05777_);
  and _14149_ (_05781_, _05780_, _05776_);
  not _14150_ (_05782_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _14151_ (_05783_, _05696_, _05782_);
  nand _14152_ (_05784_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _14153_ (_05785_, _05784_, _05783_);
  and _14154_ (_05786_, _05785_, _05781_);
  or _14155_ (_05787_, _05786_, _05728_);
  nand _14156_ (_05788_, _05787_, _05772_);
  not _14157_ (_05789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _14158_ (_05790_, _05718_, _05789_);
  not _14159_ (_05791_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _14160_ (_05792_, _05705_, _05791_);
  not _14161_ (_05793_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _14162_ (_05794_, _05711_, _05793_);
  and _14163_ (_05795_, _05794_, _05792_);
  and _14164_ (_05796_, _05795_, _05790_);
  nand _14165_ (_05797_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  not _14166_ (_05798_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _14167_ (_05799_, _05700_, _05798_);
  and _14168_ (_05800_, _05799_, _05797_);
  not _14169_ (_05801_, _05696_);
  and _14170_ (_05802_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _14171_ (_05803_, _05802_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _14172_ (_05804_, _05803_, _05800_);
  nand _14173_ (_05805_, _05804_, _05796_);
  or _14174_ (_05806_, _05805_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14175_ (_05807_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14176_ (_05808_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not _14177_ (_05809_, _05808_);
  and _14178_ (_05810_, _05809_, _05806_);
  not _14179_ (_05811_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _14180_ (_05812_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nand _14181_ (_05813_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _14182_ (_05814_, _05813_, _05812_);
  not _14183_ (_05815_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _14184_ (_05816_, _05696_, _05815_);
  not _14185_ (_05817_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or _14186_ (_05818_, _05718_, _05817_);
  and _14187_ (_05819_, _05818_, _05816_);
  nand _14188_ (_05820_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand _14189_ (_05821_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _14190_ (_05822_, _05821_, _05820_);
  and _14191_ (_05823_, _05822_, _05819_);
  nand _14192_ (_05824_, _05823_, _05814_);
  nand _14193_ (_05825_, _05824_, _05811_);
  nand _14194_ (_05826_, _05825_, _05807_);
  nor _14195_ (_05827_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _05807_);
  not _14196_ (_05828_, _05827_);
  and _14197_ (_05829_, _05828_, _05826_);
  nand _14198_ (_05830_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand _14199_ (_05831_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _14200_ (_05832_, _05831_, _05830_);
  not _14201_ (_05833_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _14202_ (_05834_, _05696_, _05833_);
  not _14203_ (_05835_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _14204_ (_05836_, _05718_, _05835_);
  and _14205_ (_05837_, _05836_, _05834_);
  nand _14206_ (_05838_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _14207_ (_05839_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and _14208_ (_05840_, _05839_, _05838_);
  and _14209_ (_05841_, _05840_, _05837_);
  nand _14210_ (_05842_, _05841_, _05832_);
  nand _14211_ (_05843_, _05842_, _05811_);
  nand _14212_ (_05844_, _05843_, _05807_);
  nor _14213_ (_05845_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not _14214_ (_05846_, _05845_);
  and _14215_ (_05847_, _05846_, _05844_);
  nor _14216_ (_05848_, _05847_, _05829_);
  and _14217_ (_05849_, _05848_, _05810_);
  and _14218_ (_05850_, _05849_, _05788_);
  and _14219_ (_05851_, _05850_, _05770_);
  not _14220_ (_05852_, _05788_);
  and _14221_ (_05853_, _05849_, _05852_);
  nor _14222_ (_05854_, _05768_, _05747_);
  and _14223_ (_05855_, _05854_, _05726_);
  and _14224_ (_05856_, _05855_, _05853_);
  not _14225_ (_05857_, _05847_);
  not _14226_ (_05858_, _05810_);
  and _14227_ (_05859_, _05829_, _05858_);
  and _14228_ (_05860_, _05859_, _05857_);
  and _14229_ (_05861_, _05860_, _05852_);
  not _14230_ (_05862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _14231_ (_05863_, _05696_, _05862_);
  and _14232_ (_05864_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not _14233_ (_05865_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _14234_ (_05866_, _05718_, _05865_);
  and _14235_ (_05867_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _14236_ (_05868_, _05867_, _05866_);
  nand _14237_ (_05869_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nand _14238_ (_05870_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _14239_ (_05871_, _05870_, _05869_);
  nand _14240_ (_05872_, _05871_, _05868_);
  or _14241_ (_05873_, _05872_, _05864_);
  or _14242_ (_05874_, _05873_, _05863_);
  or _14243_ (_05875_, _05874_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _14244_ (_05876_, _05875_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14245_ (_05878_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not _14246_ (_05879_, _05878_);
  and _14247_ (_05880_, _05879_, _05876_);
  not _14248_ (_05881_, _05880_);
  and _14249_ (_05882_, _05881_, _05769_);
  and _14250_ (_05883_, _05882_, _05861_);
  or _14251_ (_05884_, _05883_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _14252_ (_05885_, _05884_, _05856_);
  or _14253_ (_05886_, _05885_, _05851_);
  and _14254_ (_05887_, _05886_, _05691_);
  nor _14255_ (_05888_, _05690_, _05685_);
  or _14256_ (_05889_, _05888_, rst);
  or _14257_ (_00393_, _05889_, _05887_);
  and _14258_ (_05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _14259_ (_05891_, _05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _14260_ (_05892_, _05891_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _14261_ (_05893_, _05892_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _14262_ (_05894_, _05893_);
  not _14263_ (_05895_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14264_ (_05896_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05686_);
  and _14265_ (_05897_, _05896_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _14266_ (_05898_, _05897_, _05895_);
  not _14267_ (_05899_, _05898_);
  nor _14268_ (_05900_, _05892_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _14269_ (_05901_, _05900_, _05899_);
  and _14270_ (_05902_, _05901_, _05894_);
  not _14271_ (_05903_, _05902_);
  nor _14272_ (_05904_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor _14273_ (_05905_, _05904_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _14274_ (_05906_, _05905_, _05896_);
  and _14275_ (_05907_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  not _14276_ (_05908_, _05907_);
  and _14277_ (_05909_, _05897_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14278_ (_05910_, _05904_, _05896_);
  and _14279_ (_05911_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _14280_ (_05912_, _05911_, _05909_);
  and _14281_ (_05913_, _05912_, _05908_);
  not _14282_ (_05914_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _14283_ (_05915_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05686_);
  and _14284_ (_05916_, _05915_, _05914_);
  and _14285_ (_05917_, _05916_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14286_ (_05918_, _05917_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _14287_ (_05919_, _05916_, _05895_);
  and _14288_ (_05920_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  nor _14289_ (_05921_, _05920_, _05918_);
  and _14290_ (_05922_, _05921_, _05913_);
  and _14291_ (_05923_, _05922_, _05903_);
  and _14292_ (_05924_, _05893_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _14293_ (_05925_, _05924_);
  nor _14294_ (_05926_, _05893_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _14295_ (_05927_, _05926_, _05899_);
  and _14296_ (_05928_, _05927_, _05925_);
  not _14297_ (_05929_, _05928_);
  and _14298_ (_05930_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _14299_ (_05931_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _14300_ (_05932_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or _14301_ (_05933_, _05932_, _05931_);
  or _14302_ (_05934_, _05933_, _05909_);
  nor _14303_ (_05936_, _05934_, _05930_);
  and _14304_ (_05937_, _05936_, _05929_);
  and _14305_ (_05938_, _05937_, _05923_);
  and _14306_ (_05939_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _14307_ (_05940_, _05939_);
  nor _14308_ (_05941_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _14309_ (_05943_, _05941_, _05899_);
  and _14310_ (_05944_, _05943_, _05940_);
  not _14311_ (_05945_, _05944_);
  and _14312_ (_05946_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  not _14313_ (_05947_, _05946_);
  and _14314_ (_05948_, _05919_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not _14315_ (_05949_, _05948_);
  and _14316_ (_05950_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nor _14317_ (_05951_, _05950_, _05909_);
  and _14318_ (_05952_, _05951_, _05949_);
  and _14319_ (_05953_, _05952_, _05947_);
  and _14320_ (_05954_, _05953_, _05945_);
  not _14321_ (_05955_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _14322_ (_05956_, _05939_, _05955_);
  and _14323_ (_05957_, _05939_, _05955_);
  nor _14324_ (_05958_, _05957_, _05956_);
  nor _14325_ (_05959_, _05958_, _05899_);
  not _14326_ (_05960_, _05959_);
  and _14327_ (_05961_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _14328_ (_05962_, _05917_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and _14329_ (_05963_, _05919_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or _14330_ (_05964_, _05963_, _05962_);
  or _14331_ (_05965_, _05964_, _05909_);
  nor _14332_ (_05966_, _05965_, _05961_);
  and _14333_ (_05967_, _05966_, _05960_);
  nor _14334_ (_05968_, _05967_, _05954_);
  and _14335_ (_05969_, _05968_, _05938_);
  nor _14336_ (_05970_, _05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _14337_ (_05971_, _05970_, _05891_);
  and _14338_ (_05972_, _05971_, _05898_);
  and _14339_ (_05973_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _14340_ (_05975_, _05973_, _05972_);
  and _14341_ (_05976_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _14342_ (_05977_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _14343_ (_05978_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _14344_ (_05979_, _05978_, _05977_);
  nor _14345_ (_05980_, _05979_, _05976_);
  and _14346_ (_05981_, _05980_, _05975_);
  not _14347_ (_05982_, _05981_);
  nor _14348_ (_05983_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _14349_ (_05984_, _05983_, _05890_);
  and _14350_ (_05985_, _05984_, _05898_);
  and _14351_ (_05986_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _14352_ (_05987_, _05986_, _05985_);
  and _14353_ (_05988_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _14354_ (_05989_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _14355_ (_05990_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _14356_ (_05991_, _05990_, _05989_);
  nor _14357_ (_05992_, _05991_, _05988_);
  and _14358_ (_05993_, _05992_, _05987_);
  and _14359_ (_05994_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _14360_ (_05995_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _14361_ (_05996_, _05995_, _05994_);
  not _14362_ (_05997_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14363_ (_05998_, _05898_, _05997_);
  not _14364_ (_05999_, _05998_);
  and _14365_ (_06000_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _14366_ (_06001_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _14367_ (_06002_, _06001_, _06000_);
  and _14368_ (_06003_, _06002_, _05999_);
  and _14369_ (_06004_, _06003_, _05996_);
  and _14370_ (_06005_, _06004_, _05993_);
  and _14371_ (_06006_, _06005_, _05982_);
  and _14372_ (_06007_, _05896_, _05895_);
  not _14373_ (_06008_, _06007_);
  not _14374_ (_06009_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _14375_ (_06010_, \oc8051_top_1.oc8051_decoder1.wr , _05686_);
  and _14376_ (_06011_, _06010_, _06009_);
  and _14377_ (_06012_, _06011_, _06008_);
  not _14378_ (_06013_, _06012_);
  not _14379_ (_06014_, _05892_);
  nor _14380_ (_06015_, _05891_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _14381_ (_06016_, _06015_, _05899_);
  and _14382_ (_06017_, _06016_, _06014_);
  not _14383_ (_06018_, _06017_);
  and _14384_ (_06019_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _14385_ (_06020_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _14386_ (_06021_, _06020_, _06019_);
  and _14387_ (_06022_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _14388_ (_06023_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _14389_ (_06024_, _06023_, _06022_);
  and _14390_ (_06025_, _06024_, _06021_);
  and _14391_ (_06026_, _06025_, _06018_);
  nor _14392_ (_06027_, _06026_, _06013_);
  and _14393_ (_06028_, _06027_, _06006_);
  and _14394_ (_06029_, _06028_, _05969_);
  not _14395_ (_06030_, _06004_);
  and _14396_ (_06031_, _06030_, _05993_);
  and _14397_ (_06032_, _06031_, _05982_);
  and _14398_ (_06033_, _06027_, _05969_);
  and _14399_ (_06035_, _06033_, _06032_);
  nor _14400_ (_06036_, _06035_, _06029_);
  and _14401_ (_06037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _14402_ (_06038_, _06037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _14403_ (_06039_, _06038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _14404_ (_06040_, _06039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _14405_ (_06041_, _06040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _14406_ (_06042_, _06041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _14407_ (_06043_, _06042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _14408_ (_06044_, _06043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _14409_ (_06045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _14410_ (_06046_, _06045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _14411_ (_06047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _14412_ (_06048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _14413_ (_06050_, _06048_, _06047_);
  and _14414_ (_06051_, _06050_, _06046_);
  and _14415_ (_06053_, _06051_, _06044_);
  nor _14416_ (_06054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _14417_ (_06055_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _14418_ (_06056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _14419_ (_06057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _06056_);
  and _14420_ (_06058_, _06057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _14421_ (_06059_, _06058_, _06055_);
  not _14422_ (_06061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _14423_ (_06062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _14424_ (_06064_, _06062_, _06054_);
  and _14425_ (_06065_, _06064_, _06061_);
  not _14426_ (_06066_, _06065_);
  and _14427_ (_06067_, _06066_, _06059_);
  and _14428_ (_06068_, _06067_, _06054_);
  nand _14429_ (_06069_, _06068_, _06053_);
  nand _14430_ (_06070_, _06069_, _06036_);
  not _14431_ (_06071_, rst);
  or _14432_ (_06072_, _06036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _14433_ (_06073_, _06072_, _06071_);
  and _14434_ (_05877_, _06073_, _06070_);
  not _14435_ (_06075_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  not _14436_ (_06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _14437_ (_06077_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06076_);
  or _14438_ (_06078_, _06077_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _14439_ (_06079_, _06078_, _06075_);
  not _14440_ (_06080_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  not _14441_ (_06081_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _14442_ (_06082_, _06081_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _14443_ (_06083_, _06082_, _06076_);
  or _14444_ (_06084_, _06083_, _06080_);
  and _14445_ (_06085_, _06084_, _06079_);
  not _14446_ (_06086_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _14447_ (_06087_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _14448_ (_06088_, _06087_, _06081_);
  or _14449_ (_06089_, _06088_, _06086_);
  not _14450_ (_06090_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or _14451_ (_06091_, _06077_, _06081_);
  or _14452_ (_06093_, _06091_, _06090_);
  and _14453_ (_06094_, _06093_, _06089_);
  and _14454_ (_06095_, _06094_, _06085_);
  or _14455_ (_06097_, _06087_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _14456_ (_06098_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _14457_ (_06099_, _06098_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14458_ (_06100_, _06099_, ABINPUT[8]);
  nand _14459_ (_06101_, _06098_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14460_ (_06102_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _14461_ (_06103_, _06102_, _06100_);
  or _14462_ (_06104_, _06103_, _06097_);
  not _14463_ (_06105_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _14464_ (_06106_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _14465_ (_06107_, _06106_, _06081_);
  or _14466_ (_06108_, _06107_, _06105_);
  and _14467_ (_06109_, _06106_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14468_ (_06110_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and _14469_ (_06111_, _06110_, _06108_);
  and _14470_ (_06112_, _06111_, _06104_);
  and _14471_ (_06113_, _06112_, _06095_);
  and _14472_ (_06114_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _14473_ (_06115_, _06114_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor _14474_ (_06116_, _06099_, ABINPUT[0]);
  nor _14475_ (_06117_, _06101_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _14476_ (_06118_, _06117_, _06116_);
  nor _14477_ (_06119_, _06118_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _14478_ (_06120_, _06119_, _06115_);
  and _14479_ (_06121_, _06120_, _06113_);
  not _14480_ (_06122_, _06121_);
  and _14481_ (_06123_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05686_);
  and _14482_ (_06124_, _06123_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14483_ (_06125_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05686_);
  and _14484_ (_06126_, _06125_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14485_ (_06127_, _06126_, _06124_);
  not _14486_ (_06128_, _06127_);
  or _14487_ (_06129_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14488_ (_06131_, _06129_, _06103_);
  nand _14489_ (_06132_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14490_ (_06133_, _06132_, _06075_);
  not _14491_ (_06134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _14492_ (_06135_, _06134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14493_ (_06136_, _06135_, _06105_);
  and _14494_ (_06137_, _06136_, _06133_);
  and _14495_ (_06138_, _06137_, _06131_);
  not _14496_ (_06139_, _06138_);
  nor _14497_ (_06140_, _06139_, _06120_);
  nor _14498_ (_06141_, _06140_, _06128_);
  and _14499_ (_06142_, _06141_, _06122_);
  not _14500_ (_06143_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _14501_ (_06144_, _06123_, _06143_);
  and _14502_ (_06145_, _06144_, _06126_);
  not _14503_ (_06146_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  or _14504_ (_06147_, _06078_, _06146_);
  not _14505_ (_06148_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or _14506_ (_06149_, _06083_, _06148_);
  and _14507_ (_06150_, _06149_, _06147_);
  not _14508_ (_06151_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _14509_ (_06152_, _06088_, _06151_);
  not _14510_ (_06153_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or _14511_ (_06154_, _06091_, _06153_);
  and _14512_ (_06155_, _06154_, _06152_);
  and _14513_ (_06156_, _06155_, _06150_);
  or _14514_ (_06157_, _06099_, ABINPUT[5]);
  or _14515_ (_06158_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _14516_ (_06159_, _06158_, _06157_);
  or _14517_ (_06160_, _06159_, _06097_);
  not _14518_ (_06161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _14519_ (_06162_, _06107_, _06161_);
  nand _14520_ (_06163_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _14521_ (_06164_, _06163_, _06162_);
  and _14522_ (_06165_, _06164_, _06160_);
  and _14523_ (_06166_, _06165_, _06156_);
  not _14524_ (_06167_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  or _14525_ (_06168_, _06083_, _06167_);
  not _14526_ (_06169_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  or _14527_ (_06170_, _06078_, _06169_);
  and _14528_ (_06171_, _06170_, _06168_);
  not _14529_ (_06172_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _14530_ (_06173_, _06088_, _06172_);
  not _14531_ (_06174_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or _14532_ (_06175_, _06091_, _06174_);
  and _14533_ (_06176_, _06175_, _06173_);
  and _14534_ (_06177_, _06176_, _06171_);
  or _14535_ (_06178_, _06099_, ABINPUT[4]);
  or _14536_ (_06179_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _14537_ (_06180_, _06179_, _06178_);
  or _14538_ (_06181_, _06180_, _06097_);
  nand _14539_ (_06182_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _14540_ (_06183_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _14541_ (_06184_, _06107_, _06183_);
  and _14542_ (_06185_, _06184_, _06182_);
  and _14543_ (_06186_, _06185_, _06181_);
  and _14544_ (_06187_, _06186_, _06177_);
  not _14545_ (_06188_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  or _14546_ (_06189_, _06078_, _06188_);
  not _14547_ (_06190_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  or _14548_ (_06191_, _06083_, _06190_);
  and _14549_ (_06192_, _06191_, _06189_);
  not _14550_ (_06193_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _14551_ (_06194_, _06088_, _06193_);
  not _14552_ (_06195_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _14553_ (_06196_, _06091_, _06195_);
  nor _14554_ (_06197_, _06196_, _06194_);
  and _14555_ (_06198_, _06197_, _06192_);
  or _14556_ (_06200_, _06099_, ABINPUT[1]);
  or _14557_ (_06201_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _14558_ (_06202_, _06201_, _06200_);
  or _14559_ (_06203_, _06202_, _06097_);
  not _14560_ (_06204_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _14561_ (_06205_, _06107_, _06204_);
  and _14562_ (_06206_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _14563_ (_06207_, _06206_, _06205_);
  and _14564_ (_06208_, _06207_, _06203_);
  and _14565_ (_06209_, _06208_, _06198_);
  not _14566_ (_06210_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _14567_ (_06211_, _06088_, _06210_);
  nand _14568_ (_06212_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _14569_ (_06213_, _06212_, _06211_);
  not _14570_ (_06214_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or _14571_ (_06215_, _06083_, _06214_);
  not _14572_ (_06216_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _14573_ (_06217_, _06091_, _06216_);
  and _14574_ (_06218_, _06217_, _06215_);
  and _14575_ (_06219_, _06218_, _06213_);
  or _14576_ (_06220_, _06099_, ABINPUT[2]);
  or _14577_ (_06221_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _14578_ (_06222_, _06221_, _06220_);
  or _14579_ (_06223_, _06222_, _06097_);
  not _14580_ (_06224_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  or _14581_ (_06225_, _06078_, _06224_);
  not _14582_ (_06226_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _14583_ (_06227_, _06107_, _06226_);
  and _14584_ (_06228_, _06227_, _06225_);
  and _14585_ (_06229_, _06228_, _06223_);
  nand _14586_ (_06230_, _06229_, _06219_);
  not _14587_ (_06231_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or _14588_ (_06232_, _06083_, _06231_);
  not _14589_ (_06233_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  or _14590_ (_06234_, _06078_, _06233_);
  and _14591_ (_06235_, _06234_, _06232_);
  nand _14592_ (_06236_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not _14593_ (_06237_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _14594_ (_06238_, _06107_, _06237_);
  and _14595_ (_06239_, _06238_, _06236_);
  and _14596_ (_06240_, _06239_, _06235_);
  not _14597_ (_06241_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _14598_ (_06242_, _06091_, _06241_);
  not _14599_ (_06243_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _14600_ (_06244_, _06088_, _06243_);
  and _14601_ (_06245_, _06244_, _06242_);
  or _14602_ (_06246_, _06099_, ABINPUT[3]);
  or _14603_ (_06247_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _14604_ (_06248_, _06247_, _06246_);
  or _14605_ (_06249_, _06248_, _06097_);
  and _14606_ (_06250_, _06249_, _06245_);
  nand _14607_ (_06251_, _06250_, _06240_);
  nor _14608_ (_06252_, _06251_, _06230_);
  and _14609_ (_06253_, _06252_, _06209_);
  and _14610_ (_06254_, _06253_, _06187_);
  and _14611_ (_06255_, _06254_, _06166_);
  not _14612_ (_06256_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or _14613_ (_06257_, _06078_, _06256_);
  not _14614_ (_06258_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  or _14615_ (_06259_, _06083_, _06258_);
  and _14616_ (_06260_, _06259_, _06257_);
  not _14617_ (_06261_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _14618_ (_06262_, _06088_, _06261_);
  not _14619_ (_06263_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _14620_ (_06264_, _06091_, _06263_);
  and _14621_ (_06265_, _06264_, _06262_);
  and _14622_ (_06266_, _06265_, _06260_);
  or _14623_ (_06267_, _06099_, ABINPUT[7]);
  or _14624_ (_06268_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _14625_ (_06269_, _06268_, _06267_);
  or _14626_ (_06270_, _06269_, _06097_);
  not _14627_ (_06271_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _14628_ (_06272_, _06107_, _06271_);
  nand _14629_ (_06273_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _14630_ (_06274_, _06273_, _06272_);
  and _14631_ (_06275_, _06274_, _06270_);
  and _14632_ (_06276_, _06275_, _06266_);
  not _14633_ (_06277_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  or _14634_ (_06278_, _06083_, _06277_);
  not _14635_ (_06279_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or _14636_ (_06280_, _06078_, _06279_);
  and _14637_ (_06281_, _06280_, _06278_);
  not _14638_ (_06282_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or _14639_ (_06283_, _06091_, _06282_);
  not _14640_ (_06284_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _14641_ (_06285_, _06088_, _06284_);
  and _14642_ (_06286_, _06285_, _06283_);
  and _14643_ (_06287_, _06286_, _06281_);
  or _14644_ (_06288_, _06099_, ABINPUT[6]);
  or _14645_ (_06289_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _14646_ (_06290_, _06289_, _06288_);
  or _14647_ (_06291_, _06290_, _06097_);
  not _14648_ (_06292_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _14649_ (_06293_, _06107_, _06292_);
  nand _14650_ (_06294_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _14651_ (_06295_, _06294_, _06293_);
  and _14652_ (_06296_, _06295_, _06291_);
  nand _14653_ (_06297_, _06296_, _06287_);
  not _14654_ (_06298_, _06297_);
  and _14655_ (_06299_, _06298_, _06276_);
  and _14656_ (_06300_, _06299_, _06255_);
  nor _14657_ (_06301_, _06300_, _06120_);
  not _14658_ (_06302_, _06120_);
  not _14659_ (_06303_, _06276_);
  not _14660_ (_06304_, _06166_);
  not _14661_ (_06305_, _06187_);
  not _14662_ (_06306_, _06209_);
  and _14663_ (_06307_, _06230_, _06306_);
  and _14664_ (_06308_, _06251_, _06307_);
  and _14665_ (_06309_, _06308_, _06305_);
  and _14666_ (_06310_, _06309_, _06304_);
  and _14667_ (_06311_, _06297_, _06310_);
  and _14668_ (_06312_, _06311_, _06303_);
  nor _14669_ (_06313_, _06312_, _06302_);
  or _14670_ (_06314_, _06313_, _06301_);
  and _14671_ (_06315_, _06314_, _06113_);
  nor _14672_ (_06316_, _06314_, _06113_);
  nor _14673_ (_06317_, _06316_, _06315_);
  and _14674_ (_06318_, _06317_, _06145_);
  nor _14675_ (_06319_, _06318_, _06142_);
  and _14676_ (_06320_, _05686_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  nor _14677_ (_06321_, _06320_, _06123_);
  not _14678_ (_06322_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _14679_ (_06323_, _06125_, _06322_);
  and _14680_ (_06324_, _06323_, _06321_);
  and _14681_ (_06325_, _06138_, _06113_);
  nor _14682_ (_06326_, _06138_, _06113_);
  nor _14683_ (_06327_, _06326_, _06325_);
  and _14684_ (_06328_, _06327_, _06324_);
  not _14685_ (_06329_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _14686_ (_06330_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05686_);
  and _14687_ (_06331_, _06330_, _06329_);
  and _14688_ (_06332_, _06331_, _06124_);
  and _14689_ (_06333_, _06332_, _06326_);
  not _14690_ (_06334_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _14691_ (_06335_, _06320_, _06334_);
  and _14692_ (_06336_, _06335_, _06323_);
  not _14693_ (_06337_, _06336_);
  nor _14694_ (_06338_, _06337_, _06325_);
  and _14695_ (_06339_, _06331_, _06144_);
  and _14696_ (_06340_, _06339_, _06113_);
  or _14697_ (_06341_, _06340_, _06338_);
  or _14698_ (_06342_, _06341_, _06333_);
  nor _14699_ (_06343_, _06342_, _06328_);
  nor _14700_ (_06344_, _06330_, _06125_);
  and _14701_ (_06345_, _06344_, _06320_);
  and _14702_ (_06347_, _06331_, _06334_);
  nor _14703_ (_06348_, _06347_, _06345_);
  and _14704_ (_06349_, _06344_, _06321_);
  and _14705_ (_06350_, _06126_, _06334_);
  nor _14706_ (_06351_, _06350_, _06349_);
  and _14707_ (_06352_, _06323_, _06123_);
  not _14708_ (_06353_, _06352_);
  and _14709_ (_06354_, _06353_, _06351_);
  and _14710_ (_06355_, _06354_, _06348_);
  nor _14711_ (_06356_, _06355_, _06113_);
  not _14712_ (_06357_, _06356_);
  and _14713_ (_06358_, _06357_, _06343_);
  and _14714_ (_06359_, _06358_, _06319_);
  not _14715_ (_06360_, _06359_);
  and _14716_ (_06361_, _05993_, _05981_);
  and _14717_ (_06362_, _06361_, _06030_);
  and _14718_ (_06363_, _06362_, _06026_);
  not _14719_ (_06364_, _05923_);
  and _14720_ (_06365_, _05937_, _06364_);
  and _14721_ (_06366_, _05967_, _05954_);
  and _14722_ (_06367_, _06366_, _06365_);
  and _14723_ (_06368_, _06367_, _06363_);
  and _14724_ (_06369_, _06368_, _06011_);
  and _14725_ (_06370_, _06369_, _06360_);
  and _14726_ (_06371_, _06026_, _05981_);
  and _14727_ (_06372_, _06371_, _06005_);
  and _14728_ (_06373_, _06366_, _05938_);
  and _14729_ (_06374_, _06373_, _06372_);
  and _14730_ (_06375_, _06373_, _06363_);
  nor _14731_ (_06376_, _06375_, _06374_);
  and _14732_ (_06377_, _06372_, _06367_);
  not _14733_ (_06378_, _06026_);
  and _14734_ (_06380_, _06362_, _06378_);
  and _14735_ (_06381_, _06380_, _06373_);
  nor _14736_ (_06382_, _06381_, _06377_);
  and _14737_ (_06383_, _06005_, _05981_);
  and _14738_ (_06384_, _06383_, _06378_);
  and _14739_ (_06385_, _06384_, _06373_);
  not _14740_ (_06386_, _06385_);
  and _14741_ (_06387_, _06386_, _06382_);
  and _14742_ (_06388_, _06387_, _06376_);
  not _14743_ (_06389_, _06388_);
  not _14744_ (_06390_, _06011_);
  or _14745_ (_06391_, _06377_, _06368_);
  and _14746_ (_06392_, _06373_, _06361_);
  nor _14747_ (_06393_, _06392_, _06391_);
  or _14748_ (_06394_, _06393_, _06390_);
  or _14749_ (_06395_, _06394_, _06389_);
  and _14750_ (_06396_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or _14751_ (_06397_, _06396_, _06370_);
  and _14752_ (_09300_, _06397_, _06071_);
  and _14753_ (_06398_, _06380_, _06367_);
  and _14754_ (_06399_, _06398_, _06011_);
  not _14755_ (_06400_, _06399_);
  and _14756_ (_06401_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _14757_ (_06402_, _06400_, _06359_);
  or _14758_ (_06403_, _06402_, _06401_);
  and _14759_ (_12917_, _06403_, _06071_);
  or _14760_ (_06404_, _06248_, _06129_);
  or _14761_ (_06405_, _06132_, _06233_);
  or _14762_ (_06406_, _06135_, _06237_);
  and _14763_ (_06407_, _06406_, _06405_);
  nand _14764_ (_06408_, _06407_, _06404_);
  and _14765_ (_06409_, _06408_, _06127_);
  nor _14766_ (_06410_, _06209_, _06120_);
  nor _14767_ (_06411_, _06230_, _06120_);
  nor _14768_ (_06412_, _06411_, _06307_);
  nor _14769_ (_06413_, _06412_, _06410_);
  and _14770_ (_06414_, _06413_, _06251_);
  nor _14771_ (_06415_, _06413_, _06251_);
  nor _14772_ (_06416_, _06415_, _06414_);
  and _14773_ (_06417_, _06416_, _06145_);
  nor _14774_ (_06418_, _06417_, _06409_);
  nor _14775_ (_06419_, _06408_, _06251_);
  nor _14776_ (_06420_, _06419_, _06337_);
  and _14777_ (_06421_, _06408_, _06251_);
  nor _14778_ (_06422_, _06421_, _06419_);
  and _14779_ (_06423_, _06422_, _06324_);
  nor _14780_ (_06424_, _06423_, _06420_);
  and _14781_ (_06425_, _06421_, _06332_);
  not _14782_ (_06426_, _06339_);
  nor _14783_ (_06427_, _06426_, _06251_);
  nor _14784_ (_06428_, _06427_, _06425_);
  not _14785_ (_06429_, _06251_);
  nor _14786_ (_06430_, _06355_, _06429_);
  not _14787_ (_06431_, _06430_);
  and _14788_ (_06432_, _06431_, _06428_);
  and _14789_ (_06433_, _06432_, _06424_);
  and _14790_ (_06434_, _06433_, _06418_);
  not _14791_ (_06435_, _06434_);
  and _14792_ (_06436_, _06435_, _06377_);
  not _14793_ (_06437_, _06392_);
  nor _14794_ (_06438_, _06388_, _06390_);
  nand _14795_ (_06439_, _06438_, _06437_);
  and _14796_ (_06440_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _14797_ (_06441_, _06440_, _06436_);
  or _14798_ (_06442_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _14799_ (_06443_, _06442_, _06071_);
  and _14800_ (_12997_, _06443_, _06441_);
  not _14801_ (_06444_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _14802_ (_06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14803_ (_06446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _06445_);
  and _14804_ (_06447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14805_ (_06448_, _06447_, _06446_);
  and _14806_ (_06449_, _06448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _14807_ (_06450_, _06449_, _06444_);
  and _14808_ (_06451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _14809_ (_06452_, _06451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _14810_ (_06453_, _06452_);
  and _14811_ (_06454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _14812_ (_06455_, _06454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14813_ (_06456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14814_ (_06457_, _06456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor _14815_ (_06458_, _06457_, _06455_);
  and _14816_ (_06459_, _06458_, _06453_);
  nor _14817_ (_06460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  not _14818_ (_06461_, _06460_);
  and _14819_ (_06462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _14820_ (_06463_, _06462_, _06461_);
  not _14821_ (_06464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _14822_ (_06465_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _14823_ (_06466_, _06465_, _06464_);
  and _14824_ (_06467_, _06466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _14825_ (_06468_, _06467_, _06463_);
  and _14826_ (_06469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _14827_ (_06470_, _06469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _14828_ (_06471_, _06470_);
  and _14829_ (_06472_, _06471_, _06468_);
  and _14830_ (_06473_, _06472_, _06459_);
  nor _14831_ (_06474_, _06473_, _06450_);
  and _14832_ (_06475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _06444_);
  not _14833_ (_06476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _14834_ (_06477_, _06476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _14835_ (_06478_, _06477_, _06461_);
  not _14836_ (_06479_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _14837_ (_06480_, _06466_, _06479_);
  nor _14838_ (_06481_, _06480_, _06478_);
  not _14839_ (_06482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _14840_ (_06483_, _06469_, _06482_);
  not _14841_ (_06484_, _06483_);
  nand _14842_ (_06485_, _06484_, _06481_);
  and _14843_ (_06486_, _06485_, _06475_);
  or _14844_ (_06487_, _06486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not _14845_ (_06488_, _06475_);
  not _14846_ (_06489_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _14847_ (_06490_, _06451_, _06489_);
  not _14848_ (_06491_, _06490_);
  not _14849_ (_06492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14850_ (_06493_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _14851_ (_06494_, _06493_, _06492_);
  not _14852_ (_06495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14853_ (_06496_, _06454_, _06495_);
  nor _14854_ (_06497_, _06496_, _06494_);
  and _14855_ (_06498_, _06497_, _06491_);
  or _14856_ (_06499_, _06498_, _06488_);
  or _14857_ (_06500_, _06499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14858_ (_06501_, _06500_, _06487_);
  or _14859_ (_06502_, _06501_, _06474_);
  not _14860_ (_06503_, _06472_);
  or _14861_ (_06504_, _06459_, _06450_);
  or _14862_ (_06505_, _06504_, _06503_);
  and _14863_ (_06506_, _06505_, _06445_);
  or _14864_ (_06507_, _06506_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _14865_ (_06508_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _14866_ (_06509_, _06508_);
  and _14867_ (_06510_, _06509_, _06504_);
  nor _14868_ (_06511_, _06508_, _06445_);
  or _14869_ (_06512_, _06511_, _06510_);
  and _14870_ (_06513_, _06512_, _06507_);
  and _14871_ (_06514_, _06513_, _06502_);
  and _14872_ (_06515_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _14873_ (_06516_, _06515_, _06514_);
  and _14874_ (_00316_, _06516_, _06071_);
  and _14875_ (_06517_, _06498_, _06484_);
  nand _14876_ (_06518_, _06517_, _06481_);
  and _14877_ (_06519_, _06518_, _06475_);
  nand _14878_ (_06520_, _06473_, _06444_);
  or _14879_ (_06521_, _06520_, _06519_);
  nor _14880_ (_06522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06445_);
  nand _14881_ (_06523_, _06522_, _06508_);
  and _14882_ (_06524_, _06523_, _06071_);
  and _14883_ (_00503_, _06524_, _06521_);
  and _14884_ (_06525_, _05704_, _05694_);
  nor _14885_ (_06526_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and _14886_ (_06527_, _06526_, _05686_);
  not _14887_ (_06528_, _06527_);
  nor _14888_ (_06529_, _06528_, _06525_);
  nor _14889_ (_06530_, _06529_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _14890_ (_06531_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not _14891_ (_06532_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _14892_ (_06533_, _06530_, _06532_);
  and _14893_ (_06534_, _06533_, _06071_);
  and _14894_ (_00572_, _06534_, _06531_);
  and _14895_ (_06535_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _14896_ (_06536_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _14897_ (_06537_, _06059_, _06044_);
  and _14898_ (_06538_, _06537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _14899_ (_06539_, _06046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _14900_ (_06540_, _06539_, _06538_);
  and _14901_ (_06541_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _14902_ (_06542_, _06541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _14903_ (_06543_, _06540_, _06047_);
  and _14904_ (_06544_, _06543_, _06542_);
  and _14905_ (_06545_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _14906_ (_06546_, _06545_);
  and _14907_ (_06547_, _06546_, _06053_);
  and _14908_ (_06548_, _06547_, _06059_);
  and _14909_ (_06549_, _06548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _14910_ (_06550_, _06549_, _06065_);
  or _14911_ (_06551_, _06550_, _06544_);
  and _14912_ (_06552_, _06551_, _06536_);
  and _14913_ (_06553_, _06552_, _06036_);
  or _14914_ (_06554_, _06553_, _06535_);
  not _14915_ (_06555_, _06035_);
  nor _14916_ (_06556_, _06359_, _06555_);
  or _14917_ (_06557_, _06556_, _06554_);
  and _14918_ (_01048_, _06557_, _06071_);
  nor _14919_ (_06558_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _14920_ (_06559_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _14921_ (_06560_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _14922_ (_06561_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _14923_ (_01756_, _06561_, _06559_);
  nor _14924_ (_06562_, _06519_, _06474_);
  and _14925_ (_06563_, _06562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not _14926_ (_06564_, _06474_);
  and _14927_ (_06565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06445_);
  nor _14928_ (_06566_, _06565_, _06522_);
  nor _14929_ (_06567_, _06566_, _06564_);
  or _14930_ (_06568_, _06567_, _06508_);
  or _14931_ (_06569_, _06568_, _06563_);
  or _14932_ (_06570_, _06566_, _06509_);
  and _14933_ (_06571_, _06570_, _06071_);
  and _14934_ (_01890_, _06571_, _06569_);
  and _14935_ (_06572_, _06297_, _06120_);
  or _14936_ (_06573_, _06290_, _06129_);
  or _14937_ (_06574_, _06132_, _06279_);
  or _14938_ (_06575_, _06135_, _06292_);
  and _14939_ (_06576_, _06575_, _06574_);
  and _14940_ (_06577_, _06576_, _06573_);
  nor _14941_ (_06578_, _06577_, _06120_);
  or _14942_ (_06579_, _06578_, _06572_);
  and _14943_ (_06580_, _06579_, _06127_);
  and _14944_ (_06581_, _06310_, _06120_);
  and _14945_ (_06582_, _06255_, _06302_);
  nor _14946_ (_06583_, _06582_, _06581_);
  and _14947_ (_06584_, _06583_, _06298_);
  not _14948_ (_06585_, _06145_);
  nor _14949_ (_06586_, _06583_, _06298_);
  or _14950_ (_06587_, _06586_, _06585_);
  nor _14951_ (_06588_, _06587_, _06584_);
  nor _14952_ (_06590_, _06588_, _06580_);
  nor _14953_ (_06591_, _06355_, _06298_);
  not _14954_ (_06592_, _06591_);
  nand _14955_ (_06593_, _06576_, _06573_);
  and _14956_ (_06594_, _06593_, _06297_);
  nor _14957_ (_06595_, _06593_, _06297_);
  nor _14958_ (_06596_, _06595_, _06594_);
  and _14959_ (_06597_, _06596_, _06324_);
  not _14960_ (_06598_, _06597_);
  nor _14961_ (_06599_, _06595_, _06337_);
  not _14962_ (_06600_, _06599_);
  and _14963_ (_06601_, _06594_, _06332_);
  nor _14964_ (_06602_, _06426_, _06297_);
  nor _14965_ (_06603_, _06602_, _06601_);
  and _14966_ (_06605_, _06603_, _06600_);
  and _14967_ (_06607_, _06605_, _06598_);
  and _14968_ (_06608_, _06607_, _06592_);
  and _14969_ (_06609_, _06608_, _06590_);
  and _14970_ (_06610_, _06385_, _06011_);
  not _14971_ (_06611_, _06610_);
  nor _14972_ (_06612_, _06611_, _06609_);
  and _14973_ (_06613_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _14974_ (_06614_, _06613_, _06612_);
  and _14975_ (_02186_, _06614_, _06071_);
  and _14976_ (_06615_, _06344_, _06144_);
  not _14977_ (_06616_, _06615_);
  and _14978_ (_06618_, _06139_, _06113_);
  or _14979_ (_06619_, _06269_, _06129_);
  or _14980_ (_06620_, _06132_, _06256_);
  or _14981_ (_06621_, _06135_, _06271_);
  and _14982_ (_06622_, _06621_, _06620_);
  nand _14983_ (_06623_, _06622_, _06619_);
  nor _14984_ (_06624_, _06623_, _06276_);
  not _14985_ (_06625_, _06623_);
  nor _14986_ (_06626_, _06625_, _06276_);
  and _14987_ (_06627_, _06625_, _06276_);
  nor _14988_ (_06628_, _06627_, _06626_);
  and _14989_ (_06629_, _06577_, _06297_);
  or _14990_ (_06630_, _06159_, _06129_);
  or _14991_ (_06631_, _06132_, _06146_);
  or _14992_ (_06632_, _06135_, _06161_);
  and _14993_ (_06633_, _06632_, _06631_);
  nand _14994_ (_06634_, _06633_, _06630_);
  and _14995_ (_06635_, _06634_, _06166_);
  nor _14996_ (_06636_, _06635_, _06596_);
  nor _14997_ (_06637_, _06636_, _06629_);
  nor _14998_ (_06638_, _06637_, _06628_);
  nor _14999_ (_06639_, _06638_, _06624_);
  and _15000_ (_06640_, _06637_, _06628_);
  nor _15001_ (_06641_, _06640_, _06638_);
  not _15002_ (_06642_, _06641_);
  and _15003_ (_06643_, _06635_, _06596_);
  nor _15004_ (_06644_, _06643_, _06636_);
  not _15005_ (_06645_, _06644_);
  and _15006_ (_06646_, _06633_, _06630_);
  nor _15007_ (_06647_, _06646_, _06166_);
  and _15008_ (_06648_, _06646_, _06166_);
  nor _15009_ (_06649_, _06648_, _06647_);
  not _15010_ (_06650_, _06649_);
  or _15011_ (_06651_, _06180_, _06129_);
  or _15012_ (_06652_, _06132_, _06169_);
  or _15013_ (_06653_, _06135_, _06183_);
  and _15014_ (_06654_, _06653_, _06652_);
  and _15015_ (_06655_, _06654_, _06651_);
  and _15016_ (_06656_, _06655_, _06187_);
  nor _15017_ (_06657_, _06655_, _06187_);
  nor _15018_ (_06659_, _06657_, _06656_);
  and _15019_ (_06660_, _06407_, _06404_);
  and _15020_ (_06661_, _06660_, _06251_);
  or _15021_ (_06662_, _06222_, _06129_);
  or _15022_ (_06663_, _06132_, _06224_);
  or _15023_ (_06664_, _06135_, _06226_);
  and _15024_ (_06665_, _06664_, _06663_);
  nand _15025_ (_06666_, _06665_, _06662_);
  and _15026_ (_06667_, _06666_, _06230_);
  nor _15027_ (_06668_, _06666_, _06230_);
  nor _15028_ (_06669_, _06668_, _06667_);
  or _15029_ (_06670_, _06202_, _06129_);
  or _15030_ (_06671_, _06132_, _06188_);
  or _15031_ (_06672_, _06135_, _06204_);
  and _15032_ (_06673_, _06672_, _06671_);
  nand _15033_ (_06674_, _06673_, _06670_);
  and _15034_ (_06675_, _06674_, _06209_);
  nor _15035_ (_06676_, _06675_, _06669_);
  and _15036_ (_06677_, _06665_, _06662_);
  and _15037_ (_06678_, _06677_, _06230_);
  nor _15038_ (_06680_, _06678_, _06676_);
  nor _15039_ (_06681_, _06680_, _06422_);
  nor _15040_ (_06682_, _06681_, _06661_);
  nor _15041_ (_06683_, _06682_, _06659_);
  and _15042_ (_06684_, _06682_, _06659_);
  nor _15043_ (_06685_, _06684_, _06683_);
  and _15044_ (_06686_, _06680_, _06422_);
  nor _15045_ (_06687_, _06686_, _06681_);
  and _15046_ (_06688_, _06675_, _06669_);
  nor _15047_ (_06689_, _06688_, _06676_);
  and _15048_ (_06690_, _06673_, _06670_);
  nor _15049_ (_06691_, _06690_, _06209_);
  and _15050_ (_06692_, _06690_, _06209_);
  nor _15051_ (_06693_, _06692_, _06691_);
  nor _15052_ (_06694_, _06693_, _06120_);
  not _15053_ (_06695_, _06694_);
  nor _15054_ (_06696_, _06695_, _06689_);
  not _15055_ (_06697_, _06696_);
  nor _15056_ (_06698_, _06697_, _06687_);
  not _15057_ (_06699_, _06698_);
  nor _15058_ (_06700_, _06699_, _06685_);
  nand _15059_ (_06701_, _06654_, _06651_);
  or _15060_ (_06702_, _06701_, _06187_);
  and _15061_ (_06703_, _06701_, _06187_);
  or _15062_ (_06704_, _06682_, _06703_);
  and _15063_ (_06705_, _06704_, _06702_);
  or _15064_ (_06706_, _06705_, _06700_);
  and _15065_ (_06707_, _06706_, _06650_);
  and _15066_ (_06708_, _06707_, _06645_);
  and _15067_ (_06709_, _06708_, _06642_);
  nor _15068_ (_06710_, _06709_, _06639_);
  nor _15069_ (_06711_, _06710_, _06327_);
  nor _15070_ (_06712_, _06711_, _06618_);
  nor _15071_ (_06713_, _06712_, _06616_);
  not _15072_ (_06714_, _06713_);
  and _15073_ (_06715_, _06344_, _06335_);
  not _15074_ (_06716_, _06715_);
  not _15075_ (_06717_, _06326_);
  not _15076_ (_06718_, _06422_);
  and _15077_ (_06719_, _06691_, _06669_);
  nor _15078_ (_06720_, _06719_, _06667_);
  nor _15079_ (_06721_, _06720_, _06718_);
  nor _15080_ (_06722_, _06721_, _06421_);
  nor _15081_ (_06723_, _06722_, _06659_);
  and _15082_ (_06724_, _06722_, _06659_);
  nor _15083_ (_06725_, _06724_, _06723_);
  and _15084_ (_06726_, _06693_, _06302_);
  and _15085_ (_06727_, _06726_, _06669_);
  and _15086_ (_06728_, _06720_, _06718_);
  nor _15087_ (_06729_, _06728_, _06721_);
  and _15088_ (_06730_, _06729_, _06727_);
  not _15089_ (_06731_, _06730_);
  nor _15090_ (_06732_, _06731_, _06725_);
  nor _15091_ (_06733_, _06722_, _06656_);
  or _15092_ (_06734_, _06733_, _06657_);
  or _15093_ (_06735_, _06734_, _06732_);
  and _15094_ (_06736_, _06735_, _06649_);
  and _15095_ (_06737_, _06736_, _06596_);
  not _15096_ (_06738_, _06628_);
  and _15097_ (_06739_, _06647_, _06596_);
  nor _15098_ (_06740_, _06739_, _06594_);
  nor _15099_ (_06741_, _06740_, _06738_);
  and _15100_ (_06742_, _06740_, _06738_);
  nor _15101_ (_06743_, _06742_, _06741_);
  and _15102_ (_06744_, _06743_, _06737_);
  not _15103_ (_06745_, _06744_);
  nor _15104_ (_06746_, _06741_, _06626_);
  and _15105_ (_06747_, _06746_, _06745_);
  or _15106_ (_06748_, _06747_, _06325_);
  and _15107_ (_06749_, _06748_, _06717_);
  nor _15108_ (_06750_, _06749_, _06716_);
  and _15109_ (_06751_, _06335_, _06331_);
  nor _15110_ (_06752_, _06252_, _06187_);
  and _15111_ (_06753_, _06752_, _06751_);
  and _15112_ (_06754_, _06753_, _06304_);
  nor _15113_ (_06755_, _06754_, _06297_);
  and _15114_ (_06756_, _06276_, _06120_);
  and _15115_ (_06757_, _06756_, _06755_);
  nor _15116_ (_06758_, _06757_, _06121_);
  not _15117_ (_06759_, _06751_);
  and _15118_ (_06760_, _06755_, _06276_);
  nor _15119_ (_06761_, _06120_, _06113_);
  not _15120_ (_06762_, _06761_);
  nor _15121_ (_06763_, _06762_, _06760_);
  nor _15122_ (_06764_, _06763_, _06759_);
  and _15123_ (_06765_, _06764_, _06758_);
  not _15124_ (_06766_, _06118_);
  nor _15125_ (_06767_, _06753_, _06302_);
  and _15126_ (_06768_, _06767_, _06766_);
  nor _15127_ (_06769_, _06115_, _06766_);
  not _15128_ (_06770_, _06324_);
  nor _15129_ (_06771_, _06770_, _06769_);
  nor _15130_ (_06772_, _06771_, _06336_);
  not _15131_ (_06773_, _06772_);
  nor _15132_ (_06774_, _06773_, _06753_);
  nor _15133_ (_06775_, _06774_, _06768_);
  not _15134_ (_06776_, _06113_);
  and _15135_ (_06777_, _06323_, _06124_);
  and _15136_ (_06779_, _06777_, _06776_);
  and _15137_ (_06780_, _06115_, _06118_);
  and _15138_ (_06781_, _06323_, _06144_);
  and _15139_ (_06782_, _06332_, _06118_);
  nor _15140_ (_06784_, _06782_, _06781_);
  nor _15141_ (_06785_, _06784_, _06780_);
  nor _15142_ (_06786_, _06785_, _06779_);
  and _15143_ (_06787_, _06335_, _06126_);
  and _15144_ (_06788_, _06787_, _06306_);
  and _15145_ (_06789_, _06321_, _06126_);
  and _15146_ (_06790_, _06789_, _06766_);
  nor _15147_ (_06791_, _06790_, _06349_);
  and _15148_ (_06792_, _06791_, _06302_);
  and _15149_ (_06793_, _06426_, _06120_);
  nor _15150_ (_06794_, _06793_, _06792_);
  nor _15151_ (_06795_, _06794_, _06788_);
  and _15152_ (_06796_, _06795_, _06786_);
  not _15153_ (_06797_, _06796_);
  nor _15154_ (_06798_, _06797_, _06775_);
  not _15155_ (_06799_, _06798_);
  nor _15156_ (_06800_, _06799_, _06765_);
  not _15157_ (_06801_, _06800_);
  nor _15158_ (_06802_, _06801_, _06750_);
  and _15159_ (_06803_, _06802_, _06714_);
  nor _15160_ (_06804_, _06004_, _05993_);
  and _15161_ (_06805_, _06804_, _05982_);
  and _15162_ (_06806_, _05954_, _05937_);
  not _15163_ (_06807_, _05967_);
  nor _15164_ (_06808_, _06378_, _05923_);
  and _15165_ (_06809_, _06808_, _06807_);
  and _15166_ (_06810_, _06809_, _06806_);
  and _15167_ (_06812_, _06810_, _06805_);
  nand _15168_ (_06813_, _06812_, _06803_);
  and _15169_ (_06814_, _06010_, _06008_);
  and _15170_ (_06815_, _06814_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or _15171_ (_06816_, _06812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _15172_ (_06817_, _06816_, _06815_);
  and _15173_ (_06818_, _06817_, _06813_);
  not _15174_ (_06819_, _05954_);
  nor _15175_ (_06820_, _05967_, _06819_);
  and _15176_ (_06821_, _06820_, _06365_);
  and _15177_ (_06822_, _06821_, _06372_);
  nand _15178_ (_06823_, _06822_, _06359_);
  or _15179_ (_06824_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _15180_ (_06825_, _06824_, _06012_);
  and _15181_ (_06826_, _06825_, _06823_);
  not _15182_ (_06827_, _06814_);
  and _15183_ (_06828_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _15184_ (_06829_, _06828_, rst);
  or _15185_ (_06830_, _06829_, _06826_);
  or _15186_ (_03745_, _06830_, _06818_);
  nor _15187_ (_06831_, t2ex_i, rst);
  and _15188_ (_04082_, _06831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  and _15189_ (_06832_, _06026_, _05923_);
  and _15190_ (_06833_, _06832_, _06807_);
  and _15191_ (_06834_, _06833_, _06806_);
  and _15192_ (_06835_, _06834_, _06805_);
  nand _15193_ (_06836_, _06835_, _06803_);
  or _15194_ (_06837_, _06835_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _15195_ (_06838_, _06837_, _06815_);
  and _15196_ (_06839_, _06838_, _06836_);
  and _15197_ (_06840_, _06820_, _05938_);
  and _15198_ (_06841_, _06840_, _06372_);
  nand _15199_ (_06842_, _06841_, _06359_);
  or _15200_ (_06843_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _15201_ (_06844_, _06843_, _06012_);
  and _15202_ (_06845_, _06844_, _06842_);
  and _15203_ (_06846_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _15204_ (_06847_, _06846_, rst);
  or _15205_ (_06848_, _06847_, _06845_);
  or _15206_ (_05680_, _06848_, _06839_);
  or _15207_ (_06849_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not _15208_ (_06850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _15209_ (_06851_, _06530_, _06850_);
  and _15210_ (_06852_, _06851_, _06071_);
  and _15211_ (_05681_, _06852_, _06849_);
  nor _15212_ (_06853_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _15213_ (_06854_, _06853_);
  and _15214_ (_06855_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  not _15215_ (_06856_, _06230_);
  not _15216_ (_06857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _15217_ (_06858_, _06857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _15218_ (_06859_, _06858_);
  or _15219_ (_06860_, _06859_, _06660_);
  not _15220_ (_06861_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _15221_ (_06862_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _06861_);
  not _15222_ (_06863_, _06862_);
  or _15223_ (_06864_, _06863_, _06646_);
  and _15224_ (_06865_, _06864_, _06860_);
  or _15225_ (_06866_, _06862_, _06858_);
  or _15226_ (_06867_, _06866_, _06690_);
  and _15227_ (_06868_, _06867_, _06854_);
  nand _15228_ (_06869_, _06868_, _06865_);
  or _15229_ (_06870_, _06854_, _06623_);
  nand _15230_ (_06871_, _06870_, _06869_);
  or _15231_ (_06872_, _06871_, _06856_);
  or _15232_ (_06873_, _06859_, _06655_);
  or _15233_ (_06874_, _06863_, _06577_);
  and _15234_ (_06875_, _06874_, _06873_);
  or _15235_ (_06876_, _06866_, _06677_);
  and _15236_ (_06877_, _06876_, _06854_);
  nand _15237_ (_06878_, _06877_, _06875_);
  nand _15238_ (_06879_, _06853_, _06138_);
  nand _15239_ (_06880_, _06879_, _06878_);
  or _15240_ (_06881_, _06880_, _06209_);
  nor _15241_ (_06882_, _06881_, _06872_);
  and _15242_ (_06883_, _06879_, _06878_);
  and _15243_ (_06884_, _06883_, _06230_);
  and _15244_ (_06885_, _06870_, _06869_);
  and _15245_ (_06886_, _06885_, _06251_);
  nand _15246_ (_06887_, _06886_, _06884_);
  or _15247_ (_06888_, _06886_, _06884_);
  and _15248_ (_06889_, _06888_, _06887_);
  and _15249_ (_06890_, _06889_, _06882_);
  and _15250_ (_06891_, _06885_, _06305_);
  and _15251_ (_06892_, _06883_, _06251_);
  and _15252_ (_06893_, _06892_, _06872_);
  nand _15253_ (_06894_, _06893_, _06891_);
  or _15254_ (_06895_, _06893_, _06891_);
  and _15255_ (_06896_, _06895_, _06894_);
  and _15256_ (_06897_, _06896_, _06890_);
  nand _15257_ (_06898_, _06894_, _06887_);
  or _15258_ (_06899_, _06880_, _06187_);
  or _15259_ (_06900_, _06871_, _06166_);
  or _15260_ (_06901_, _06900_, _06899_);
  nand _15261_ (_06902_, _06900_, _06899_);
  and _15262_ (_06903_, _06902_, _06901_);
  nand _15263_ (_06904_, _06903_, _06898_);
  or _15264_ (_06905_, _06903_, _06898_);
  and _15265_ (_06906_, _06905_, _06904_);
  nand _15266_ (_06907_, _06906_, _06897_);
  or _15267_ (_06908_, _06906_, _06897_);
  and _15268_ (_06910_, _06908_, _06907_);
  nand _15269_ (_06911_, _06910_, _06855_);
  and _15270_ (_06912_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand _15271_ (_06913_, _06896_, _06890_);
  or _15272_ (_06914_, _06896_, _06890_);
  and _15273_ (_06915_, _06914_, _06913_);
  nand _15274_ (_06916_, _06915_, _06912_);
  and _15275_ (_06917_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _15276_ (_06918_, _06889_, _06882_);
  nor _15277_ (_06919_, _06918_, _06890_);
  nand _15278_ (_06920_, _06919_, _06917_);
  or _15279_ (_06921_, _06915_, _06912_);
  nand _15280_ (_06922_, _06921_, _06916_);
  or _15281_ (_06923_, _06922_, _06920_);
  and _15282_ (_06924_, _06923_, _06916_);
  or _15283_ (_06925_, _06910_, _06855_);
  nand _15284_ (_06926_, _06925_, _06911_);
  or _15285_ (_06927_, _06926_, _06924_);
  and _15286_ (_06928_, _06927_, _06911_);
  and _15287_ (_06929_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  and _15288_ (_06930_, _06906_, _06897_);
  and _15289_ (_06931_, _06903_, _06898_);
  and _15290_ (_06932_, _06883_, _06304_);
  and _15291_ (_06933_, _06932_, _06891_);
  or _15292_ (_06934_, _06880_, _06298_);
  or _15293_ (_06935_, _06934_, _06900_);
  and _15294_ (_06936_, _06885_, _06297_);
  or _15295_ (_06937_, _06936_, _06932_);
  and _15296_ (_06938_, _06937_, _06935_);
  nand _15297_ (_06939_, _06938_, _06933_);
  or _15298_ (_06940_, _06938_, _06933_);
  and _15299_ (_06941_, _06940_, _06939_);
  nand _15300_ (_06942_, _06941_, _06931_);
  or _15301_ (_06943_, _06941_, _06931_);
  and _15302_ (_06944_, _06943_, _06942_);
  nand _15303_ (_06945_, _06944_, _06930_);
  or _15304_ (_06946_, _06944_, _06930_);
  and _15305_ (_06947_, _06946_, _06945_);
  nand _15306_ (_06948_, _06947_, _06929_);
  or _15307_ (_06949_, _06947_, _06929_);
  nand _15308_ (_06951_, _06949_, _06948_);
  or _15309_ (_06952_, _06951_, _06928_);
  not _15310_ (_06954_, _06952_);
  and _15311_ (_06955_, _06951_, _06928_);
  nor _15312_ (_06956_, _06955_, _06954_);
  and _15313_ (_05682_, _06956_, _06071_);
  or _15314_ (_06957_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not _15315_ (_06958_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _15316_ (_06959_, _06530_, _06958_);
  and _15317_ (_06960_, _06959_, _06071_);
  and _15318_ (_05683_, _06960_, _06957_);
  or _15319_ (_06961_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not _15320_ (_06962_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _15321_ (_06963_, _06530_, _06962_);
  and _15322_ (_06964_, _06963_, _06071_);
  and _15323_ (_05684_, _06964_, _06961_);
  and _15324_ (_06965_, _06384_, _06367_);
  and _15325_ (_06966_, _06965_, _06011_);
  not _15326_ (_06967_, _06966_);
  and _15327_ (_06968_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor _15328_ (_06969_, _06166_, _06302_);
  nor _15329_ (_06970_, _06646_, _06120_);
  or _15330_ (_06971_, _06970_, _06969_);
  and _15331_ (_06972_, _06971_, _06127_);
  nor _15332_ (_06973_, _06309_, _06302_);
  nor _15333_ (_06974_, _06254_, _06120_);
  nor _15334_ (_06975_, _06974_, _06973_);
  and _15335_ (_06976_, _06975_, _06304_);
  nor _15336_ (_06977_, _06975_, _06304_);
  nor _15337_ (_06978_, _06977_, _06976_);
  and _15338_ (_06979_, _06978_, _06145_);
  nor _15339_ (_06980_, _06979_, _06972_);
  nor _15340_ (_06981_, _06355_, _06166_);
  not _15341_ (_06982_, _06981_);
  and _15342_ (_06983_, _06649_, _06324_);
  not _15343_ (_06984_, _06983_);
  nor _15344_ (_06985_, _06648_, _06337_);
  not _15345_ (_06986_, _06985_);
  and _15346_ (_06987_, _06647_, _06332_);
  and _15347_ (_06988_, _06339_, _06166_);
  nor _15348_ (_06989_, _06988_, _06987_);
  and _15349_ (_06990_, _06989_, _06986_);
  and _15350_ (_06991_, _06990_, _06984_);
  and _15351_ (_06992_, _06991_, _06982_);
  and _15352_ (_06993_, _06992_, _06980_);
  nor _15353_ (_06994_, _06993_, _06967_);
  or _15354_ (_06995_, _06994_, _06968_);
  and _15355_ (_05750_, _06995_, _06071_);
  not _15356_ (_06996_, _06375_);
  nor _15357_ (_06997_, _06434_, _06996_);
  and _15358_ (_06998_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _15359_ (_06999_, _06998_, _06390_);
  or _15360_ (_07000_, _06999_, _06997_);
  or _15361_ (_07001_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _15362_ (_07002_, _07001_, _06071_);
  and _15363_ (_05935_, _07002_, _07000_);
  and _15364_ (_07003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _06071_);
  not _15365_ (_07004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor _15366_ (_07005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor _15367_ (_07006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _15368_ (_07007_, _07006_, _07005_);
  or _15369_ (_07008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _15370_ (_07009_, _07008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _15371_ (_07010_, _07009_, _07007_);
  and _15372_ (_07011_, _07010_, _07004_);
  and _15373_ (_07012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _06071_);
  and _15374_ (_07013_, _07012_, _07011_);
  or _15375_ (_05942_, _07013_, _07003_);
  and _15376_ (_07014_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _15377_ (_07015_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _15378_ (_07016_, _06939_);
  not _15379_ (_07017_, _06934_);
  and _15380_ (_07018_, _06885_, _06303_);
  not _15381_ (_07019_, _07018_);
  nand _15382_ (_07020_, _07019_, _06935_);
  or _15383_ (_07021_, _06935_, _06276_);
  and _15384_ (_07022_, _07021_, _07020_);
  nand _15385_ (_07023_, _07022_, _07017_);
  or _15386_ (_07024_, _07018_, _07017_);
  and _15387_ (_07025_, _07024_, _07023_);
  and _15388_ (_07026_, _07025_, _07016_);
  or _15389_ (_07027_, _06871_, _06113_);
  or _15390_ (_07028_, _06880_, _06276_);
  or _15391_ (_07029_, _07028_, _07027_);
  nand _15392_ (_07030_, _07028_, _07027_);
  and _15393_ (_07031_, _07030_, _07029_);
  not _15394_ (_07032_, _07031_);
  or _15395_ (_07033_, _07032_, _07021_);
  or _15396_ (_07034_, _07032_, _07023_);
  nand _15397_ (_07035_, _07032_, _07023_);
  nand _15398_ (_07036_, _07035_, _07034_);
  nand _15399_ (_07037_, _07036_, _07021_);
  and _15400_ (_07038_, _07037_, _07033_);
  nand _15401_ (_07039_, _07038_, _07026_);
  or _15402_ (_07040_, _07038_, _07026_);
  and _15403_ (_07041_, _07040_, _07039_);
  nand _15404_ (_07042_, _07024_, _07023_);
  or _15405_ (_07043_, _07042_, _06942_);
  not _15406_ (_07044_, _06945_);
  and _15407_ (_07045_, _06942_, _06939_);
  nand _15408_ (_07046_, _07045_, _07042_);
  or _15409_ (_07047_, _07045_, _07042_);
  and _15410_ (_07048_, _07047_, _07046_);
  nand _15411_ (_07049_, _07048_, _07044_);
  nand _15412_ (_07050_, _07049_, _07043_);
  nand _15413_ (_07051_, _07050_, _07041_);
  nand _15414_ (_07053_, _07051_, _07039_);
  and _15415_ (_07054_, _06883_, _06776_);
  and _15416_ (_07055_, _07054_, _07019_);
  and _15417_ (_07056_, _07033_, _07034_);
  not _15418_ (_07057_, _07056_);
  nand _15419_ (_07058_, _07057_, _07055_);
  or _15420_ (_07059_, _07057_, _07055_);
  and _15421_ (_07060_, _07059_, _07058_);
  nand _15422_ (_07061_, _07060_, _07053_);
  and _15423_ (_07062_, _07058_, _07029_);
  nand _15424_ (_07063_, _07062_, _07061_);
  nand _15425_ (_07064_, _07063_, _07015_);
  or _15426_ (_07065_, _07063_, _07015_);
  nand _15427_ (_07067_, _07065_, _07064_);
  and _15428_ (_07068_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or _15429_ (_07070_, _07060_, _07053_);
  and _15430_ (_07071_, _07070_, _07061_);
  nand _15431_ (_07073_, _07071_, _07068_);
  and _15432_ (_07075_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or _15433_ (_07076_, _07050_, _07041_);
  and _15434_ (_07078_, _07076_, _07051_);
  nand _15435_ (_07079_, _07078_, _07075_);
  or _15436_ (_07081_, _07078_, _07075_);
  nand _15437_ (_07083_, _07081_, _07079_);
  and _15438_ (_07084_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or _15439_ (_07085_, _07048_, _07044_);
  and _15440_ (_07086_, _07085_, _07049_);
  nand _15441_ (_07087_, _07086_, _07084_);
  or _15442_ (_07088_, _07086_, _07084_);
  nand _15443_ (_07089_, _07088_, _07087_);
  and _15444_ (_07090_, _06952_, _06948_);
  or _15445_ (_07091_, _07090_, _07089_);
  and _15446_ (_07092_, _07091_, _07087_);
  or _15447_ (_07093_, _07092_, _07083_);
  and _15448_ (_07094_, _07093_, _07079_);
  or _15449_ (_07095_, _07071_, _07068_);
  nand _15450_ (_07096_, _07095_, _07073_);
  or _15451_ (_07097_, _07096_, _07094_);
  and _15452_ (_07098_, _07097_, _07073_);
  or _15453_ (_07099_, _07098_, _07067_);
  nand _15454_ (_07100_, _07099_, _07064_);
  nand _15455_ (_07101_, _07100_, _07014_);
  or _15456_ (_07102_, _07100_, _07014_);
  and _15457_ (_07103_, _07102_, _07101_);
  and _15458_ (_05974_, _07103_, _06071_);
  and _15459_ (_07104_, _06026_, _06012_);
  and _15460_ (_07105_, _06804_, _05981_);
  and _15461_ (_07106_, _06840_, _07105_);
  nand _15462_ (_07107_, _07106_, _07104_);
  and _15463_ (_07108_, _06331_, _06321_);
  and _15464_ (_07109_, _06625_, _06138_);
  nor _15465_ (_07110_, _07109_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _15466_ (_07112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15467_ (_07113_, _06634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _15468_ (_07114_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15469_ (_07115_, _06623_, _07114_);
  nand _15470_ (_07116_, _07115_, _07113_);
  or _15471_ (_07117_, _06593_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15472_ (_07118_, _06138_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15473_ (_07119_, _07118_, _07117_);
  and _15474_ (_07120_, _07119_, _07116_);
  or _15475_ (_07121_, _06701_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15476_ (_07122_, _06593_, _07114_);
  nand _15477_ (_07123_, _07122_, _07121_);
  or _15478_ (_07124_, _06408_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15479_ (_07126_, _06634_, _07114_);
  nand _15480_ (_07127_, _07126_, _07124_);
  and _15481_ (_07128_, _07127_, _07123_);
  nand _15482_ (_07129_, _07128_, _07120_);
  and _15483_ (_07130_, _07129_, _07112_);
  nor _15484_ (_07132_, _07130_, _07110_);
  or _15485_ (_07133_, _06666_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15486_ (_07134_, _06701_, _07114_);
  nand _15487_ (_07135_, _07134_, _07133_);
  and _15488_ (_07136_, _07135_, _07112_);
  and _15489_ (_07137_, _07119_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15490_ (_07138_, _07137_, _07136_);
  nor _15491_ (_07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15492_ (_07140_, _07139_, _06113_);
  nor _15493_ (_07141_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _15494_ (_07142_, _07141_);
  and _15495_ (_07143_, _07142_, _07140_);
  not _15496_ (_07144_, _07143_);
  or _15497_ (_07145_, _06674_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15498_ (_07146_, _06408_, _07114_);
  and _15499_ (_07147_, _07146_, _07145_);
  or _15500_ (_07148_, _07147_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15501_ (_07149_, _07116_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _15502_ (_07150_, _07149_, _07148_);
  or _15503_ (_07151_, _07150_, _07144_);
  nor _15504_ (_07152_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _15505_ (_07153_, _07152_);
  nand _15506_ (_07154_, _07139_, _06276_);
  and _15507_ (_07155_, _07154_, _07153_);
  not _15508_ (_07156_, _07155_);
  and _15509_ (_07157_, _06666_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15510_ (_07158_, _07157_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15511_ (_07159_, _07123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _15512_ (_07160_, _07159_, _07158_);
  or _15513_ (_07161_, _07160_, _07156_);
  nand _15514_ (_07162_, _07149_, _07148_);
  or _15515_ (_07163_, _07162_, _07143_);
  and _15516_ (_07164_, _07163_, _07151_);
  not _15517_ (_07165_, _07164_);
  or _15518_ (_07166_, _07165_, _07161_);
  and _15519_ (_07167_, _07166_, _07151_);
  nand _15520_ (_07168_, _07159_, _07158_);
  or _15521_ (_07169_, _07168_, _07155_);
  and _15522_ (_07170_, _07169_, _07161_);
  and _15523_ (_07171_, _07170_, _07164_);
  not _15524_ (_07172_, _07139_);
  or _15525_ (_07173_, _07172_, _06297_);
  nor _15526_ (_07174_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _15527_ (_07175_, _07174_);
  nand _15528_ (_07176_, _07175_, _07173_);
  and _15529_ (_07177_, _06674_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15530_ (_07178_, _07177_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15531_ (_07179_, _07127_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _15532_ (_07180_, _07179_, _07178_);
  or _15533_ (_07181_, _07180_, _07176_);
  nor _15534_ (_07182_, _07135_, _07112_);
  nor _15535_ (_07183_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _15536_ (_07184_, _07183_);
  nand _15537_ (_07185_, _07139_, _06166_);
  and _15538_ (_07186_, _07185_, _07184_);
  not _15539_ (_07187_, _07186_);
  or _15540_ (_07188_, _07187_, _07182_);
  and _15541_ (_07189_, _07175_, _07173_);
  nand _15542_ (_07190_, _07179_, _07178_);
  or _15543_ (_07191_, _07190_, _07189_);
  nand _15544_ (_07192_, _07191_, _07181_);
  or _15545_ (_07193_, _07192_, _07188_);
  nand _15546_ (_07194_, _07193_, _07181_);
  nand _15547_ (_07195_, _07194_, _07171_);
  and _15548_ (_07196_, _07195_, _07167_);
  and _15549_ (_07197_, _07147_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15550_ (_07198_, _07197_);
  nor _15551_ (_07199_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _15552_ (_07200_, _07199_);
  nand _15553_ (_07201_, _07139_, _06187_);
  and _15554_ (_07202_, _07201_, _07200_);
  nand _15555_ (_07203_, _07202_, _07198_);
  or _15556_ (_07204_, _07202_, _07198_);
  nand _15557_ (_07205_, _07204_, _07203_);
  nand _15558_ (_07206_, _07157_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15559_ (_07207_, _07172_, _06251_);
  nor _15560_ (_07208_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _15561_ (_07209_, _07208_);
  and _15562_ (_07210_, _07209_, _07207_);
  nand _15563_ (_07211_, _07210_, _07206_);
  and _15564_ (_07212_, _07177_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15565_ (_07213_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _15566_ (_07214_, _07213_);
  or _15567_ (_07215_, _07172_, _06230_);
  nand _15568_ (_07216_, _07215_, _07214_);
  and _15569_ (_07217_, _07216_, _07212_);
  or _15570_ (_07218_, _07210_, _07206_);
  nand _15571_ (_07219_, _07218_, _07211_);
  or _15572_ (_07220_, _07219_, _07217_);
  and _15573_ (_07221_, _07220_, _07211_);
  or _15574_ (_07222_, _07221_, _07205_);
  nand _15575_ (_07223_, _07222_, _07203_);
  not _15576_ (_07224_, _07182_);
  or _15577_ (_07225_, _07186_, _07224_);
  and _15578_ (_07226_, _07225_, _07188_);
  and _15579_ (_07227_, _07191_, _07181_);
  and _15580_ (_07228_, _07227_, _07226_);
  and _15581_ (_07229_, _07228_, _07171_);
  nand _15582_ (_07230_, _07229_, _07223_);
  nand _15583_ (_07231_, _07230_, _07196_);
  not _15584_ (_07232_, _07138_);
  and _15585_ (_07233_, _07232_, _07132_);
  nand _15586_ (_07235_, _07233_, _07231_);
  and _15587_ (_07236_, _07235_, _07143_);
  not _15588_ (_07237_, _07236_);
  and _15589_ (_07239_, _07233_, _07231_);
  and _15590_ (_07240_, _07180_, _07176_);
  not _15591_ (_07241_, _07188_);
  and _15592_ (_07242_, _07226_, _07223_);
  nor _15593_ (_07243_, _07242_, _07241_);
  or _15594_ (_07244_, _07243_, _07240_);
  and _15595_ (_07245_, _07244_, _07181_);
  not _15596_ (_07246_, _07245_);
  nand _15597_ (_07247_, _07246_, _07170_);
  and _15598_ (_07248_, _07247_, _07161_);
  nand _15599_ (_07249_, _07248_, _07164_);
  or _15600_ (_07250_, _07248_, _07164_);
  nand _15601_ (_07251_, _07250_, _07249_);
  nand _15602_ (_07252_, _07251_, _07239_);
  and _15603_ (_07253_, _07252_, _07237_);
  or _15604_ (_07254_, _07253_, _07138_);
  or _15605_ (_07255_, _07246_, _07170_);
  nand _15606_ (_07256_, _07255_, _07247_);
  nand _15607_ (_07257_, _07256_, _07239_);
  and _15608_ (_07259_, _07235_, _07156_);
  not _15609_ (_07261_, _07259_);
  and _15610_ (_07262_, _07261_, _07257_);
  nand _15611_ (_07263_, _07262_, _07162_);
  nand _15612_ (_07264_, _07253_, _07138_);
  nand _15613_ (_07265_, _07264_, _07254_);
  or _15614_ (_07266_, _07265_, _07263_);
  and _15615_ (_07267_, _07266_, _07254_);
  and _15616_ (_07268_, _07264_, _07254_);
  or _15617_ (_07269_, _07262_, _07162_);
  and _15618_ (_07270_, _07269_, _07263_);
  and _15619_ (_07271_, _07270_, _07268_);
  nand _15620_ (_07272_, _07192_, _07243_);
  or _15621_ (_07273_, _07192_, _07243_);
  nand _15622_ (_07274_, _07273_, _07272_);
  nand _15623_ (_07275_, _07274_, _07239_);
  and _15624_ (_07276_, _07235_, _07176_);
  not _15625_ (_07277_, _07276_);
  and _15626_ (_07278_, _07277_, _07275_);
  and _15627_ (_07279_, _07278_, _07168_);
  nor _15628_ (_07280_, _07226_, _07223_);
  or _15629_ (_07281_, _07280_, _07242_);
  and _15630_ (_07282_, _07281_, _07239_);
  and _15631_ (_07283_, _07235_, _07187_);
  nor _15632_ (_07284_, _07283_, _07282_);
  and _15633_ (_07285_, _07284_, _07190_);
  nor _15634_ (_07286_, _07278_, _07168_);
  or _15635_ (_07287_, _07286_, _07279_);
  not _15636_ (_07288_, _07287_);
  and _15637_ (_07289_, _07288_, _07285_);
  nor _15638_ (_07290_, _07289_, _07279_);
  and _15639_ (_07291_, _07221_, _07205_);
  not _15640_ (_07292_, _07291_);
  and _15641_ (_07293_, _07292_, _07222_);
  or _15642_ (_07294_, _07293_, _07235_);
  or _15643_ (_07295_, _07239_, _07202_);
  and _15644_ (_07296_, _07295_, _07294_);
  nor _15645_ (_07297_, _07296_, _07224_);
  not _15646_ (_07298_, _07297_);
  not _15647_ (_07299_, _07212_);
  or _15648_ (_07300_, _07235_, _07299_);
  nand _15649_ (_07301_, _07300_, _07216_);
  or _15650_ (_07302_, _07300_, _07216_);
  and _15651_ (_07303_, _07302_, _07301_);
  nand _15652_ (_07304_, _07303_, _07206_);
  or _15653_ (_07305_, _07303_, _07206_);
  and _15654_ (_07306_, _07305_, _07304_);
  and _15655_ (_07307_, _07139_, _06209_);
  nor _15656_ (_07308_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _15657_ (_07309_, _07308_, _07307_);
  nor _15658_ (_07310_, _07309_, _07299_);
  not _15659_ (_07311_, _07310_);
  nand _15660_ (_07312_, _07311_, _07306_);
  nand _15661_ (_07313_, _07312_, _07304_);
  and _15662_ (_07314_, _07219_, _07217_);
  not _15663_ (_07315_, _07314_);
  and _15664_ (_07316_, _07315_, _07220_);
  or _15665_ (_07317_, _07316_, _07235_);
  or _15666_ (_07318_, _07239_, _07210_);
  and _15667_ (_07319_, _07318_, _07317_);
  nand _15668_ (_07320_, _07319_, _07198_);
  or _15669_ (_07321_, _07319_, _07198_);
  and _15670_ (_07322_, _07321_, _07320_);
  nand _15671_ (_07323_, _07322_, _07313_);
  and _15672_ (_07324_, _07296_, _07224_);
  not _15673_ (_07325_, _07324_);
  and _15674_ (_07326_, _07325_, _07320_);
  nand _15675_ (_07327_, _07326_, _07323_);
  and _15676_ (_07328_, _07327_, _07298_);
  nor _15677_ (_07329_, _07284_, _07190_);
  nor _15678_ (_07330_, _07329_, _07285_);
  and _15679_ (_07331_, _07288_, _07330_);
  nand _15680_ (_07332_, _07331_, _07328_);
  nand _15681_ (_07333_, _07332_, _07290_);
  nand _15682_ (_07334_, _07333_, _07271_);
  nand _15683_ (_07335_, _07334_, _07267_);
  and _15684_ (_07336_, _07335_, _07132_);
  nand _15685_ (_07337_, _07333_, _07270_);
  or _15686_ (_07338_, _07333_, _07270_);
  nand _15687_ (_07339_, _07338_, _07337_);
  nand _15688_ (_07340_, _07339_, _07336_);
  or _15689_ (_07341_, _07336_, _07262_);
  and _15690_ (_07342_, _07341_, _07340_);
  nand _15691_ (_07343_, _07342_, _07108_);
  and _15692_ (_07344_, _06344_, _06124_);
  and _15693_ (_07345_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not _15694_ (_07346_, _07345_);
  or _15695_ (_07347_, _07073_, _07067_);
  nand _15696_ (_07348_, _07347_, _07064_);
  and _15697_ (_07349_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _15698_ (_07350_, _07349_, _07014_);
  and _15699_ (_07351_, _07350_, _07348_);
  nor _15700_ (_07352_, _07096_, _07067_);
  nand _15701_ (_07353_, _07350_, _07352_);
  nor _15702_ (_07354_, _07353_, _07094_);
  or _15703_ (_07355_, _07354_, _07351_);
  and _15704_ (_07356_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  not _15705_ (_07357_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _15706_ (_07358_, _06853_, _07357_);
  and _15707_ (_07360_, _07358_, _07356_);
  and _15708_ (_07361_, _07360_, _07355_);
  and _15709_ (_07362_, _07361_, _07346_);
  nand _15710_ (_07363_, _07360_, _07355_);
  and _15711_ (_07364_, _07363_, _07345_);
  or _15712_ (_07365_, _07364_, _07362_);
  nand _15713_ (_07366_, _07365_, _07344_);
  nor _15714_ (_07367_, _06708_, _06642_);
  nor _15715_ (_07368_, _07367_, _06709_);
  nor _15716_ (_07369_, _07368_, _06616_);
  not _15717_ (_07370_, _07369_);
  nor _15718_ (_07371_, _06743_, _06737_);
  nor _15719_ (_07372_, _07371_, _06716_);
  and _15720_ (_07373_, _07372_, _06745_);
  not _15721_ (_07374_, _06756_);
  nor _15722_ (_07375_, _06623_, _06120_);
  nor _15723_ (_07376_, _07375_, _06128_);
  and _15724_ (_07377_, _07376_, _07374_);
  and _15725_ (_07378_, _06311_, _06120_);
  nor _15726_ (_07379_, _06297_, _06120_);
  and _15727_ (_07380_, _07379_, _06255_);
  nor _15728_ (_07381_, _07380_, _07378_);
  nor _15729_ (_07383_, _07381_, _06276_);
  not _15730_ (_07384_, _07383_);
  and _15731_ (_07385_, _07381_, _06276_);
  nor _15732_ (_07386_, _07385_, _06585_);
  and _15733_ (_07387_, _07386_, _07384_);
  nor _15734_ (_07388_, _07387_, _07377_);
  nor _15735_ (_07389_, _06299_, _06113_);
  not _15736_ (_07390_, _07389_);
  and _15737_ (_07391_, _06767_, _07390_);
  not _15738_ (_07392_, _07391_);
  and _15739_ (_07393_, _06754_, _06297_);
  nor _15740_ (_07394_, _07393_, _06303_);
  nor _15741_ (_07395_, _07394_, _07392_);
  not _15742_ (_07396_, _07395_);
  and _15743_ (_07397_, _07392_, _06760_);
  nor _15744_ (_07398_, _07391_, _06755_);
  and _15745_ (_07399_, _07398_, _06303_);
  nor _15746_ (_07400_, _07399_, _07397_);
  and _15747_ (_07401_, _07400_, _07396_);
  nor _15748_ (_07402_, _07401_, _06759_);
  and _15749_ (_07403_, _06628_, _06324_);
  and _15750_ (_07404_, _06626_, _06332_);
  nor _15751_ (_07405_, _06627_, _06337_);
  and _15752_ (_07406_, _06339_, _06276_);
  or _15753_ (_07407_, _07406_, _07405_);
  or _15754_ (_07409_, _07407_, _07404_);
  nor _15755_ (_07410_, _07409_, _07403_);
  not _15756_ (_07411_, _06350_);
  or _15757_ (_07412_, _07411_, _06113_);
  and _15758_ (_07413_, _06352_, _06297_);
  and _15759_ (_07414_, _06349_, _06303_);
  nor _15760_ (_07415_, _07414_, _07413_);
  and _15761_ (_07416_, _07415_, _07412_);
  and _15762_ (_07417_, _07416_, _07410_);
  not _15763_ (_07418_, _07417_);
  nor _15764_ (_07419_, _07418_, _07402_);
  and _15765_ (_07420_, _07419_, _07388_);
  not _15766_ (_07421_, _07420_);
  nor _15767_ (_07422_, _07421_, _07373_);
  and _15768_ (_07423_, _07422_, _07370_);
  and _15769_ (_07424_, _07423_, _07366_);
  nand _15770_ (_07425_, _07424_, _07343_);
  not _15771_ (_07426_, _07425_);
  nor _15772_ (_07427_, _07426_, _07107_);
  and _15773_ (_07428_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05686_);
  and _15774_ (_07429_, _07428_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15775_ (_07430_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _15776_ (_07431_, _07430_, _07429_);
  or _15777_ (_07432_, _07431_, _07427_);
  not _15778_ (_07433_, _07429_);
  and _15779_ (_07434_, _06623_, _06349_);
  and _15780_ (_07435_, _06777_, _06251_);
  and _15781_ (_07437_, _06646_, _06120_);
  not _15782_ (_07438_, _07437_);
  nor _15783_ (_07439_, _06690_, _06113_);
  and _15784_ (_07440_, _07439_, _06312_);
  and _15785_ (_07441_, _07440_, _06666_);
  and _15786_ (_07442_, _07441_, _06408_);
  and _15787_ (_07443_, _07442_, _06701_);
  or _15788_ (_07444_, _07443_, _06302_);
  and _15789_ (_07445_, _07444_, _07438_);
  and _15790_ (_07446_, _06300_, _06113_);
  and _15791_ (_07447_, _06690_, _06677_);
  and _15792_ (_07448_, _06655_, _06660_);
  and _15793_ (_07449_, _07448_, _07447_);
  and _15794_ (_07450_, _07449_, _07446_);
  nor _15795_ (_07451_, _07450_, _06120_);
  not _15796_ (_07452_, _07451_);
  and _15797_ (_07453_, _06577_, _06120_);
  and _15798_ (_07454_, _06646_, _06577_);
  nor _15799_ (_07455_, _07454_, _06120_);
  nor _15800_ (_07456_, _07455_, _07453_);
  and _15801_ (_07457_, _07456_, _07452_);
  and _15802_ (_07458_, _07457_, _07445_);
  and _15803_ (_07459_, _07458_, _06623_);
  nor _15804_ (_07460_, _07458_, _06623_);
  nor _15805_ (_07461_, _07460_, _07459_);
  and _15806_ (_07462_, _07461_, _06145_);
  and _15807_ (_07463_, _06623_, _06120_);
  nor _15808_ (_07464_, _06276_, _06120_);
  or _15809_ (_07465_, _07464_, _07463_);
  and _15810_ (_07466_, _07465_, _06127_);
  or _15811_ (_07467_, _07466_, _07462_);
  or _15812_ (_07468_, _07467_, _07435_);
  and _15813_ (_07469_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _15814_ (_07470_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15815_ (_07471_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06284_);
  nor _15816_ (_07473_, _07471_, _07470_);
  not _15817_ (_07474_, _07473_);
  nor _15818_ (_07475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15819_ (_07477_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06172_);
  nor _15820_ (_07478_, _07477_, _07475_);
  not _15821_ (_07479_, _07478_);
  nor _15822_ (_07480_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _15823_ (_07481_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06193_);
  nor _15824_ (_07483_, _07481_, _07480_);
  not _15825_ (_07484_, _07483_);
  nor _15826_ (_07486_, _07484_, _06749_);
  nor _15827_ (_07487_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _15828_ (_07488_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06210_);
  nor _15829_ (_07489_, _07488_, _07487_);
  and _15830_ (_07490_, _07489_, _07486_);
  nor _15831_ (_07491_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15832_ (_07492_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06243_);
  nor _15833_ (_07493_, _07492_, _07491_);
  nand _15834_ (_07494_, _07493_, _07490_);
  or _15835_ (_07495_, _07494_, _07479_);
  nor _15836_ (_07496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15837_ (_07497_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06151_);
  nor _15838_ (_07498_, _07497_, _07496_);
  not _15839_ (_07499_, _07498_);
  or _15840_ (_07500_, _07499_, _07495_);
  or _15841_ (_07501_, _07500_, _07474_);
  nor _15842_ (_07502_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _15843_ (_07503_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06261_);
  nor _15844_ (_07504_, _07503_, _07502_);
  not _15845_ (_07505_, _07504_);
  and _15846_ (_07506_, _07505_, _07501_);
  not _15847_ (_07507_, _07506_);
  nor _15848_ (_07508_, _07505_, _07501_);
  nor _15849_ (_07509_, _07508_, _06716_);
  and _15850_ (_07511_, _07509_, _07507_);
  and _15851_ (_07512_, _07090_, _07089_);
  not _15852_ (_07514_, _07512_);
  and _15853_ (_07515_, _07514_, _07091_);
  and _15854_ (_07516_, _07515_, _07344_);
  or _15855_ (_07517_, _07516_, _07511_);
  or _15856_ (_07518_, _07517_, _07469_);
  or _15857_ (_07519_, _07518_, _07468_);
  or _15858_ (_07520_, _07519_, _07434_);
  or _15859_ (_07521_, _07520_, _07433_);
  and _15860_ (_07523_, _07521_, _06071_);
  and _15861_ (_06034_, _07523_, _07432_);
  and _15862_ (_07525_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _15863_ (_07526_, _06804_, _06371_);
  and _15864_ (_07527_, _07526_, _06840_);
  and _15865_ (_07528_, _07527_, _06814_);
  and _15866_ (_07530_, _07528_, _06009_);
  nand _15867_ (_07531_, _07335_, _07132_);
  or _15868_ (_07532_, _07322_, _07313_);
  and _15869_ (_07533_, _07532_, _07323_);
  or _15870_ (_07534_, _07533_, _07531_);
  or _15871_ (_07535_, _07336_, _07319_);
  and _15872_ (_07536_, _07535_, _07534_);
  and _15873_ (_07537_, _07536_, _07108_);
  and _15874_ (_07538_, _07103_, _07344_);
  or _15875_ (_07540_, _06729_, _06727_);
  nor _15876_ (_07541_, _06730_, _06716_);
  and _15877_ (_07542_, _07541_, _07540_);
  and _15878_ (_07543_, _06697_, _06687_);
  or _15879_ (_07544_, _07543_, _06698_);
  and _15880_ (_07545_, _07544_, _06615_);
  and _15881_ (_07546_, _06252_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _15882_ (_07547_, _06752_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _15883_ (_07548_, _07547_, _06230_);
  nor _15884_ (_07549_, _07548_, _06429_);
  or _15885_ (_07550_, _07549_, _07546_);
  and _15886_ (_07551_, _07550_, _06751_);
  nor _15887_ (_07552_, _07411_, _06187_);
  and _15888_ (_07553_, _06349_, _06251_);
  and _15889_ (_07554_, _06352_, _06230_);
  or _15890_ (_07555_, _07554_, _07553_);
  nor _15891_ (_07556_, _07555_, _07552_);
  and _15892_ (_07557_, _07556_, _06428_);
  and _15893_ (_07558_, _07557_, _06424_);
  nand _15894_ (_07559_, _07558_, _06418_);
  or _15895_ (_07560_, _07559_, _07551_);
  or _15896_ (_07561_, _07560_, _07545_);
  or _15897_ (_07562_, _07561_, _07542_);
  or _15898_ (_07563_, _07562_, _07538_);
  or _15899_ (_07564_, _07563_, _07537_);
  and _15900_ (_07565_, _07564_, _07530_);
  or _15901_ (_07566_, _07565_, _07525_);
  or _15902_ (_07567_, _07566_, _07429_);
  or _15903_ (_07569_, _07493_, _07490_);
  and _15904_ (_07570_, _07494_, _06715_);
  and _15905_ (_07571_, _07570_, _07569_);
  nor _15906_ (_07572_, _07441_, _06302_);
  and _15907_ (_07573_, _07447_, _07446_);
  nor _15908_ (_07574_, _07573_, _06120_);
  nor _15909_ (_07575_, _07574_, _07572_);
  nand _15910_ (_07576_, _07575_, _06408_);
  or _15911_ (_07577_, _07575_, _06408_);
  and _15912_ (_07578_, _07577_, _06145_);
  and _15913_ (_07579_, _07578_, _07576_);
  or _15914_ (_07580_, _06919_, _06917_);
  and _15915_ (_07581_, _07580_, _06920_);
  and _15916_ (_07583_, _07581_, _07344_);
  and _15917_ (_07584_, _06777_, _06303_);
  and _15918_ (_07585_, _06251_, _06127_);
  and _15919_ (_07586_, _06408_, _06349_);
  and _15920_ (_07587_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or _15921_ (_07588_, _07587_, _07586_);
  or _15922_ (_07590_, _07588_, _07585_);
  or _15923_ (_07591_, _07590_, _07584_);
  or _15924_ (_07592_, _07591_, _07583_);
  or _15925_ (_07593_, _07592_, _07579_);
  or _15926_ (_07594_, _07593_, _07571_);
  or _15927_ (_07595_, _07594_, _07433_);
  and _15928_ (_07596_, _07595_, _06071_);
  and _15929_ (_06049_, _07596_, _07567_);
  and _15930_ (_07597_, _07330_, _07328_);
  nor _15931_ (_07598_, _07597_, _07285_);
  nand _15932_ (_07599_, _07287_, _07598_);
  or _15933_ (_07600_, _07287_, _07598_);
  nand _15934_ (_07601_, _07600_, _07599_);
  nand _15935_ (_07602_, _07601_, _07336_);
  or _15936_ (_07603_, _07336_, _07278_);
  and _15937_ (_07604_, _07603_, _07602_);
  nand _15938_ (_07605_, _07604_, _07108_);
  nand _15939_ (_07606_, _07356_, _07355_);
  nor _15940_ (_07607_, _07358_, _07606_);
  and _15941_ (_07608_, _07358_, _07606_);
  or _15942_ (_07609_, _07608_, _07607_);
  nand _15943_ (_07610_, _07609_, _07344_);
  nor _15944_ (_07611_, _06707_, _06645_);
  nor _15945_ (_07612_, _07611_, _06708_);
  nor _15946_ (_07613_, _07612_, _06616_);
  not _15947_ (_07614_, _07613_);
  nor _15948_ (_07615_, _06647_, _06596_);
  or _15949_ (_07616_, _07615_, _06739_);
  not _15950_ (_07617_, _07616_);
  nor _15951_ (_07618_, _07617_, _06736_);
  or _15952_ (_07619_, _07618_, _06716_);
  nor _15953_ (_07621_, _07619_, _06737_);
  nor _15954_ (_07622_, _07393_, _06755_);
  nor _15955_ (_07623_, _07622_, _07392_);
  and _15956_ (_07624_, _07622_, _07392_);
  or _15957_ (_07625_, _07624_, _06759_);
  nor _15958_ (_07626_, _07625_, _07623_);
  and _15959_ (_07627_, _06349_, _06297_);
  not _15960_ (_07628_, _07627_);
  nor _15961_ (_07630_, _06353_, _06166_);
  nor _15962_ (_07631_, _07411_, _06276_);
  nor _15963_ (_07632_, _07631_, _07630_);
  and _15964_ (_07633_, _07632_, _07628_);
  and _15965_ (_07634_, _07633_, _06607_);
  not _15966_ (_07635_, _07634_);
  nor _15967_ (_07636_, _07635_, _07626_);
  and _15968_ (_07637_, _07636_, _06590_);
  not _15969_ (_07638_, _07637_);
  nor _15970_ (_07639_, _07638_, _07621_);
  and _15971_ (_07641_, _07639_, _07614_);
  and _15972_ (_07642_, _07641_, _07610_);
  and _15973_ (_07643_, _07642_, _07605_);
  nor _15974_ (_07644_, _07643_, _07107_);
  and _15975_ (_07645_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _15976_ (_07646_, _07645_, _07429_);
  or _15977_ (_07647_, _07646_, _07644_);
  and _15978_ (_07648_, _06593_, _06349_);
  and _15979_ (_07650_, _06777_, _06230_);
  and _15980_ (_07651_, _07450_, _06646_);
  nor _15981_ (_07652_, _07651_, _06120_);
  not _15982_ (_07653_, _07652_);
  and _15983_ (_07654_, _07653_, _07445_);
  and _15984_ (_07655_, _07654_, _06577_);
  nor _15985_ (_07656_, _07654_, _06577_);
  nor _15986_ (_07657_, _07656_, _07655_);
  nor _15987_ (_07658_, _07657_, _06585_);
  not _15988_ (_07659_, _07379_);
  nor _15989_ (_07660_, _07453_, _06128_);
  and _15990_ (_07661_, _07660_, _07659_);
  or _15991_ (_07662_, _07661_, _07658_);
  or _15992_ (_07663_, _07662_, _07650_);
  and _15993_ (_07664_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  and _15994_ (_07665_, _07500_, _07474_);
  not _15995_ (_07666_, _07665_);
  and _15996_ (_07667_, _07501_, _06715_);
  and _15997_ (_07668_, _07667_, _07666_);
  and _15998_ (_07669_, _06956_, _07344_);
  or _15999_ (_07670_, _07669_, _07668_);
  or _16000_ (_07671_, _07670_, _07664_);
  or _16001_ (_07672_, _07671_, _07663_);
  nor _16002_ (_07673_, _07672_, _07648_);
  nand _16003_ (_07674_, _07673_, _07429_);
  and _16004_ (_07675_, _07674_, _06071_);
  and _16005_ (_06052_, _07675_, _07647_);
  and _16006_ (_06060_, _07609_, _06071_);
  nor _16007_ (_07676_, _07330_, _07328_);
  or _16008_ (_07677_, _07676_, _07597_);
  nand _16009_ (_07678_, _07677_, _07336_);
  or _16010_ (_07679_, _07336_, _07284_);
  and _16011_ (_07680_, _07679_, _07678_);
  nand _16012_ (_07681_, _07680_, _07108_);
  or _16013_ (_07682_, _07356_, _07355_);
  and _16014_ (_07683_, _07682_, _07606_);
  nand _16015_ (_07684_, _07683_, _07344_);
  nor _16016_ (_07685_, _06706_, _06649_);
  and _16017_ (_07686_, _06706_, _06649_);
  nor _16018_ (_07687_, _07686_, _07685_);
  and _16019_ (_07688_, _07687_, _06615_);
  not _16020_ (_07689_, _07688_);
  nor _16021_ (_07690_, _06735_, _06649_);
  not _16022_ (_07691_, _07690_);
  nor _16023_ (_07692_, _06736_, _06716_);
  and _16024_ (_07693_, _07692_, _07691_);
  and _16025_ (_07694_, _06753_, _06166_);
  not _16026_ (_07695_, _07694_);
  nor _16027_ (_07696_, _06752_, _06759_);
  and _16028_ (_07697_, _07696_, _06304_);
  not _16029_ (_07698_, _07697_);
  nor _16030_ (_07699_, _06353_, _06187_);
  not _16031_ (_07700_, _07699_);
  nand _16032_ (_07701_, _06350_, _06297_);
  not _16033_ (_07702_, _07701_);
  and _16034_ (_07703_, _06349_, _06304_);
  nor _16035_ (_07704_, _07703_, _07702_);
  and _16036_ (_07705_, _07704_, _07700_);
  and _16037_ (_07706_, _07705_, _07698_);
  and _16038_ (_07707_, _07706_, _07695_);
  and _16039_ (_07709_, _07707_, _06991_);
  and _16040_ (_07710_, _07709_, _06980_);
  not _16041_ (_07711_, _07710_);
  nor _16042_ (_07712_, _07711_, _07693_);
  and _16043_ (_07713_, _07712_, _07689_);
  and _16044_ (_07714_, _07713_, _07684_);
  and _16045_ (_07715_, _07714_, _07681_);
  nor _16046_ (_07716_, _07715_, _07107_);
  and _16047_ (_07717_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _16048_ (_07718_, _07717_, _07429_);
  or _16049_ (_07719_, _07718_, _07716_);
  and _16050_ (_07720_, _06634_, _06349_);
  and _16051_ (_07721_, _06777_, _06306_);
  and _16052_ (_07722_, _07452_, _07444_);
  nor _16053_ (_07723_, _07722_, _06634_);
  and _16054_ (_07724_, _07722_, _06634_);
  or _16055_ (_07725_, _07724_, _06585_);
  nor _16056_ (_07726_, _07725_, _07723_);
  and _16057_ (_07727_, _06166_, _06302_);
  not _16058_ (_07728_, _07727_);
  nor _16059_ (_07729_, _07437_, _06128_);
  and _16060_ (_07730_, _07729_, _07728_);
  or _16061_ (_07731_, _07730_, _07726_);
  or _16062_ (_07732_, _07731_, _07721_);
  and _16063_ (_07733_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and _16064_ (_07734_, _07499_, _07495_);
  not _16065_ (_07735_, _07734_);
  and _16066_ (_07737_, _07500_, _06715_);
  and _16067_ (_07738_, _07737_, _07735_);
  and _16068_ (_07739_, _06926_, _06924_);
  not _16069_ (_07740_, _07739_);
  and _16070_ (_07741_, _07740_, _06927_);
  and _16071_ (_07742_, _07741_, _07344_);
  or _16072_ (_07743_, _07742_, _07738_);
  or _16073_ (_07744_, _07743_, _07733_);
  or _16074_ (_07745_, _07744_, _07732_);
  nor _16075_ (_07746_, _07745_, _07720_);
  nand _16076_ (_07747_, _07746_, _07429_);
  and _16077_ (_07748_, _07747_, _06071_);
  and _16078_ (_06063_, _07748_, _07719_);
  and _16079_ (_06074_, _07683_, _06071_);
  not _16080_ (_07749_, _07349_);
  and _16081_ (_07750_, _07749_, _07101_);
  or _16082_ (_07751_, _07750_, _07355_);
  nor _16083_ (_06092_, _07751_, rst);
  not _16084_ (_07752_, _05993_);
  and _16085_ (_07753_, _06004_, _05981_);
  and _16086_ (_07754_, _07753_, _07752_);
  and _16087_ (_07755_, _07104_, _07754_);
  and _16088_ (_07756_, _07755_, _06840_);
  nor _16089_ (_07757_, _07756_, _07429_);
  or _16090_ (_07758_, _07757_, _07564_);
  not _16091_ (_07759_, _07757_);
  or _16092_ (_07760_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _16093_ (_07761_, _07760_, _06071_);
  and _16094_ (_06096_, _07761_, _07758_);
  nand _16095_ (_07762_, _07759_, _07643_);
  or _16096_ (_07763_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _16097_ (_07764_, _07763_, _06071_);
  and _16098_ (_06130_, _07764_, _07762_);
  not _16099_ (_07765_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _16100_ (_07766_, _07428_, _07765_);
  not _16101_ (_07767_, _05937_);
  and _16102_ (_07768_, _07767_, _05923_);
  and _16103_ (_07769_, _07768_, _05968_);
  and _16104_ (_07770_, _07769_, _06372_);
  and _16105_ (_07771_, _07770_, _06012_);
  nor _16106_ (_07772_, _07771_, _07766_);
  not _16107_ (_07773_, _07772_);
  or _16108_ (_07774_, _07336_, _07253_);
  and _16109_ (_07775_, _07337_, _07263_);
  nand _16110_ (_07776_, _07775_, _07268_);
  or _16111_ (_07777_, _07775_, _07268_);
  nand _16112_ (_07778_, _07777_, _07776_);
  nand _16113_ (_07779_, _07778_, _07336_);
  nand _16114_ (_07781_, _07779_, _07774_);
  nand _16115_ (_07782_, _07781_, _07108_);
  and _16116_ (_07783_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or _16117_ (_07784_, _07363_, _07346_);
  nand _16118_ (_07785_, _07784_, _07783_);
  or _16119_ (_07786_, _07784_, _07783_);
  nand _16120_ (_07787_, _07786_, _07785_);
  nand _16121_ (_07788_, _07787_, _07344_);
  not _16122_ (_07789_, _06327_);
  and _16123_ (_07790_, _06710_, _07789_);
  nor _16124_ (_07791_, _06710_, _07789_);
  nor _16125_ (_07792_, _07791_, _07790_);
  and _16126_ (_07793_, _07792_, _06615_);
  not _16127_ (_07794_, _07793_);
  nor _16128_ (_07795_, _06747_, _07789_);
  and _16129_ (_07796_, _06747_, _07789_);
  or _16130_ (_07797_, _07796_, _07795_);
  nor _16131_ (_07798_, _07797_, _06716_);
  nor _16132_ (_07799_, _07391_, _06760_);
  nor _16133_ (_07800_, _07799_, _06113_);
  and _16134_ (_07801_, _07799_, _06113_);
  nor _16135_ (_07802_, _07801_, _07800_);
  nor _16136_ (_07803_, _07802_, _06759_);
  nor _16137_ (_07804_, _06353_, _06276_);
  and _16138_ (_07805_, _06787_, _06302_);
  nor _16139_ (_07806_, _07805_, _07804_);
  and _16140_ (_07807_, _06349_, _06776_);
  and _16141_ (_07808_, _06789_, _06306_);
  nor _16142_ (_07809_, _07808_, _07807_);
  and _16143_ (_07810_, _07809_, _07806_);
  and _16144_ (_07811_, _07810_, _06343_);
  not _16145_ (_07812_, _07811_);
  nor _16146_ (_07813_, _07812_, _07803_);
  and _16147_ (_07814_, _07813_, _06319_);
  not _16148_ (_07815_, _07814_);
  nor _16149_ (_07816_, _07815_, _07798_);
  and _16150_ (_07817_, _07816_, _07794_);
  and _16151_ (_07818_, _07817_, _07788_);
  nand _16152_ (_07819_, _07818_, _07782_);
  nand _16153_ (_07820_, _07819_, _07773_);
  not _16154_ (_07821_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _16155_ (_07822_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05686_);
  and _16156_ (_07823_, _07822_, _07821_);
  nor _16157_ (_07824_, _05954_, _05937_);
  and _16158_ (_07825_, _07824_, _06833_);
  and _16159_ (_07826_, _07825_, _06815_);
  and _16160_ (_07827_, _07826_, _06805_);
  and _16161_ (_07828_, _07827_, _06803_);
  nor _16162_ (_07829_, _07827_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _16163_ (_07830_, _07823_);
  and _16164_ (_07831_, _07830_, _07772_);
  not _16165_ (_07832_, _07831_);
  nor _16166_ (_07833_, _07832_, _07829_);
  not _16167_ (_07834_, _07833_);
  nor _16168_ (_07835_, _07834_, _07828_);
  nor _16169_ (_07836_, _07835_, _07823_);
  nand _16170_ (_07837_, _07836_, _07820_);
  nor _16171_ (_07838_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _16172_ (_07839_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06086_);
  nor _16173_ (_07840_, _07839_, _07838_);
  and _16174_ (_07841_, _07840_, _07508_);
  nor _16175_ (_07843_, _07840_, _07508_);
  or _16176_ (_07844_, _07843_, _06716_);
  or _16177_ (_07845_, _07844_, _07841_);
  and _16178_ (_07846_, _07092_, _07083_);
  not _16179_ (_07847_, _07846_);
  and _16180_ (_07848_, _07847_, _07093_);
  and _16181_ (_07849_, _07848_, _07344_);
  nor _16182_ (_07850_, _07463_, _07375_);
  not _16183_ (_07851_, _07850_);
  and _16184_ (_07852_, _07851_, _07458_);
  nor _16185_ (_07853_, _07852_, _06139_);
  and _16186_ (_07854_, _07852_, _06139_);
  nor _16187_ (_07855_, _07854_, _07853_);
  and _16188_ (_07856_, _07855_, _06145_);
  and _16189_ (_07857_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and _16190_ (_07858_, _06127_, _06120_);
  or _16191_ (_07859_, _07858_, _06349_);
  and _16192_ (_07860_, _07859_, _06139_);
  or _16193_ (_07861_, _07860_, _07857_);
  and _16194_ (_07862_, _06777_, _06305_);
  and _16195_ (_07863_, _06761_, _06127_);
  or _16196_ (_07864_, _07863_, _07862_);
  nor _16197_ (_07865_, _07864_, _07861_);
  not _16198_ (_07866_, _07865_);
  nor _16199_ (_07867_, _07866_, _07856_);
  not _16200_ (_07868_, _07867_);
  nor _16201_ (_07869_, _07868_, _07849_);
  nand _16202_ (_07870_, _07869_, _07845_);
  or _16203_ (_07871_, _07870_, _07830_);
  and _16204_ (_07872_, _07871_, _07837_);
  and _16205_ (_06199_, _07872_, _06071_);
  and _16206_ (_07873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _16207_ (_07874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _16208_ (_07875_, _07874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _16209_ (_07876_, _07875_);
  nor _16210_ (_07877_, _07876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not _16211_ (_07878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _16212_ (_07879_, _07878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _16213_ (_07880_, _07879_, _07877_);
  nor _16214_ (_07881_, _07880_, _07873_);
  or _16215_ (_07882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _16216_ (_07883_, _07882_, _06071_);
  nor _16217_ (_06346_, _07883_, _07881_);
  and _16218_ (_07884_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _16219_ (_07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _16220_ (_07886_, _07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _16221_ (_07887_, _07886_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _16222_ (_07888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _16223_ (_07889_, _07885_, _07888_);
  and _16224_ (_07890_, _07889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _16225_ (_07891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _16226_ (_07892_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _07891_);
  not _16227_ (_07893_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _16228_ (_07894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _07893_);
  and _16229_ (_07895_, _07894_, _07892_);
  and _16230_ (_07896_, _07895_, _07890_);
  nor _16231_ (_07897_, _07896_, _07887_);
  not _16232_ (_07898_, _07897_);
  and _16233_ (_07899_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  not _16234_ (_07900_, _07890_);
  nor _16235_ (_07901_, _07895_, _07900_);
  not _16236_ (_07902_, _07885_);
  and _16237_ (_07903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _16238_ (_07904_, _07903_, _07902_);
  not _16239_ (_07905_, _07904_);
  and _16240_ (_07906_, _07888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not _16241_ (_07907_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _16242_ (_07908_, _07885_, _07907_);
  and _16243_ (_07909_, _07908_, _07906_);
  nor _16244_ (_07910_, _07909_, _07890_);
  and _16245_ (_07911_, _07910_, _07905_);
  nor _16246_ (_07912_, _07911_, _07901_);
  not _16247_ (_07913_, _07887_);
  nand _16248_ (_07914_, _07913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _16249_ (_07915_, _07914_, _07912_);
  or _16250_ (_07916_, _07915_, _07899_);
  and _16251_ (_07917_, _07916_, _06560_);
  or _16252_ (_06379_, _07917_, _07884_);
  and _16253_ (_07918_, _06922_, _06920_);
  not _16254_ (_07919_, _07918_);
  and _16255_ (_07920_, _07919_, _06923_);
  and _16256_ (_06589_, _07920_, _06071_);
  and _16257_ (_06604_, _07581_, _06071_);
  and _16258_ (_07922_, _06881_, _06872_);
  nor _16259_ (_07923_, _07922_, _06882_);
  and _16260_ (_06606_, _07923_, _06071_);
  and _16261_ (_07924_, _06885_, _06306_);
  and _16262_ (_06617_, _07924_, _06071_);
  and _16263_ (_07925_, _06701_, _06127_);
  nor _16264_ (_07926_, _06253_, _06120_);
  nor _16265_ (_07927_, _06308_, _06302_);
  nor _16266_ (_07928_, _07927_, _07926_);
  and _16267_ (_07929_, _07928_, _06305_);
  not _16268_ (_07930_, _07929_);
  nor _16269_ (_07931_, _07928_, _06305_);
  nor _16270_ (_07932_, _07931_, _06585_);
  and _16271_ (_07933_, _07932_, _07930_);
  nor _16272_ (_07934_, _07933_, _07925_);
  nor _16273_ (_07935_, _06656_, _06337_);
  and _16274_ (_07936_, _06659_, _06324_);
  nor _16275_ (_07937_, _07936_, _07935_);
  and _16276_ (_07938_, _06657_, _06332_);
  and _16277_ (_07939_, _06339_, _06187_);
  nor _16278_ (_07940_, _07939_, _07938_);
  nor _16279_ (_07941_, _06355_, _06187_);
  not _16280_ (_07942_, _07941_);
  and _16281_ (_07943_, _07942_, _07940_);
  and _16282_ (_07944_, _07943_, _07937_);
  and _16283_ (_07945_, _07944_, _07934_);
  and _16284_ (_07946_, _06374_, _06011_);
  nand _16285_ (_07947_, _07946_, _07945_);
  or _16286_ (_07948_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _16287_ (_07949_, _07948_, _06071_);
  and _16288_ (_06658_, _07949_, _07947_);
  and _16289_ (_07950_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  not _16290_ (_07951_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _16291_ (_07952_, _07897_, _07951_);
  nand _16292_ (_07953_, _07913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor _16293_ (_07954_, _07953_, _07912_);
  or _16294_ (_07955_, _07954_, _07952_);
  and _16295_ (_07956_, _07955_, _06560_);
  or _16296_ (_06679_, _07956_, _07950_);
  not _16297_ (_07957_, _06374_);
  nand _16298_ (_07958_, _06438_, _07957_);
  and _16299_ (_07959_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _16300_ (_07960_, _06691_, _06332_);
  and _16301_ (_07961_, _06339_, _06209_);
  nor _16302_ (_07962_, _07961_, _07960_);
  and _16303_ (_07963_, _06674_, _06127_);
  and _16304_ (_07964_, _06145_, _06209_);
  nor _16305_ (_07965_, _07964_, _07963_);
  nor _16306_ (_07966_, _07808_, _06788_);
  and _16307_ (_07967_, _07966_, _07965_);
  and _16308_ (_07968_, _07967_, _07962_);
  nor _16309_ (_07969_, _06691_, _06770_);
  nor _16310_ (_07970_, _07969_, _06336_);
  or _16311_ (_07971_, _07970_, _06692_);
  nor _16312_ (_07972_, _06352_, _06349_);
  and _16313_ (_07973_, _07972_, _06348_);
  nor _16314_ (_07974_, _07973_, _06209_);
  not _16315_ (_07975_, _07974_);
  and _16316_ (_07976_, _07975_, _07971_);
  and _16317_ (_07977_, _07976_, _07968_);
  not _16318_ (_07978_, _07977_);
  and _16319_ (_07979_, _06377_, _06011_);
  and _16320_ (_07980_, _07979_, _07978_);
  or _16321_ (_07981_, _06384_, _06362_);
  and _16322_ (_07983_, _07981_, _06373_);
  and _16323_ (_07984_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _16324_ (_07985_, _07984_, _07983_);
  or _16325_ (_07986_, _07985_, _07980_);
  or _16326_ (_07988_, _07986_, _07959_);
  and _16327_ (_06778_, _07988_, _06071_);
  and _16328_ (_07989_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _16329_ (_07990_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _16330_ (_07991_, _07901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _16331_ (_07992_, _07904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _16332_ (_07993_, _07992_, _07910_);
  or _16333_ (_07994_, _07993_, _07991_);
  and _16334_ (_07996_, _07994_, _07913_);
  or _16335_ (_07997_, _07996_, _07990_);
  and _16336_ (_07998_, _07997_, _06560_);
  or _16337_ (_06783_, _07998_, _07989_);
  and _16338_ (_07999_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _16339_ (_08000_, _06993_, _06611_);
  or _16340_ (_08001_, _08000_, _07999_);
  and _16341_ (_06811_, _08001_, _06071_);
  and _16342_ (_08002_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _16343_ (_06909_, _08002_, _07884_);
  and _16344_ (_06950_, _05768_, _06071_);
  not _16345_ (_08003_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and _16346_ (_08004_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08003_);
  and _16347_ (_08005_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [1]);
  or _16348_ (_08006_, _08005_, _08004_);
  and _16349_ (_06953_, _08006_, _06071_);
  nor _16350_ (_08007_, _07344_, _06857_);
  and _16351_ (_08008_, _07344_, _06857_);
  or _16352_ (_08009_, _08008_, _08007_);
  and _16353_ (_07052_, _08009_, _06071_);
  and _16354_ (_07066_, _05788_, _06071_);
  and _16355_ (_07069_, _05810_, _06071_);
  and _16356_ (_07072_, _05829_, _06071_);
  and _16357_ (_07074_, _05847_, _06071_);
  and _16358_ (_07077_, _05880_, _06071_);
  and _16359_ (_07080_, _05726_, _06071_);
  and _16360_ (_07082_, _05747_, _06071_);
  nor _16361_ (_08010_, _06609_, _06996_);
  and _16362_ (_08011_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _16363_ (_08012_, _08011_, _06390_);
  or _16364_ (_08013_, _08012_, _08010_);
  or _16365_ (_08014_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _16366_ (_08015_, _08014_, _06071_);
  and _16367_ (_07111_, _08015_, _08013_);
  and _16368_ (_08016_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _16369_ (_08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _16370_ (_08018_, _08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _16371_ (_08019_, _08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _16372_ (_08020_, _08019_, _08018_);
  or _16373_ (_08021_, _08020_, _08016_);
  and _16374_ (_07125_, _08021_, _06071_);
  and _16375_ (_08022_, _08003_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _16376_ (_08023_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _16377_ (_08024_, _08023_, _08022_);
  and _16378_ (_07131_, _08024_, _06071_);
  nand _16379_ (_08025_, _07336_, _07212_);
  and _16380_ (_08026_, _08025_, _07309_);
  nor _16381_ (_08027_, _08025_, _07309_);
  or _16382_ (_08028_, _08027_, _08026_);
  nand _16383_ (_08029_, _08028_, _07108_);
  not _16384_ (_08030_, _07097_);
  and _16385_ (_08031_, _07096_, _07094_);
  nor _16386_ (_08032_, _08031_, _08030_);
  and _16387_ (_08033_, _08032_, _07344_);
  and _16388_ (_08034_, _06350_, _06230_);
  nor _16389_ (_08035_, _06751_, _06349_);
  nor _16390_ (_08036_, _08035_, _06209_);
  nor _16391_ (_08037_, _08036_, _08034_);
  nor _16392_ (_08038_, _06693_, _06302_);
  nor _16393_ (_08039_, _08038_, _06726_);
  nor _16394_ (_08040_, _06715_, _06615_);
  not _16395_ (_08041_, _08040_);
  and _16396_ (_08042_, _08041_, _08039_);
  and _16397_ (_08043_, _06781_, _06776_);
  and _16398_ (_08044_, _06777_, _06302_);
  nor _16399_ (_08045_, _08044_, _08043_);
  and _16400_ (_08046_, _08045_, _07965_);
  nand _16401_ (_08047_, _08046_, _07962_);
  nor _16402_ (_08048_, _08047_, _08042_);
  and _16403_ (_08049_, _08048_, _08037_);
  and _16404_ (_08050_, _08049_, _07971_);
  not _16405_ (_08051_, _08050_);
  nor _16406_ (_08052_, _08051_, _08033_);
  and _16407_ (_08053_, _08052_, _08029_);
  nand _16408_ (_08054_, _08053_, _07759_);
  or _16409_ (_08056_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _16410_ (_08057_, _08056_, _06071_);
  and _16411_ (_07234_, _08057_, _08054_);
  or _16412_ (_08058_, _07311_, _07306_);
  and _16413_ (_08059_, _08058_, _07312_);
  or _16414_ (_08060_, _08059_, _07531_);
  or _16415_ (_08061_, _07336_, _07303_);
  and _16416_ (_08062_, _08061_, _08060_);
  nand _16417_ (_08063_, _08062_, _07108_);
  nand _16418_ (_08064_, _07098_, _07067_);
  and _16419_ (_08065_, _08064_, _07099_);
  nand _16420_ (_08066_, _08065_, _07344_);
  and _16421_ (_08067_, _06695_, _06689_);
  nor _16422_ (_08068_, _08067_, _06696_);
  nor _16423_ (_08069_, _08068_, _06616_);
  not _16424_ (_08070_, _08069_);
  and _16425_ (_08071_, _06666_, _06127_);
  nor _16426_ (_08072_, _06230_, _06209_);
  and _16427_ (_08073_, _06230_, _06209_);
  nor _16428_ (_08074_, _08073_, _08072_);
  nor _16429_ (_08075_, _08074_, _06302_);
  and _16430_ (_08076_, _08074_, _06302_);
  nor _16431_ (_08077_, _08076_, _08075_);
  nor _16432_ (_08078_, _08077_, _06585_);
  nor _16433_ (_08079_, _08078_, _08071_);
  nand _16434_ (_08080_, _06350_, _06251_);
  nor _16435_ (_08081_, _06353_, _06209_);
  and _16436_ (_08082_, _06349_, _06230_);
  nor _16437_ (_08083_, _08082_, _08081_);
  and _16438_ (_08084_, _08083_, _08080_);
  and _16439_ (_08086_, _06669_, _06324_);
  nor _16440_ (_08087_, _06668_, _06337_);
  not _16441_ (_08088_, _08087_);
  and _16442_ (_08090_, _06667_, _06332_);
  nor _16443_ (_08091_, _06426_, _06230_);
  nor _16444_ (_08092_, _08091_, _08090_);
  nand _16445_ (_08093_, _08092_, _08088_);
  nor _16446_ (_08094_, _08093_, _08086_);
  and _16447_ (_08095_, _08094_, _08084_);
  and _16448_ (_08096_, _08095_, _08079_);
  and _16449_ (_08097_, _07547_, _06230_);
  nor _16450_ (_08098_, _08097_, _07548_);
  nor _16451_ (_08099_, _08098_, _06759_);
  nor _16452_ (_08100_, _06691_, _06669_);
  or _16453_ (_08101_, _08100_, _06719_);
  and _16454_ (_08102_, _08101_, _06726_);
  nor _16455_ (_08103_, _08101_, _06726_);
  or _16456_ (_08104_, _08103_, _08102_);
  and _16457_ (_08105_, _08104_, _06715_);
  nor _16458_ (_08106_, _08105_, _08099_);
  and _16459_ (_08107_, _08106_, _08096_);
  and _16460_ (_08108_, _08107_, _08070_);
  and _16461_ (_08109_, _08108_, _08066_);
  and _16462_ (_08110_, _08109_, _08063_);
  nand _16463_ (_08111_, _08110_, _07759_);
  or _16464_ (_08112_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _16465_ (_08113_, _08112_, _06071_);
  and _16466_ (_07238_, _08113_, _08111_);
  nor _16467_ (_08114_, _08053_, _07107_);
  and _16468_ (_08115_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _16469_ (_08116_, _08115_, _07429_);
  or _16470_ (_08117_, _08116_, _08114_);
  and _16471_ (_08118_, _07484_, _06749_);
  nor _16472_ (_08119_, _08118_, _07486_);
  and _16473_ (_08120_, _08119_, _06715_);
  nand _16474_ (_08121_, _07336_, _07108_);
  nor _16475_ (_08122_, _06761_, _06121_);
  not _16476_ (_08123_, _08122_);
  nor _16477_ (_08124_, _08123_, _06314_);
  and _16478_ (_08125_, _08124_, _06674_);
  nor _16479_ (_08126_, _08124_, _06674_);
  nor _16480_ (_08127_, _08126_, _08125_);
  and _16481_ (_08128_, _08127_, _06145_);
  and _16482_ (_08129_, _06674_, _06349_);
  and _16483_ (_08130_, _07924_, _07344_);
  and _16484_ (_08131_, _06777_, _06304_);
  nor _16485_ (_08132_, _06209_, _06128_);
  or _16486_ (_08133_, _08132_, _08131_);
  or _16487_ (_08134_, _08133_, _08130_);
  nor _16488_ (_08135_, _08134_, _08129_);
  not _16489_ (_08136_, _08135_);
  nor _16490_ (_08137_, _08136_, _08128_);
  nand _16491_ (_08138_, _08137_, _08121_);
  or _16492_ (_08139_, _08138_, _08120_);
  or _16493_ (_08140_, _08139_, _07433_);
  and _16494_ (_08141_, _08140_, _06071_);
  and _16495_ (_07258_, _08141_, _08117_);
  nor _16496_ (_08142_, _08110_, _07107_);
  and _16497_ (_08143_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _16498_ (_08144_, _08143_, _07429_);
  or _16499_ (_08145_, _08144_, _08142_);
  and _16500_ (_08146_, _06666_, _06349_);
  and _16501_ (_08147_, _06777_, _06297_);
  nor _16502_ (_08148_, _07440_, _06302_);
  and _16503_ (_08150_, _06690_, _07446_);
  nor _16504_ (_08151_, _08150_, _06120_);
  or _16505_ (_08152_, _08151_, _08148_);
  nor _16506_ (_08153_, _08152_, _06666_);
  and _16507_ (_08154_, _08152_, _06666_);
  nor _16508_ (_08155_, _08154_, _08153_);
  nor _16509_ (_08156_, _08155_, _06585_);
  and _16510_ (_08158_, _06230_, _06127_);
  or _16511_ (_08159_, _08158_, _08156_);
  or _16512_ (_08160_, _08159_, _08147_);
  and _16513_ (_08161_, _07239_, _07108_);
  nor _16514_ (_08162_, _07489_, _07486_);
  nor _16515_ (_08163_, _08162_, _07490_);
  and _16516_ (_08164_, _08163_, _06715_);
  and _16517_ (_08165_, _07923_, _07344_);
  or _16518_ (_08166_, _08165_, _08164_);
  or _16519_ (_08167_, _08166_, _08161_);
  or _16520_ (_08168_, _08167_, _08160_);
  nor _16521_ (_08169_, _08168_, _08146_);
  nand _16522_ (_08170_, _08169_, _07429_);
  and _16523_ (_08171_, _08170_, _06071_);
  and _16524_ (_07260_, _08171_, _08145_);
  nor _16525_ (_08172_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _16526_ (_08173_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor _16527_ (_08174_, _08173_, _08172_);
  not _16528_ (_08175_, _08174_);
  not _16529_ (_08176_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _16530_ (_08177_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _16531_ (_08178_, _06530_, _08177_);
  nor _16532_ (_08179_, _08178_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _16533_ (_08180_, _08178_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16534_ (_08181_, _08180_, _08179_);
  nor _16535_ (_08182_, _08181_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16536_ (_08183_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor _16537_ (_08184_, _08183_, _08182_);
  nor _16538_ (_08185_, _08184_, _08176_);
  and _16539_ (_08186_, _08184_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _16540_ (_08187_, _08186_, _08185_);
  nor _16541_ (_08188_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _16542_ (_08189_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor _16543_ (_08190_, _08189_, _08188_);
  and _16544_ (_08191_, _06530_, _08177_);
  nor _16545_ (_08192_, _08191_, _08178_);
  nor _16546_ (_08193_, _08192_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16547_ (_08194_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor _16548_ (_08195_, _08194_, _08193_);
  nor _16549_ (_08196_, _08195_, _08190_);
  not _16550_ (_08197_, _08196_);
  nor _16551_ (_08198_, _08197_, _08187_);
  or _16552_ (_08199_, _08198_, _08175_);
  and _16553_ (_08200_, _08195_, _08190_);
  not _16554_ (_08201_, _08200_);
  nor _16555_ (_08202_, _08184_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _16556_ (_08203_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _16557_ (_08204_, _08184_, _08203_);
  or _16558_ (_08205_, _08204_, _08202_);
  nor _16559_ (_08206_, _08205_, _08201_);
  not _16560_ (_08207_, _08190_);
  nor _16561_ (_08208_, _08195_, _08207_);
  not _16562_ (_08209_, _08208_);
  not _16563_ (_08210_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16564_ (_08211_, _08184_, _08210_);
  and _16565_ (_08212_, _08184_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16566_ (_08213_, _08212_, _08211_);
  nor _16567_ (_08214_, _08213_, _08209_);
  not _16568_ (_08215_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _16569_ (_08217_, _08184_, _08215_);
  nor _16570_ (_08218_, _08184_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16571_ (_08219_, _08218_, _08217_);
  not _16572_ (_08220_, _08219_);
  and _16573_ (_08221_, _08195_, _08207_);
  and _16574_ (_08222_, _08221_, _08220_);
  or _16575_ (_08223_, _08222_, _08214_);
  or _16576_ (_08224_, _08223_, _08206_);
  nor _16577_ (_08225_, _08224_, _08199_);
  nor _16578_ (_08227_, _08184_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not _16579_ (_08228_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16580_ (_08229_, _08184_, _08228_);
  or _16581_ (_08230_, _08229_, _08227_);
  nor _16582_ (_08231_, _08230_, _08201_);
  nor _16583_ (_08232_, _08231_, _08174_);
  not _16584_ (_08233_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16585_ (_08234_, _08184_, _08233_);
  nor _16586_ (_08235_, _08184_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16587_ (_08236_, _08235_, _08234_);
  not _16588_ (_08237_, _08236_);
  nand _16589_ (_08238_, _08237_, _08221_);
  and _16590_ (_08239_, _08184_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _16591_ (_08240_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _16592_ (_08241_, _08184_, _08240_);
  nor _16593_ (_08242_, _08241_, _08239_);
  nor _16594_ (_08243_, _08242_, _08209_);
  nor _16595_ (_08244_, _08184_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _16596_ (_08245_, _08244_);
  not _16597_ (_08246_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16598_ (_08247_, _08184_, _08246_);
  nor _16599_ (_08248_, _08247_, _08197_);
  and _16600_ (_08249_, _08248_, _08245_);
  nor _16601_ (_08250_, _08249_, _08243_);
  and _16602_ (_08251_, _08250_, _08238_);
  and _16603_ (_08252_, _08251_, _08232_);
  nor _16604_ (_08253_, _08252_, _08225_);
  not _16605_ (_08254_, _08253_);
  and _16606_ (_08255_, _08254_, word_in[7]);
  not _16607_ (_08256_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16608_ (_08257_, _08174_, _08256_);
  or _16609_ (_08258_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16610_ (_08259_, _08258_, _08257_);
  and _16611_ (_08260_, _08259_, _08196_);
  or _16612_ (_08261_, _08260_, _08184_);
  not _16613_ (_08262_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16614_ (_08263_, _08174_, _08262_);
  or _16615_ (_08264_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16616_ (_08266_, _08264_, _08263_);
  and _16617_ (_08267_, _08266_, _08221_);
  not _16618_ (_08268_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16619_ (_08269_, _08174_, _08268_);
  or _16620_ (_08270_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16621_ (_08271_, _08270_, _08269_);
  and _16622_ (_08272_, _08271_, _08200_);
  or _16623_ (_08273_, _08272_, _08267_);
  not _16624_ (_08274_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16625_ (_08275_, _08174_, _08274_);
  or _16626_ (_08276_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16627_ (_08277_, _08276_, _08275_);
  and _16628_ (_08278_, _08277_, _08208_);
  or _16629_ (_08279_, _08278_, _08273_);
  or _16630_ (_08280_, _08279_, _08261_);
  not _16631_ (_08281_, _08184_);
  not _16632_ (_08282_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16633_ (_08283_, _08174_, _08282_);
  or _16634_ (_08284_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16635_ (_08285_, _08284_, _08283_);
  and _16636_ (_08286_, _08285_, _08196_);
  or _16637_ (_08287_, _08286_, _08281_);
  not _16638_ (_08288_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16639_ (_08289_, _08174_, _08288_);
  or _16640_ (_08290_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16641_ (_08291_, _08290_, _08289_);
  and _16642_ (_08292_, _08291_, _08221_);
  not _16643_ (_08293_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16644_ (_08294_, _08174_, _08293_);
  or _16645_ (_08295_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16646_ (_08296_, _08295_, _08294_);
  and _16647_ (_08297_, _08296_, _08200_);
  or _16648_ (_08298_, _08297_, _08292_);
  not _16649_ (_08299_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16650_ (_08300_, _08174_, _08299_);
  or _16651_ (_08301_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16652_ (_08302_, _08301_, _08300_);
  and _16653_ (_08303_, _08302_, _08208_);
  or _16654_ (_08304_, _08303_, _08298_);
  or _16655_ (_08305_, _08304_, _08287_);
  and _16656_ (_08306_, _08305_, _08280_);
  and _16657_ (_08307_, _08306_, _08253_);
  or _16658_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08307_, _08255_);
  and _16659_ (_08308_, _08207_, _08174_);
  not _16660_ (_08309_, _08308_);
  and _16661_ (_08310_, _08190_, _08174_);
  and _16662_ (_08311_, _08310_, _08195_);
  nor _16663_ (_08312_, _08310_, _08195_);
  nor _16664_ (_08313_, _08312_, _08311_);
  not _16665_ (_08314_, _08313_);
  nor _16666_ (_08315_, _08314_, _08230_);
  nor _16667_ (_08316_, _08311_, _08281_);
  not _16668_ (_08317_, _08195_);
  nor _16669_ (_08318_, _08317_, _08184_);
  and _16670_ (_08319_, _08310_, _08318_);
  nor _16671_ (_08320_, _08319_, _08316_);
  and _16672_ (_08321_, _08320_, _08314_);
  and _16673_ (_08322_, _08321_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _16674_ (_08323_, _08320_, _08313_);
  and _16675_ (_08324_, _08323_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16676_ (_08325_, _08324_, _08322_);
  nor _16677_ (_08326_, _08325_, _08315_);
  nor _16678_ (_08327_, _08326_, _08309_);
  nor _16679_ (_08328_, _08190_, _08174_);
  not _16680_ (_08329_, _08328_);
  nor _16681_ (_08330_, _08314_, _08219_);
  and _16682_ (_08331_, _08321_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _16683_ (_08332_, _08323_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16684_ (_08333_, _08332_, _08331_);
  nor _16685_ (_08334_, _08333_, _08330_);
  nor _16686_ (_08335_, _08334_, _08329_);
  nor _16687_ (_08336_, _08335_, _08327_);
  not _16688_ (_08337_, _08310_);
  nor _16689_ (_08338_, _08314_, _08236_);
  and _16690_ (_08339_, _08321_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16691_ (_08340_, _08323_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _16692_ (_08341_, _08340_, _08339_);
  nor _16693_ (_08342_, _08341_, _08338_);
  nor _16694_ (_08343_, _08342_, _08337_);
  and _16695_ (_08344_, _08190_, _08175_);
  not _16696_ (_08345_, _08344_);
  and _16697_ (_08346_, _08313_, _08281_);
  and _16698_ (_08347_, _08346_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _16699_ (_08348_, _08323_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16700_ (_08349_, _08321_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _16701_ (_08350_, _08313_, _08184_);
  and _16702_ (_08351_, _08350_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or _16703_ (_08352_, _08351_, _08349_);
  or _16704_ (_08353_, _08352_, _08348_);
  nor _16705_ (_08354_, _08353_, _08347_);
  nor _16706_ (_08355_, _08354_, _08345_);
  nor _16707_ (_08356_, _08355_, _08343_);
  and _16708_ (_08357_, _08356_, _08336_);
  or _16709_ (_08358_, _08328_, _08310_);
  not _16710_ (_08359_, _08358_);
  not _16711_ (_08360_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16712_ (_08361_, _08174_, _08360_);
  or _16713_ (_08362_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16714_ (_08363_, _08362_, _08361_);
  and _16715_ (_08364_, _08363_, _08359_);
  not _16716_ (_08365_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16717_ (_08366_, _08174_, _08365_);
  or _16718_ (_08367_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16719_ (_08368_, _08367_, _08366_);
  and _16720_ (_08369_, _08368_, _08358_);
  or _16721_ (_08370_, _08369_, _08364_);
  and _16722_ (_08371_, _08370_, _08323_);
  not _16723_ (_08372_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16724_ (_08373_, _08174_, _08372_);
  or _16725_ (_08374_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16726_ (_08375_, _08374_, _08373_);
  and _16727_ (_08376_, _08375_, _08359_);
  not _16728_ (_08377_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _16729_ (_08378_, _08174_, _08377_);
  or _16730_ (_08379_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _16731_ (_08380_, _08379_, _08378_);
  and _16732_ (_08381_, _08380_, _08358_);
  or _16733_ (_08382_, _08381_, _08376_);
  and _16734_ (_08383_, _08382_, _08321_);
  not _16735_ (_08384_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16736_ (_08386_, _08174_, _08384_);
  or _16737_ (_08387_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16738_ (_08388_, _08387_, _08386_);
  and _16739_ (_08389_, _08388_, _08359_);
  not _16740_ (_08390_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16741_ (_08391_, _08174_, _08390_);
  or _16742_ (_08392_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16743_ (_08393_, _08392_, _08391_);
  and _16744_ (_08394_, _08393_, _08358_);
  or _16745_ (_08395_, _08394_, _08389_);
  and _16746_ (_08396_, _08395_, _08346_);
  not _16747_ (_08397_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16748_ (_08398_, _08174_, _08397_);
  or _16749_ (_08399_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16750_ (_08400_, _08399_, _08398_);
  and _16751_ (_08401_, _08400_, _08359_);
  not _16752_ (_08402_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16753_ (_08403_, _08174_, _08402_);
  or _16754_ (_08404_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16755_ (_08405_, _08404_, _08403_);
  and _16756_ (_08406_, _08405_, _08358_);
  or _16757_ (_08407_, _08406_, _08401_);
  and _16758_ (_08408_, _08407_, _08350_);
  or _16759_ (_08409_, _08408_, _08396_);
  or _16760_ (_08410_, _08409_, _08383_);
  nor _16761_ (_08411_, _08410_, _08371_);
  nor _16762_ (_08412_, _08411_, _08357_);
  and _16763_ (_08413_, _08357_, word_in[15]);
  or _16764_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08413_, _08412_);
  nor _16765_ (_08414_, _08200_, _08196_);
  not _16766_ (_08415_, _08414_);
  nor _16767_ (_08416_, _08415_, _08205_);
  and _16768_ (_08417_, _08200_, _08184_);
  nor _16769_ (_08418_, _08200_, _08184_);
  nor _16770_ (_08419_, _08418_, _08417_);
  and _16771_ (_08420_, _08415_, _08419_);
  and _16772_ (_08421_, _08420_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16773_ (_08422_, _08414_, _08419_);
  and _16774_ (_08423_, _08422_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _16775_ (_08424_, _08423_, _08421_);
  nor _16776_ (_08425_, _08424_, _08416_);
  nor _16777_ (_08426_, _08425_, _08309_);
  not _16778_ (_08427_, _08426_);
  and _16779_ (_08428_, _08344_, _08318_);
  nand _16780_ (_08429_, _08428_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _16781_ (_08430_, _08415_, _08236_);
  and _16782_ (_08431_, _08422_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16783_ (_08432_, _08431_, _08430_);
  or _16784_ (_08433_, _08432_, _08345_);
  and _16785_ (_08434_, _08433_, _08429_);
  and _16786_ (_08435_, _08434_, _08427_);
  nor _16787_ (_08436_, _08415_, _08230_);
  and _16788_ (_08437_, _08420_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16789_ (_08438_, _08422_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16790_ (_08439_, _08438_, _08437_);
  nor _16791_ (_08440_, _08439_, _08436_);
  nor _16792_ (_08441_, _08440_, _08329_);
  nor _16793_ (_08442_, _08415_, _08219_);
  and _16794_ (_08443_, _08420_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16795_ (_08444_, _08422_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16796_ (_08445_, _08444_, _08443_);
  nor _16797_ (_08446_, _08445_, _08442_);
  nor _16798_ (_08448_, _08446_, _08337_);
  nor _16799_ (_08449_, _08448_, _08441_);
  and _16800_ (_08450_, _08449_, _08435_);
  and _16801_ (_08451_, _08450_, word_in[23]);
  and _16802_ (_08452_, _08266_, _08208_);
  and _16803_ (_08453_, _08277_, _08196_);
  or _16804_ (_08454_, _08453_, _08452_);
  and _16805_ (_08455_, _08271_, _08221_);
  and _16806_ (_08456_, _08259_, _08200_);
  or _16807_ (_08457_, _08456_, _08455_);
  or _16808_ (_08458_, _08457_, _08454_);
  or _16809_ (_08459_, _08458_, _08419_);
  not _16810_ (_08460_, _08419_);
  and _16811_ (_08461_, _08291_, _08208_);
  and _16812_ (_08462_, _08302_, _08196_);
  or _16813_ (_08463_, _08462_, _08461_);
  and _16814_ (_08464_, _08296_, _08221_);
  and _16815_ (_08465_, _08285_, _08200_);
  or _16816_ (_08466_, _08465_, _08464_);
  or _16817_ (_08467_, _08466_, _08463_);
  or _16818_ (_08468_, _08467_, _08460_);
  nand _16819_ (_08469_, _08468_, _08459_);
  nor _16820_ (_08470_, _08469_, _08450_);
  or _16821_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08470_, _08451_);
  nor _16822_ (_08471_, _08329_, _08195_);
  nand _16823_ (_08472_, _08329_, _08195_);
  not _16824_ (_08473_, _08472_);
  nor _16825_ (_08474_, _08473_, _08471_);
  not _16826_ (_08475_, _08474_);
  nor _16827_ (_08476_, _08475_, _08236_);
  nor _16828_ (_08477_, _08472_, _08184_);
  and _16829_ (_08478_, _08472_, _08184_);
  nor _16830_ (_08479_, _08478_, _08477_);
  and _16831_ (_08480_, _08479_, _08475_);
  and _16832_ (_08481_, _08480_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16833_ (_08482_, _08479_, _08474_);
  and _16834_ (_08483_, _08482_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _16835_ (_08484_, _08483_, _08481_);
  nor _16836_ (_08485_, _08484_, _08476_);
  nor _16837_ (_08486_, _08485_, _08309_);
  and _16838_ (_08487_, _08471_, _08211_);
  nor _16839_ (_08488_, _08475_, _08205_);
  and _16840_ (_08489_, _08482_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16841_ (_08490_, _08489_, _08488_);
  and _16842_ (_08491_, _08490_, _08328_);
  nor _16843_ (_08492_, _08491_, _08487_);
  not _16844_ (_08493_, _08492_);
  nor _16845_ (_08494_, _08493_, _08486_);
  nor _16846_ (_08495_, _08475_, _08230_);
  and _16847_ (_08496_, _08480_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _16848_ (_08497_, _08482_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16849_ (_08498_, _08497_, _08496_);
  nor _16850_ (_08499_, _08498_, _08495_);
  nor _16851_ (_08500_, _08499_, _08337_);
  nor _16852_ (_08501_, _08475_, _08219_);
  and _16853_ (_08502_, _08480_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _16854_ (_08503_, _08482_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16855_ (_08504_, _08503_, _08502_);
  nor _16856_ (_08505_, _08504_, _08501_);
  nor _16857_ (_08506_, _08505_, _08345_);
  nor _16858_ (_08507_, _08506_, _08500_);
  and _16859_ (_08508_, _08507_, _08494_);
  and _16860_ (_08509_, _08368_, _08359_);
  and _16861_ (_08510_, _08363_, _08358_);
  or _16862_ (_08511_, _08510_, _08509_);
  and _16863_ (_08512_, _08511_, _08482_);
  and _16864_ (_08513_, _08380_, _08359_);
  and _16865_ (_08514_, _08375_, _08358_);
  or _16866_ (_08515_, _08514_, _08513_);
  and _16867_ (_08516_, _08515_, _08480_);
  and _16868_ (_08517_, _08474_, _08281_);
  and _16869_ (_08518_, _08393_, _08359_);
  and _16870_ (_08519_, _08388_, _08358_);
  or _16871_ (_08520_, _08519_, _08518_);
  and _16872_ (_08521_, _08520_, _08517_);
  and _16873_ (_08522_, _08474_, _08184_);
  and _16874_ (_08523_, _08405_, _08359_);
  and _16875_ (_08524_, _08400_, _08358_);
  or _16876_ (_08525_, _08524_, _08523_);
  and _16877_ (_08526_, _08525_, _08522_);
  or _16878_ (_08527_, _08526_, _08521_);
  or _16879_ (_08528_, _08527_, _08516_);
  nor _16880_ (_08529_, _08528_, _08512_);
  nor _16881_ (_08530_, _08529_, _08508_);
  and _16882_ (_08531_, _08508_, word_in[31]);
  or _16883_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08531_, _08530_);
  and _16884_ (_08532_, _08195_, _08184_);
  nor _16885_ (_08533_, _08417_, _08203_);
  or _16886_ (_08534_, _08533_, _08532_);
  and _16887_ (_07359_, _08534_, _06071_);
  not _16888_ (_08535_, _06526_);
  or _16889_ (_08536_, _08535_, _05810_);
  or _16890_ (_08537_, _06526_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _16891_ (_08538_, _08537_, _06071_);
  and _16892_ (_07382_, _08538_, _08536_);
  and _16893_ (_08539_, _08508_, _06071_);
  and _16894_ (_08540_, _08539_, word_in[31]);
  and _16895_ (_08541_, _08532_, _08328_);
  and _16896_ (_08542_, _08539_, _08541_);
  and _16897_ (_08543_, _08542_, _08540_);
  not _16898_ (_08544_, _08542_);
  and _16899_ (_08545_, _08450_, _06071_);
  and _16900_ (_08546_, _08545_, _08414_);
  and _16901_ (_08547_, _08546_, _08419_);
  and _16902_ (_08548_, _08547_, _08308_);
  not _16903_ (_08549_, _08548_);
  and _16904_ (_08550_, _08357_, _06071_);
  and _16905_ (_08551_, _08550_, _08344_);
  and _16906_ (_08552_, _08551_, _08350_);
  and _16907_ (_08553_, _08225_, _06071_);
  and _16908_ (_08554_, _08553_, _08190_);
  nor _16909_ (_08555_, _08253_, rst);
  and _16910_ (_08556_, _08555_, _08532_);
  and _16911_ (_08557_, _08556_, _08554_);
  and _16912_ (_08558_, _08555_, word_in[7]);
  and _16913_ (_08559_, _08558_, _08557_);
  nor _16914_ (_08560_, _08557_, _08293_);
  nor _16915_ (_08561_, _08560_, _08559_);
  nor _16916_ (_08562_, _08561_, _08552_);
  and _16917_ (_08563_, _08552_, word_in[15]);
  or _16918_ (_08564_, _08563_, _08562_);
  and _16919_ (_08565_, _08564_, _08549_);
  and _16920_ (_08566_, _08545_, word_in[23]);
  and _16921_ (_08567_, _08566_, _08548_);
  or _16922_ (_08568_, _08567_, _08565_);
  and _16923_ (_08569_, _08568_, _08544_);
  or _16924_ (_14025_, _08569_, _08543_);
  or _16925_ (_08570_, _08480_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16926_ (_07408_, _08570_, _06071_);
  or _16927_ (_08571_, _08197_, _08184_);
  nor _16928_ (_08572_, _08417_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand _16929_ (_08573_, _08572_, _08571_);
  and _16930_ (_07436_, _08573_, _06071_);
  and _16931_ (_08574_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _16932_ (_08575_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _16933_ (_08576_, _08575_, _07912_);
  or _16934_ (_08577_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _16935_ (_08578_, _08577_, _06560_);
  and _16936_ (_08579_, _08578_, _08576_);
  or _16937_ (_07472_, _08579_, _08574_);
  and _16938_ (_08580_, _08311_, _08184_);
  not _16939_ (_08581_, _08571_);
  nor _16940_ (_08582_, _08581_, _08580_);
  not _16941_ (_08583_, _08312_);
  or _16942_ (_08584_, _08583_, _08184_);
  nor _16943_ (_08585_, _08584_, _08207_);
  nor _16944_ (_08586_, _08585_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _16945_ (_08587_, _08586_, _08582_);
  and _16946_ (_07476_, _08587_, _06071_);
  and _16947_ (_08588_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _16948_ (_08589_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _16949_ (_08590_, _08589_, _07912_);
  or _16950_ (_08591_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _16951_ (_08592_, _08591_, _06560_);
  and _16952_ (_08593_, _08592_, _08590_);
  or _16953_ (_07482_, _08593_, _08588_);
  or _16954_ (_08594_, _08535_, _05880_);
  or _16955_ (_08595_, _06526_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _16956_ (_08596_, _08595_, _06071_);
  and _16957_ (_07485_, _08596_, _08594_);
  and _16958_ (_08597_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _16959_ (_08598_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _16960_ (_08599_, _08598_, _07912_);
  or _16961_ (_08600_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _16962_ (_08601_, _08600_, _06560_);
  and _16963_ (_08602_, _08601_, _08599_);
  or _16964_ (_07510_, _08602_, _08597_);
  and _16965_ (_08603_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _16966_ (_08604_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _16967_ (_08605_, _08604_, _07912_);
  or _16968_ (_08606_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _16969_ (_08607_, _08606_, _06560_);
  and _16970_ (_08608_, _08607_, _08605_);
  or _16971_ (_07513_, _08608_, _08603_);
  or _16972_ (_08609_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _16973_ (_08611_, _08609_, _07912_);
  or _16974_ (_08612_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _16975_ (_08613_, _08612_, _06560_);
  and _16976_ (_08614_, _08613_, _08611_);
  or _16977_ (_07522_, _08614_, _06559_);
  not _16978_ (_08615_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor _16979_ (_08616_, _08016_, _08615_);
  nor _16980_ (_08617_, _08616_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _16981_ (_08618_, _08616_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _16982_ (_08619_, _08618_, _08617_);
  nor _16983_ (_07524_, _08619_, rst);
  not _16984_ (_08620_, _08321_);
  and _16985_ (_08621_, _08517_, _08310_);
  or _16986_ (_08622_, _08195_, _08184_);
  or _16987_ (_08623_, _08622_, _08344_);
  and _16988_ (_08624_, _08623_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _16989_ (_08625_, _08624_, _08621_);
  and _16990_ (_08626_, _08625_, _08620_);
  and _16991_ (_08627_, _08211_, _08196_);
  or _16992_ (_08628_, _08627_, _08585_);
  or _16993_ (_08629_, _08628_, _08626_);
  and _16994_ (_08630_, _08629_, _08582_);
  or _16995_ (_08631_, _08627_, _08625_);
  and _16996_ (_08632_, _08631_, _08580_);
  or _16997_ (_08633_, _08632_, _08581_);
  or _16998_ (_08634_, _08633_, _08630_);
  and _16999_ (_07529_, _08634_, _06071_);
  or _17000_ (_08635_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17001_ (_08636_, _08635_, _07912_);
  and _17002_ (_08637_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17003_ (_08638_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17004_ (_08639_, _08638_, _06560_);
  or _17005_ (_08640_, _08639_, _08637_);
  and _17006_ (_07539_, _08640_, _08636_);
  or _17007_ (_08641_, _08535_, _05788_);
  or _17008_ (_08642_, _06526_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _17009_ (_08643_, _08642_, _06071_);
  and _17010_ (_07568_, _08643_, _08641_);
  and _17011_ (_08644_, _08328_, _08318_);
  or _17012_ (_08645_, _08644_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17013_ (_08646_, _08645_, _08622_);
  or _17014_ (_08647_, _08646_, _08621_);
  and _17015_ (_08648_, _08647_, _08620_);
  and _17016_ (_08649_, _08645_, _08580_);
  nand _17017_ (_08650_, _08195_, _08174_);
  nand _17018_ (_08651_, _08418_, _08650_);
  nor _17019_ (_08652_, _08651_, _08309_);
  and _17020_ (_08653_, _08471_, _08281_);
  and _17021_ (_08654_, _08653_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _17022_ (_08655_, _08654_, _08652_);
  or _17023_ (_08656_, _08655_, _08649_);
  or _17024_ (_08657_, _08656_, _08585_);
  or _17025_ (_08658_, _08657_, _08648_);
  and _17026_ (_07582_, _08658_, _06071_);
  and _17027_ (_08659_, _08016_, _08615_);
  nor _17028_ (_08660_, _08659_, _08616_);
  and _17029_ (_07589_, _08660_, _06071_);
  or _17030_ (_08661_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17031_ (_08662_, _08661_, _07912_);
  and _17032_ (_08663_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17033_ (_08664_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and _17034_ (_08665_, _08664_, _06560_);
  or _17035_ (_08666_, _08665_, _08663_);
  and _17036_ (_07620_, _08666_, _08662_);
  or _17037_ (_08667_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _17038_ (_08668_, _08667_, _07912_);
  and _17039_ (_08669_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _17040_ (_08670_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and _17041_ (_08671_, _08670_, _06560_);
  or _17042_ (_08672_, _08671_, _08669_);
  and _17043_ (_07629_, _08672_, _08668_);
  not _17044_ (_08673_, _08417_);
  and _17045_ (_08674_, _08584_, _08673_);
  and _17046_ (_08675_, _08201_, _08184_);
  or _17047_ (_08676_, _08675_, _08318_);
  not _17048_ (_08677_, _08418_);
  or _17049_ (_08678_, _08644_, _08621_);
  or _17050_ (_08679_, _08678_, _08677_);
  and _17051_ (_08680_, _08679_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17052_ (_08681_, _08585_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17053_ (_08682_, _08308_, _08318_);
  and _17054_ (_08683_, _08581_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17055_ (_08684_, _08683_, _08682_);
  or _17056_ (_08685_, _08684_, _08681_);
  or _17057_ (_08686_, _08685_, _08680_);
  or _17058_ (_08687_, _08316_, _08477_);
  and _17059_ (_08688_, _08687_, _08686_);
  and _17060_ (_08689_, _08517_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17061_ (_08690_, _08689_, _08644_);
  or _17062_ (_08691_, _08690_, _08688_);
  and _17063_ (_08692_, _08691_, _08676_);
  and _17064_ (_08693_, _08686_, _08580_);
  or _17065_ (_08694_, _08683_, _08621_);
  or _17066_ (_08695_, _08694_, _08681_);
  or _17067_ (_08696_, _08695_, _08693_);
  or _17068_ (_08697_, _08696_, _08692_);
  and _17069_ (_08698_, _08697_, _08674_);
  and _17070_ (_08699_, _08532_, _08344_);
  and _17071_ (_08700_, _08691_, _08699_);
  or _17072_ (_08701_, _08683_, _08585_);
  or _17073_ (_08702_, _08701_, _08693_);
  or _17074_ (_08703_, _08702_, _08700_);
  or _17075_ (_08704_, _08703_, _08698_);
  and _17076_ (_07640_, _08704_, _06071_);
  and _17077_ (_08705_, _06527_, _05689_);
  not _17078_ (_08706_, _08705_);
  or _17079_ (_08707_, _08706_, _05829_);
  not _17080_ (_08708_, _05689_);
  nor _17081_ (_08709_, _06527_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _17082_ (_08710_, _08709_, _08708_);
  nand _17083_ (_08711_, _08710_, _08707_);
  or _17084_ (_08712_, _08706_, _05847_);
  nor _17085_ (_08713_, _06527_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _17086_ (_08714_, _08713_, _08708_);
  nand _17087_ (_08715_, _08714_, _08712_);
  and _17088_ (_08717_, _08715_, _08711_);
  or _17089_ (_08718_, _08706_, _05788_);
  nor _17090_ (_08719_, _06527_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _17091_ (_08720_, _08719_, _08708_);
  nand _17092_ (_08721_, _08720_, _08718_);
  or _17093_ (_08722_, _08706_, _05810_);
  nor _17094_ (_08723_, _06527_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _17095_ (_08724_, _08723_, _08708_);
  and _17096_ (_08725_, _08724_, _08722_);
  not _17097_ (_08726_, _08725_);
  and _17098_ (_08727_, _08726_, _08721_);
  and _17099_ (_08728_, _08727_, _08717_);
  or _17100_ (_08729_, _08706_, _05880_);
  nor _17101_ (_08730_, _06527_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _17102_ (_08731_, _08730_, _08708_);
  and _17103_ (_08732_, _08731_, _08729_);
  or _17104_ (_08733_, _08706_, _05768_);
  nor _17105_ (_08734_, _06527_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _17106_ (_08735_, _08734_, _08708_);
  and _17107_ (_08736_, _08735_, _08733_);
  or _17108_ (_08737_, _08706_, _05747_);
  nor _17109_ (_08739_, _06527_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _17110_ (_08740_, _08739_, _08708_);
  nand _17111_ (_08741_, _08740_, _08737_);
  or _17112_ (_08742_, _08706_, _05726_);
  nor _17113_ (_08744_, _06527_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _17114_ (_08745_, _08744_, _08708_);
  nand _17115_ (_08746_, _08745_, _08742_);
  nor _17116_ (_08748_, _08746_, _08741_);
  and _17117_ (_08749_, _08748_, _08736_);
  and _17118_ (_08750_, _08749_, _08732_);
  nand _17119_ (_08752_, _08750_, _08728_);
  and _17120_ (_08753_, _08720_, _08718_);
  and _17121_ (_08754_, _08725_, _08711_);
  and _17122_ (_08756_, _08754_, _08715_);
  and _17123_ (_08757_, _08756_, _08753_);
  and _17124_ (_08758_, _08746_, _08741_);
  and _17125_ (_08760_, _08758_, _08736_);
  and _17126_ (_08761_, _08760_, _08757_);
  not _17127_ (_08762_, _08761_);
  not _17128_ (_08764_, _08732_);
  and _17129_ (_08765_, _08749_, _08764_);
  and _17130_ (_08767_, _08765_, _08728_);
  and _17131_ (_08768_, _08765_, _08756_);
  nor _17132_ (_08769_, _08768_, _08767_);
  and _17133_ (_08770_, _08769_, _08762_);
  and _17134_ (_08771_, _08770_, _08752_);
  and _17135_ (_08772_, _08732_, _08715_);
  and _17136_ (_08773_, _08772_, _08749_);
  and _17137_ (_08774_, _08773_, _08754_);
  and _17138_ (_08775_, _06527_, _06071_);
  not _17139_ (_08776_, _08775_);
  or _17140_ (_08777_, _08776_, _08768_);
  or _17141_ (_08778_, _08777_, _08774_);
  or _17142_ (_07649_, _08778_, _08771_);
  or _17143_ (_08779_, _08428_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17144_ (_08780_, _08779_, _08651_);
  and _17145_ (_08781_, _08780_, _08677_);
  and _17146_ (_08782_, _08678_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17147_ (_08783_, _08782_, _08682_);
  or _17148_ (_08784_, _08783_, _08781_);
  and _17149_ (_08785_, _08784_, _08687_);
  and _17150_ (_08786_, _08779_, _08580_);
  and _17151_ (_08787_, _08585_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17152_ (_08788_, _08581_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17153_ (_08789_, _08788_, _08621_);
  or _17154_ (_08790_, _08789_, _08787_);
  or _17155_ (_08791_, _08790_, _08644_);
  or _17156_ (_08792_, _08791_, _08786_);
  or _17157_ (_08793_, _08792_, _08785_);
  and _17158_ (_07708_, _08793_, _06071_);
  nand _17159_ (_08794_, _07823_, _07520_);
  or _17160_ (_08795_, _07772_, _07425_);
  nor _17161_ (_08796_, _07826_, _06271_);
  nor _17162_ (_08797_, _08796_, _07773_);
  not _17163_ (_08798_, _08797_);
  not _17164_ (_08799_, _06803_);
  and _17165_ (_08800_, _06004_, _07752_);
  and _17166_ (_08801_, _08800_, _05982_);
  and _17167_ (_08802_, _08801_, _08799_);
  nor _17168_ (_08803_, _08801_, _06271_);
  nor _17169_ (_08804_, _08803_, _08802_);
  and _17170_ (_08805_, _07831_, _07826_);
  not _17171_ (_08806_, _08805_);
  nor _17172_ (_08807_, _08806_, _08804_);
  nor _17173_ (_08808_, _08807_, _08798_);
  nor _17174_ (_08809_, _08808_, _07823_);
  nand _17175_ (_08810_, _08809_, _08795_);
  nand _17176_ (_08811_, _08810_, _08794_);
  and _17177_ (_07736_, _08811_, _06071_);
  not _17178_ (_08812_, _08320_);
  and _17179_ (_08813_, _08653_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17180_ (_08814_, _08517_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17181_ (_08815_, _08814_, _08329_);
  or _17182_ (_08816_, _08815_, _08813_);
  or _17183_ (_08817_, _08428_, _08184_);
  and _17184_ (_08818_, _08817_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _17185_ (_08819_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _17186_ (_08820_, _08190_, _08819_);
  and _17187_ (_08821_, _08820_, _08318_);
  or _17188_ (_08822_, _08821_, _08319_);
  or _17189_ (_08823_, _08822_, _08818_);
  or _17190_ (_08824_, _08823_, _08816_);
  and _17191_ (_08825_, _08824_, _08812_);
  or _17192_ (_08826_, _08821_, _08428_);
  or _17193_ (_08827_, _08826_, _08815_);
  or _17194_ (_08828_, _08827_, _08825_);
  and _17195_ (_08829_, _08828_, _08677_);
  and _17196_ (_08830_, _08824_, _08580_);
  or _17197_ (_08831_, _08813_, _08644_);
  or _17198_ (_08832_, _08831_, _08814_);
  or _17199_ (_08833_, _08832_, _08682_);
  or _17200_ (_08834_, _08833_, _08830_);
  or _17201_ (_08835_, _08834_, _08829_);
  and _17202_ (_07780_, _08835_, _06071_);
  nor _17203_ (_08836_, _08482_, _08281_);
  and _17204_ (_08837_, _08836_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17205_ (_08838_, _08471_, _08184_);
  nor _17206_ (_08839_, _08195_, _08246_);
  or _17207_ (_08840_, _08839_, _08311_);
  and _17208_ (_08841_, _08840_, _08281_);
  and _17209_ (_08842_, _08644_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17210_ (_08843_, _08842_, _08682_);
  or _17211_ (_08844_, _08843_, _08841_);
  or _17212_ (_08845_, _08844_, _08428_);
  or _17213_ (_08847_, _08845_, _08838_);
  or _17214_ (_08848_, _08847_, _08837_);
  and _17215_ (_07842_, _08848_, _06071_);
  and _17216_ (_08849_, _08478_, _08308_);
  nor _17217_ (_08851_, _08675_, _08311_);
  nor _17218_ (_08852_, _08851_, _08849_);
  or _17219_ (_08854_, _08682_, _08653_);
  or _17220_ (_08856_, _08854_, _08852_);
  or _17221_ (_08857_, _08856_, _08699_);
  or _17222_ (_08859_, _08857_, _08517_);
  and _17223_ (_08861_, _08859_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17224_ (_08862_, _08861_, _08420_);
  and _17225_ (_07921_, _08862_, _06071_);
  and _17226_ (_08864_, _06381_, _06011_);
  not _17227_ (_08865_, _08864_);
  and _17228_ (_08867_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _17229_ (_08869_, _08865_, _07945_);
  or _17230_ (_08871_, _08869_, _08867_);
  and _17231_ (_07982_, _08871_, _06071_);
  or _17232_ (_08873_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _17233_ (_08874_, _06530_, _05815_);
  and _17234_ (_08876_, _08874_, _06071_);
  and _17235_ (_07987_, _08876_, _08873_);
  and _17236_ (_08877_, _08532_, _08308_);
  or _17237_ (_08878_, _08877_, _08522_);
  or _17238_ (_08879_, _08878_, _08699_);
  and _17239_ (_08880_, _08316_, _08197_);
  and _17240_ (_08881_, _08428_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17241_ (_08882_, _08678_, _08682_);
  and _17242_ (_08883_, _08882_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17243_ (_08884_, _08883_, _08881_);
  and _17244_ (_08885_, _08849_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _17245_ (_08886_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17246_ (_08887_, _08358_, _08886_);
  and _17247_ (_08888_, _08887_, _08517_);
  and _17248_ (_08889_, _08653_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17249_ (_08891_, _08522_, _08344_);
  and _17250_ (_08892_, _08583_, _08239_);
  or _17251_ (_08893_, _08892_, _08891_);
  or _17252_ (_08895_, _08893_, _08889_);
  or _17253_ (_08896_, _08895_, _08888_);
  or _17254_ (_08897_, _08896_, _08885_);
  or _17255_ (_08898_, _08897_, _08884_);
  and _17256_ (_08899_, _08898_, _08880_);
  or _17257_ (_08900_, _08319_, _08838_);
  and _17258_ (_08901_, _08900_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17259_ (_08902_, _08901_, _08849_);
  or _17260_ (_08903_, _08902_, _08899_);
  and _17261_ (_08904_, _08903_, _08879_);
  or _17262_ (_08905_, _08901_, _08898_);
  and _17263_ (_08906_, _08905_, _08580_);
  and _17264_ (_08907_, _08414_, _08281_);
  and _17265_ (_08908_, _08907_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _17266_ (_08909_, _08571_, _08886_);
  or _17267_ (_08910_, _08909_, _08319_);
  or _17268_ (_08911_, _08910_, _08881_);
  or _17269_ (_08912_, _08911_, _08908_);
  or _17270_ (_08913_, _08912_, _08838_);
  or _17271_ (_08914_, _08913_, _08906_);
  or _17272_ (_08915_, _08914_, _08904_);
  and _17273_ (_07995_, _08915_, _06071_);
  and _17274_ (_08916_, _08532_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17275_ (_08917_, _08208_, _08184_);
  or _17276_ (_08918_, _08174_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17277_ (_08919_, _08918_, _08917_);
  and _17278_ (_08920_, _08208_, _08281_);
  and _17279_ (_08921_, _08920_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17280_ (_08922_, _08921_, _08919_);
  or _17281_ (_08923_, _08922_, _08916_);
  and _17282_ (_08924_, _08212_, _08196_);
  not _17283_ (_08925_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17284_ (_08926_, _08184_, _08925_);
  and _17285_ (_08927_, _08926_, _08209_);
  or _17286_ (_08928_, _08927_, _08924_);
  or _17287_ (_08929_, _08928_, _08923_);
  and _17288_ (_08930_, _08929_, _08350_);
  or _17289_ (_08931_, _08924_, _08891_);
  or _17290_ (_08932_, _08931_, _08930_);
  and _17291_ (_08933_, _08932_, _08197_);
  and _17292_ (_08934_, _08929_, _08580_);
  or _17293_ (_08935_, _08934_, _08838_);
  or _17294_ (_08936_, _08935_, _08849_);
  or _17295_ (_08937_, _08936_, _08926_);
  or _17296_ (_08938_, _08937_, _08933_);
  and _17297_ (_08055_, _08938_, _06071_);
  or _17298_ (_08939_, _07772_, _07643_);
  not _17299_ (_08940_, _07826_);
  and _17300_ (_08941_, _07831_, _08940_);
  and _17301_ (_08942_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _17302_ (_08943_, _08799_, _06032_);
  nor _17303_ (_08944_, _06032_, _06292_);
  nor _17304_ (_08945_, _08944_, _08943_);
  nor _17305_ (_08946_, _08945_, _08806_);
  nor _17306_ (_08947_, _08946_, _08942_);
  and _17307_ (_08948_, _08947_, _07830_);
  nand _17308_ (_08949_, _08948_, _08939_);
  and _17309_ (_08950_, _07823_, _07673_);
  not _17310_ (_08951_, _08950_);
  and _17311_ (_08952_, _08951_, _08949_);
  and _17312_ (_08085_, _08952_, _06071_);
  or _17313_ (_08953_, _08053_, _07772_);
  and _17314_ (_08954_, _07826_, _06383_);
  and _17315_ (_08955_, _08954_, _06803_);
  nor _17316_ (_08956_, _08954_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _17317_ (_08957_, _08956_, _07832_);
  not _17318_ (_08958_, _08957_);
  nor _17319_ (_08959_, _08958_, _08955_);
  nor _17320_ (_08961_, _08959_, _07823_);
  nand _17321_ (_08962_, _08961_, _08953_);
  or _17322_ (_08963_, _08139_, _07830_);
  and _17323_ (_08964_, _08963_, _08962_);
  and _17324_ (_08089_, _08964_, _06071_);
  and _17325_ (_08966_, _08532_, _08329_);
  and _17326_ (_08967_, _08966_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17327_ (_08968_, _08190_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17328_ (_08970_, _08968_, _08517_);
  and _17329_ (_08971_, _08838_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor _17330_ (_08973_, _08571_, _08233_);
  and _17331_ (_08974_, _08318_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17332_ (_08975_, _08974_, _08973_);
  or _17333_ (_08977_, _08975_, _08971_);
  or _17334_ (_08978_, _08977_, _08522_);
  or _17335_ (_08979_, _08978_, _08970_);
  or _17336_ (_08980_, _08979_, _08967_);
  and _17337_ (_08149_, _08980_, _06071_);
  and _17338_ (_08982_, _07104_, _06383_);
  and _17339_ (_08984_, _08982_, _05968_);
  nand _17340_ (_08985_, _08984_, _06365_);
  and _17341_ (_08986_, _08985_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _17342_ (_08987_, _06365_, _05968_);
  and _17343_ (_08988_, _08987_, _08982_);
  not _17344_ (_08989_, _08988_);
  nor _17345_ (_08990_, _08989_, _06993_);
  nor _17346_ (_08991_, _08990_, _08986_);
  nor _17347_ (_08157_, _08991_, rst);
  not _17348_ (_08992_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _17349_ (_08993_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _17350_ (_08994_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08993_);
  not _17351_ (_08995_, _08994_);
  and _17352_ (_08996_, _07902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17353_ (_08997_, _08996_, _08995_);
  and _17354_ (_08998_, _08997_, _07900_);
  nor _17355_ (_08999_, _08998_, _08992_);
  and _17356_ (_09000_, _08998_, rxd_i);
  or _17357_ (_09001_, _09000_, rst);
  or _17358_ (_08216_, _09001_, _08999_);
  not _17359_ (_09002_, rxd_i);
  nor _17360_ (_09003_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _17361_ (_09004_, _09003_, _07892_);
  and _17362_ (_09005_, _07890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17363_ (_09006_, _09005_, _09004_);
  nand _17364_ (_09007_, _09006_, _09002_);
  or _17365_ (_09008_, _09006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _17366_ (_09009_, _09008_, _06071_);
  and _17367_ (_08226_, _09009_, _09007_);
  and _17368_ (_09010_, _08190_, _08184_);
  or _17369_ (_09011_, _08346_, _09010_);
  and _17370_ (_09012_, _09011_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _17371_ (_09013_, _09012_, _08207_);
  and _17372_ (_09014_, _09013_, _08966_);
  or _17373_ (_09015_, _08541_, _08917_);
  nor _17374_ (_09016_, _09010_, _08532_);
  and _17375_ (_09017_, _09016_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _17376_ (_09018_, _09017_, _09015_);
  or _17377_ (_09019_, _09018_, _09014_);
  and _17378_ (_08265_, _09019_, _06071_);
  or _17379_ (_09020_, _08350_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _17380_ (_08385_, _09020_, _06071_);
  or _17381_ (_09021_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not _17382_ (_09022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _17383_ (_09023_, _06530_, _09022_);
  and _17384_ (_09024_, _09023_, _06071_);
  and _17385_ (_08447_, _09024_, _09021_);
  not _17386_ (_09025_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nor _17387_ (_09026_, _05954_, _07767_);
  and _17388_ (_09027_, _09026_, _06809_);
  and _17389_ (_09028_, _09027_, _06815_);
  nand _17390_ (_09029_, _09028_, _06362_);
  nand _17391_ (_09030_, _09029_, _09025_);
  and _17392_ (_09031_, _09030_, _08989_);
  or _17393_ (_09032_, _09029_, _08799_);
  and _17394_ (_09033_, _09032_, _09031_);
  nor _17395_ (_09034_, _06355_, _06856_);
  not _17396_ (_09035_, _09034_);
  and _17397_ (_09036_, _09035_, _08094_);
  and _17398_ (_09037_, _09036_, _08079_);
  nor _17399_ (_09038_, _09037_, _08989_);
  or _17400_ (_09039_, _09038_, _09033_);
  and _17401_ (_08610_, _09039_, _06071_);
  nand _17402_ (_09040_, _07946_, _06434_);
  or _17403_ (_09041_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _17404_ (_09042_, _09041_, _06071_);
  and _17405_ (_08716_, _09042_, _09040_);
  and _17406_ (_09043_, _08539_, word_in[24]);
  and _17407_ (_09044_, _08539_, _08877_);
  and _17408_ (_09045_, _09044_, _09043_);
  and _17409_ (_09046_, _08545_, _08699_);
  not _17410_ (_09047_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _17411_ (_09048_, _08555_, _08190_);
  nor _17412_ (_09049_, _09048_, _08553_);
  and _17413_ (_09050_, _08555_, _08622_);
  not _17414_ (_09051_, _09050_);
  and _17415_ (_09052_, _09051_, _09049_);
  and _17416_ (_09053_, _09052_, _08555_);
  nor _17417_ (_09054_, _09053_, _09047_);
  and _17418_ (_09056_, _08555_, word_in[0]);
  and _17419_ (_09057_, _09056_, _09052_);
  or _17420_ (_09059_, _09057_, _09054_);
  and _17421_ (_09061_, _08550_, _08580_);
  not _17422_ (_09062_, _09061_);
  and _17423_ (_09063_, _09062_, _09059_);
  and _17424_ (_09064_, _09061_, word_in[8]);
  or _17425_ (_09066_, _09064_, _09063_);
  or _17426_ (_09067_, _09066_, _09046_);
  not _17427_ (_09068_, _09044_);
  not _17428_ (_09070_, _09046_);
  or _17429_ (_09071_, _09070_, word_in[16]);
  and _17430_ (_09072_, _09071_, _09068_);
  and _17431_ (_09073_, _09072_, _09067_);
  or _17432_ (_08738_, _09073_, _09045_);
  and _17433_ (_09075_, _08539_, word_in[25]);
  and _17434_ (_09076_, _09075_, _09044_);
  not _17435_ (_09078_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _17436_ (_09079_, _09053_, _09078_);
  and _17437_ (_09080_, _08555_, word_in[1]);
  and _17438_ (_09081_, _09080_, _09052_);
  or _17439_ (_09082_, _09081_, _09079_);
  or _17440_ (_09083_, _09082_, _09061_);
  or _17441_ (_09084_, _09062_, word_in[9]);
  and _17442_ (_09085_, _09084_, _09070_);
  and _17443_ (_09086_, _09085_, _09083_);
  and _17444_ (_09088_, _09046_, word_in[17]);
  or _17445_ (_09089_, _09088_, _09086_);
  and _17446_ (_09090_, _09089_, _09068_);
  or _17447_ (_08743_, _09090_, _09076_);
  or _17448_ (_09091_, _09062_, word_in[10]);
  and _17449_ (_09092_, _09091_, _09070_);
  not _17450_ (_09093_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _17451_ (_09094_, _09053_, _09093_);
  and _17452_ (_09095_, _09053_, word_in[2]);
  or _17453_ (_09096_, _09095_, _09094_);
  or _17454_ (_09097_, _09096_, _09061_);
  and _17455_ (_09098_, _09097_, _09092_);
  and _17456_ (_09099_, _09046_, word_in[18]);
  or _17457_ (_09100_, _09099_, _09044_);
  or _17458_ (_09101_, _09100_, _09098_);
  or _17459_ (_09102_, _09068_, word_in[26]);
  and _17460_ (_08747_, _09102_, _09101_);
  and _17461_ (_09103_, _08539_, word_in[27]);
  and _17462_ (_09104_, _09103_, _09044_);
  not _17463_ (_09105_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _17464_ (_09106_, _09053_, _09105_);
  and _17465_ (_09107_, _09053_, word_in[3]);
  or _17466_ (_09108_, _09107_, _09106_);
  and _17467_ (_09109_, _09108_, _09062_);
  and _17468_ (_09110_, _09061_, word_in[11]);
  or _17469_ (_09111_, _09110_, _09109_);
  and _17470_ (_09112_, _09111_, _09070_);
  and _17471_ (_09113_, _08545_, word_in[19]);
  and _17472_ (_09114_, _09113_, _08699_);
  or _17473_ (_09115_, _09114_, _09112_);
  and _17474_ (_09116_, _09115_, _09068_);
  or _17475_ (_08751_, _09116_, _09104_);
  or _17476_ (_09117_, _09062_, word_in[12]);
  and _17477_ (_09118_, _09117_, _09070_);
  and _17478_ (_09119_, _09053_, word_in[4]);
  not _17479_ (_09120_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _17480_ (_09121_, _09053_, _09120_);
  or _17481_ (_09122_, _09121_, _09119_);
  or _17482_ (_09123_, _09122_, _09061_);
  and _17483_ (_09124_, _09123_, _09118_);
  and _17484_ (_09125_, _09046_, word_in[20]);
  or _17485_ (_09126_, _09125_, _09044_);
  or _17486_ (_09127_, _09126_, _09124_);
  or _17487_ (_09128_, _09068_, word_in[28]);
  and _17488_ (_08755_, _09128_, _09127_);
  or _17489_ (_09129_, _09062_, word_in[13]);
  and _17490_ (_09130_, _09129_, _09070_);
  not _17491_ (_09131_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _17492_ (_09132_, _09053_, _09131_);
  and _17493_ (_09133_, _09053_, word_in[5]);
  or _17494_ (_09134_, _09133_, _09132_);
  or _17495_ (_09135_, _09134_, _09061_);
  and _17496_ (_09136_, _09135_, _09130_);
  and _17497_ (_09137_, _09046_, word_in[21]);
  or _17498_ (_09138_, _09137_, _09136_);
  and _17499_ (_09139_, _09138_, _09068_);
  and _17500_ (_09140_, _08539_, word_in[29]);
  and _17501_ (_09141_, _09140_, _09044_);
  or _17502_ (_08759_, _09141_, _09139_);
  or _17503_ (_09142_, _09062_, word_in[14]);
  and _17504_ (_09143_, _09142_, _09070_);
  not _17505_ (_09144_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _17506_ (_09145_, _09053_, _09144_);
  and _17507_ (_09146_, _09053_, word_in[6]);
  or _17508_ (_09147_, _09146_, _09145_);
  or _17509_ (_09149_, _09147_, _09061_);
  and _17510_ (_09150_, _09149_, _09143_);
  and _17511_ (_09151_, _09046_, word_in[22]);
  or _17512_ (_09152_, _09151_, _09044_);
  or _17513_ (_09153_, _09152_, _09150_);
  or _17514_ (_09154_, _09068_, word_in[30]);
  and _17515_ (_08763_, _09154_, _09153_);
  or _17516_ (_09155_, _09068_, word_in[31]);
  nor _17517_ (_09156_, _09053_, _08377_);
  and _17518_ (_09157_, _09053_, _08558_);
  or _17519_ (_09158_, _09157_, _09156_);
  or _17520_ (_09159_, _09158_, _09061_);
  or _17521_ (_09160_, _09062_, word_in[15]);
  and _17522_ (_09162_, _09160_, _09070_);
  and _17523_ (_09163_, _09162_, _09159_);
  and _17524_ (_09165_, _08566_, _08699_);
  or _17525_ (_09166_, _09165_, _09044_);
  or _17526_ (_09167_, _09166_, _09163_);
  and _17527_ (_08766_, _09167_, _09155_);
  and _17528_ (_09168_, _08545_, word_in[16]);
  and _17529_ (_09169_, _08545_, _08310_);
  and _17530_ (_09170_, _09169_, _08422_);
  and _17531_ (_09171_, _09170_, _09168_);
  not _17532_ (_09172_, _09170_);
  and _17533_ (_09173_, _08550_, _08328_);
  and _17534_ (_09174_, _09173_, _08321_);
  not _17535_ (_09175_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _17536_ (_09177_, _08553_, _08207_);
  and _17537_ (_09178_, _09177_, _09051_);
  nor _17538_ (_09180_, _09178_, _09175_);
  and _17539_ (_09181_, _09178_, _09056_);
  nor _17540_ (_09182_, _09181_, _09180_);
  nor _17541_ (_09183_, _09182_, _09174_);
  and _17542_ (_09184_, _09174_, word_in[8]);
  or _17543_ (_09185_, _09184_, _09183_);
  and _17544_ (_09187_, _09185_, _09172_);
  or _17545_ (_09188_, _09187_, _09171_);
  and _17546_ (_09189_, _08539_, _08699_);
  not _17547_ (_09190_, _09189_);
  and _17548_ (_09191_, _09190_, _09188_);
  and _17549_ (_09192_, _09189_, word_in[24]);
  or _17550_ (_08846_, _09192_, _09191_);
  and _17551_ (_09194_, _08545_, word_in[17]);
  and _17552_ (_09195_, _09170_, _09194_);
  and _17553_ (_09196_, _09178_, _09080_);
  not _17554_ (_09197_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _17555_ (_09198_, _09178_, _09197_);
  nor _17556_ (_09199_, _09198_, _09196_);
  nor _17557_ (_09200_, _09199_, _09174_);
  and _17558_ (_09201_, _09174_, word_in[9]);
  or _17559_ (_09202_, _09201_, _09200_);
  and _17560_ (_09203_, _09202_, _09172_);
  or _17561_ (_09204_, _09203_, _09195_);
  and _17562_ (_09205_, _09204_, _09190_);
  and _17563_ (_09206_, _09189_, word_in[25]);
  or _17564_ (_08850_, _09206_, _09205_);
  nor _17565_ (_09207_, t2_i, rst);
  and _17566_ (_08853_, _09207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not _17567_ (_09208_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _17568_ (_09209_, _09178_, _09208_);
  and _17569_ (_09210_, _08555_, word_in[2]);
  and _17570_ (_09211_, _09178_, _09210_);
  nor _17571_ (_09212_, _09211_, _09209_);
  nor _17572_ (_09213_, _09212_, _09174_);
  and _17573_ (_09214_, _09174_, word_in[10]);
  or _17574_ (_09215_, _09214_, _09213_);
  and _17575_ (_09216_, _09215_, _09172_);
  and _17576_ (_09217_, _08545_, word_in[18]);
  and _17577_ (_09218_, _09170_, _09217_);
  or _17578_ (_09219_, _09218_, _09216_);
  and _17579_ (_09220_, _09219_, _09190_);
  and _17580_ (_09221_, _09189_, word_in[26]);
  or _17581_ (_08855_, _09221_, _09220_);
  not _17582_ (_09222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _17583_ (_09223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _09222_);
  not _17584_ (_09224_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and _17585_ (_09225_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _17586_ (_09226_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _06445_);
  nor _17587_ (_09227_, _09226_, _09225_);
  nor _17588_ (_09228_, _09227_, _06444_);
  nor _17589_ (_09229_, _09228_, _09224_);
  and _17590_ (_09230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _17591_ (_09231_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _06445_);
  nor _17592_ (_09232_, _09231_, _09230_);
  nor _17593_ (_09233_, _09232_, _06444_);
  not _17594_ (_09234_, _09233_);
  and _17595_ (_09236_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _17596_ (_09237_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _06445_);
  nor _17597_ (_09238_, _09237_, _09236_);
  nor _17598_ (_09239_, _09238_, _06444_);
  and _17599_ (_09240_, _09239_, _09234_);
  nand _17600_ (_09241_, _09240_, _09229_);
  and _17601_ (_09242_, _09241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _17602_ (_09243_, _09242_, _09223_);
  and _17603_ (_09244_, _06032_, _06378_);
  and _17604_ (_09245_, _06840_, _09244_);
  and _17605_ (_09246_, _09245_, _06815_);
  or _17606_ (_09247_, _09246_, _09243_);
  and _17607_ (_09248_, _06383_, _06027_);
  and _17608_ (_09249_, _09248_, _06840_);
  not _17609_ (_09250_, _09249_);
  and _17610_ (_09251_, _09250_, _09247_);
  nand _17611_ (_09252_, _09246_, _06803_);
  and _17612_ (_09254_, _09252_, _09251_);
  nor _17613_ (_09255_, _09250_, _06609_);
  or _17614_ (_09256_, _09255_, _09254_);
  and _17615_ (_08858_, _09256_, _06071_);
  not _17616_ (_09258_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _17617_ (_09259_, _09178_, _09258_);
  and _17618_ (_09260_, _08555_, word_in[3]);
  and _17619_ (_09262_, _09178_, _09260_);
  nor _17620_ (_09263_, _09262_, _09259_);
  nor _17621_ (_09264_, _09263_, _09174_);
  and _17622_ (_09265_, _09174_, word_in[11]);
  or _17623_ (_09267_, _09265_, _09264_);
  and _17624_ (_09268_, _09267_, _09172_);
  and _17625_ (_09269_, _09170_, _09113_);
  or _17626_ (_09271_, _09269_, _09268_);
  and _17627_ (_09272_, _09271_, _09190_);
  and _17628_ (_09273_, _09189_, word_in[27]);
  or _17629_ (_08860_, _09273_, _09272_);
  not _17630_ (_09275_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _17631_ (_09276_, _09178_, _09275_);
  and _17632_ (_09277_, _08555_, word_in[4]);
  and _17633_ (_09279_, _09178_, _09277_);
  or _17634_ (_09280_, _09279_, _09276_);
  or _17635_ (_09282_, _09280_, _09174_);
  not _17636_ (_09283_, _09174_);
  or _17637_ (_09284_, _09283_, word_in[12]);
  and _17638_ (_09285_, _09284_, _09282_);
  and _17639_ (_09286_, _09285_, _09172_);
  and _17640_ (_09287_, _08545_, word_in[20]);
  and _17641_ (_09288_, _09170_, _09287_);
  or _17642_ (_09289_, _09288_, _09286_);
  or _17643_ (_09290_, _09289_, _09189_);
  or _17644_ (_09291_, _09190_, word_in[28]);
  and _17645_ (_08863_, _09291_, _09290_);
  and _17646_ (_09292_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor _17647_ (_09293_, _06967_, _06609_);
  or _17648_ (_09294_, _09293_, _09292_);
  and _17649_ (_08866_, _09294_, _06071_);
  not _17650_ (_09295_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _17651_ (_09296_, _09178_, _09295_);
  and _17652_ (_09297_, _08555_, word_in[5]);
  and _17653_ (_09298_, _09178_, _09297_);
  or _17654_ (_09299_, _09298_, _09296_);
  or _17655_ (_09301_, _09299_, _09174_);
  or _17656_ (_09302_, _09283_, word_in[13]);
  and _17657_ (_09303_, _09302_, _09301_);
  or _17658_ (_09304_, _09303_, _09170_);
  and _17659_ (_09305_, _08545_, word_in[21]);
  or _17660_ (_09306_, _09172_, _09305_);
  and _17661_ (_09307_, _09306_, _09304_);
  or _17662_ (_09308_, _09307_, _09189_);
  or _17663_ (_09309_, _09190_, word_in[29]);
  and _17664_ (_08868_, _09309_, _09308_);
  nor _17665_ (_09310_, _06434_, _06400_);
  and _17666_ (_09311_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _17667_ (_09312_, _09311_, _09310_);
  and _17668_ (_08870_, _09312_, _06071_);
  not _17669_ (_09313_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _17670_ (_09314_, _09178_, _09313_);
  and _17671_ (_09315_, _08555_, word_in[6]);
  and _17672_ (_09316_, _09178_, _09315_);
  nor _17673_ (_09317_, _09316_, _09314_);
  nor _17674_ (_09318_, _09317_, _09174_);
  and _17675_ (_09319_, _09174_, word_in[14]);
  or _17676_ (_09320_, _09319_, _09318_);
  and _17677_ (_09321_, _09320_, _09172_);
  and _17678_ (_09322_, _08545_, word_in[22]);
  and _17679_ (_09323_, _09170_, _09322_);
  or _17680_ (_09324_, _09323_, _09321_);
  and _17681_ (_09325_, _09324_, _09190_);
  and _17682_ (_09326_, _09189_, word_in[30]);
  or _17683_ (_08872_, _09326_, _09325_);
  and _17684_ (_09327_, _09170_, _08566_);
  and _17685_ (_09328_, _09178_, _08558_);
  nor _17686_ (_09329_, _09178_, _08256_);
  nor _17687_ (_09330_, _09329_, _09328_);
  nor _17688_ (_09331_, _09330_, _09174_);
  and _17689_ (_09332_, _09174_, word_in[15]);
  or _17690_ (_09333_, _09332_, _09331_);
  and _17691_ (_09334_, _09333_, _09172_);
  or _17692_ (_09335_, _09334_, _09327_);
  and _17693_ (_09336_, _09335_, _09190_);
  and _17694_ (_09337_, _09189_, word_in[31]);
  or _17695_ (_08875_, _09337_, _09336_);
  nor _17696_ (_09338_, _06355_, _06276_);
  not _17697_ (_09339_, _09338_);
  and _17698_ (_09340_, _09339_, _07410_);
  and _17699_ (_09341_, _09340_, _07388_);
  nor _17700_ (_09342_, _09341_, _06967_);
  and _17701_ (_09343_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _17702_ (_09344_, _09343_, _09342_);
  and _17703_ (_08890_, _09344_, _06071_);
  or _17704_ (_09345_, _06965_, _06391_);
  nor _17705_ (_09346_, _09345_, _06392_);
  or _17706_ (_09347_, _09346_, _06390_);
  and _17707_ (_09348_, _09347_, _06400_);
  or _17708_ (_09349_, _09348_, _06392_);
  and _17709_ (_09350_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _17710_ (_09351_, _07945_, _06400_);
  and _17711_ (_09352_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _17712_ (_09353_, _09352_, _09345_);
  or _17713_ (_09354_, _09353_, _09351_);
  or _17714_ (_09355_, _09354_, _09350_);
  and _17715_ (_08894_, _09355_, _06071_);
  and _17716_ (_09357_, _08545_, _08328_);
  and _17717_ (_09358_, _09357_, _08422_);
  not _17718_ (_09359_, _09358_);
  and _17719_ (_09361_, _08550_, _08308_);
  and _17720_ (_09362_, _09361_, _08321_);
  not _17721_ (_09364_, _08553_);
  and _17722_ (_09365_, _09048_, _09364_);
  and _17723_ (_09367_, _09365_, _09051_);
  and _17724_ (_09368_, _09367_, _09056_);
  not _17725_ (_09369_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _17726_ (_09370_, _09367_, _09369_);
  nor _17727_ (_09372_, _09370_, _09368_);
  nor _17728_ (_09374_, _09372_, _09362_);
  and _17729_ (_09375_, _09362_, word_in[8]);
  or _17730_ (_09377_, _09375_, _09374_);
  and _17731_ (_09378_, _09377_, _09359_);
  and _17732_ (_09380_, _08539_, _08580_);
  and _17733_ (_09381_, _09358_, _09168_);
  or _17734_ (_09382_, _09381_, _09380_);
  or _17735_ (_09383_, _09382_, _09378_);
  not _17736_ (_09384_, _09380_);
  or _17737_ (_09385_, _09384_, word_in[24]);
  and _17738_ (_08960_, _09385_, _09383_);
  not _17739_ (_09386_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _17740_ (_09387_, _09367_, _09386_);
  and _17741_ (_09388_, _09367_, _09080_);
  or _17742_ (_09389_, _09388_, _09387_);
  or _17743_ (_09390_, _09389_, _09362_);
  not _17744_ (_09391_, _09362_);
  or _17745_ (_09392_, _09391_, word_in[9]);
  and _17746_ (_09393_, _09392_, _09390_);
  or _17747_ (_09394_, _09393_, _09358_);
  or _17748_ (_09395_, _09359_, _09194_);
  and _17749_ (_09396_, _09395_, _09384_);
  and _17750_ (_09397_, _09396_, _09394_);
  and _17751_ (_09398_, _09380_, word_in[25]);
  or _17752_ (_08965_, _09398_, _09397_);
  and _17753_ (_09399_, _09367_, _09210_);
  not _17754_ (_09400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _17755_ (_09401_, _09367_, _09400_);
  nor _17756_ (_09402_, _09401_, _09399_);
  nor _17757_ (_09403_, _09402_, _09362_);
  and _17758_ (_09404_, _09362_, word_in[10]);
  or _17759_ (_09405_, _09404_, _09403_);
  and _17760_ (_09406_, _09405_, _09359_);
  and _17761_ (_09407_, _09358_, _09217_);
  or _17762_ (_09408_, _09407_, _09380_);
  or _17763_ (_09409_, _09408_, _09406_);
  or _17764_ (_09410_, _09384_, word_in[26]);
  and _17765_ (_08969_, _09410_, _09409_);
  and _17766_ (_09411_, _09358_, _09113_);
  and _17767_ (_09412_, _09367_, _09260_);
  not _17768_ (_09413_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _17769_ (_09414_, _09367_, _09413_);
  nor _17770_ (_09415_, _09414_, _09412_);
  nor _17771_ (_09416_, _09415_, _09362_);
  and _17772_ (_09417_, _09362_, word_in[11]);
  or _17773_ (_09418_, _09417_, _09416_);
  and _17774_ (_09419_, _09418_, _09359_);
  or _17775_ (_09420_, _09419_, _09411_);
  and _17776_ (_09421_, _09420_, _09384_);
  and _17777_ (_09422_, _09380_, word_in[27]);
  or _17778_ (_08972_, _09422_, _09421_);
  and _17779_ (_09423_, _09367_, _09277_);
  not _17780_ (_09424_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _17781_ (_09425_, _09367_, _09424_);
  nor _17782_ (_09426_, _09425_, _09423_);
  nor _17783_ (_09427_, _09426_, _09362_);
  and _17784_ (_09428_, _09362_, word_in[12]);
  or _17785_ (_09429_, _09428_, _09427_);
  and _17786_ (_09430_, _09429_, _09359_);
  and _17787_ (_09431_, _09358_, _09287_);
  or _17788_ (_09432_, _09431_, _09380_);
  or _17789_ (_09433_, _09432_, _09430_);
  or _17790_ (_09434_, _09384_, word_in[28]);
  and _17791_ (_08976_, _09434_, _09433_);
  not _17792_ (_09435_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _17793_ (_09436_, _09367_, _09435_);
  and _17794_ (_09437_, _09367_, _09297_);
  or _17795_ (_09438_, _09437_, _09436_);
  or _17796_ (_09439_, _09438_, _09362_);
  or _17797_ (_09440_, _09391_, word_in[13]);
  and _17798_ (_09441_, _09440_, _09439_);
  or _17799_ (_09442_, _09441_, _09358_);
  or _17800_ (_09443_, _09359_, _09305_);
  and _17801_ (_09444_, _09443_, _09384_);
  and _17802_ (_09445_, _09444_, _09442_);
  and _17803_ (_09446_, _09380_, word_in[29]);
  or _17804_ (_14026_, _09446_, _09445_);
  and _17805_ (_09447_, _09367_, _09315_);
  not _17806_ (_09448_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _17807_ (_09449_, _09367_, _09448_);
  nor _17808_ (_09450_, _09449_, _09447_);
  nor _17809_ (_09451_, _09450_, _09362_);
  and _17810_ (_09452_, _09362_, word_in[14]);
  or _17811_ (_09453_, _09452_, _09451_);
  and _17812_ (_09454_, _09453_, _09359_);
  and _17813_ (_09455_, _09358_, _09322_);
  or _17814_ (_09456_, _09455_, _09380_);
  or _17815_ (_09457_, _09456_, _09454_);
  or _17816_ (_09458_, _09384_, word_in[30]);
  and _17817_ (_08981_, _09458_, _09457_);
  and _17818_ (_09459_, _09358_, _08566_);
  and _17819_ (_09460_, _09367_, _08558_);
  nor _17820_ (_09461_, _09367_, _08372_);
  nor _17821_ (_09462_, _09461_, _09460_);
  nor _17822_ (_09463_, _09462_, _09362_);
  and _17823_ (_09464_, _09362_, word_in[15]);
  or _17824_ (_09465_, _09464_, _09463_);
  and _17825_ (_09466_, _09465_, _09359_);
  or _17826_ (_09467_, _09466_, _09459_);
  and _17827_ (_09468_, _09467_, _09384_);
  and _17828_ (_09469_, _09380_, word_in[31]);
  or _17829_ (_08983_, _09469_, _09468_);
  and _17830_ (_09470_, _08539_, _08653_);
  not _17831_ (_09471_, _09470_);
  and _17832_ (_09472_, _08545_, _08308_);
  and _17833_ (_09473_, _09472_, _08422_);
  not _17834_ (_09474_, _09473_);
  and _17835_ (_09475_, _08551_, _08321_);
  not _17836_ (_09476_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _17837_ (_09477_, _09051_, _08554_);
  nor _17838_ (_09478_, _09477_, _09476_);
  and _17839_ (_09479_, _09477_, _09056_);
  nor _17840_ (_09480_, _09479_, _09478_);
  nor _17841_ (_09481_, _09480_, _09475_);
  and _17842_ (_09482_, _09475_, word_in[8]);
  or _17843_ (_09483_, _09482_, _09481_);
  and _17844_ (_09484_, _09483_, _09474_);
  and _17845_ (_09485_, _09473_, _09168_);
  or _17846_ (_09486_, _09485_, _09484_);
  and _17847_ (_09487_, _09486_, _09471_);
  and _17848_ (_09488_, _09470_, word_in[24]);
  or _17849_ (_14027_, _09488_, _09487_);
  and _17850_ (_09489_, _09477_, _09080_);
  not _17851_ (_09490_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _17852_ (_09491_, _09477_, _09490_);
  nor _17853_ (_09492_, _09491_, _09489_);
  nor _17854_ (_09493_, _09492_, _09475_);
  and _17855_ (_09494_, _09475_, word_in[9]);
  or _17856_ (_09495_, _09494_, _09493_);
  and _17857_ (_09496_, _09495_, _09474_);
  and _17858_ (_09497_, _09473_, _09194_);
  or _17859_ (_09498_, _09497_, _09496_);
  and _17860_ (_09499_, _09498_, _09471_);
  and _17861_ (_09500_, _09470_, word_in[25]);
  or _17862_ (_09055_, _09500_, _09499_);
  and _17863_ (_09501_, _09477_, _09210_);
  not _17864_ (_09502_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _17865_ (_09503_, _09477_, _09502_);
  nor _17866_ (_09504_, _09503_, _09501_);
  nor _17867_ (_09505_, _09504_, _09475_);
  and _17868_ (_09506_, _09475_, word_in[10]);
  or _17869_ (_09507_, _09506_, _09505_);
  and _17870_ (_09508_, _09507_, _09474_);
  and _17871_ (_09509_, _09473_, _09217_);
  or _17872_ (_09510_, _09509_, _09508_);
  and _17873_ (_09511_, _09510_, _09471_);
  and _17874_ (_09512_, _09470_, word_in[26]);
  or _17875_ (_09058_, _09512_, _09511_);
  not _17876_ (_09513_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _17877_ (_09514_, _09477_, _09513_);
  and _17878_ (_09515_, _09477_, _09260_);
  nor _17879_ (_09516_, _09515_, _09514_);
  nor _17880_ (_09517_, _09516_, _09475_);
  and _17881_ (_09518_, _09475_, word_in[11]);
  or _17882_ (_09519_, _09518_, _09517_);
  and _17883_ (_09520_, _09519_, _09474_);
  and _17884_ (_09521_, _09473_, _09113_);
  or _17885_ (_09522_, _09521_, _09520_);
  and _17886_ (_09523_, _09522_, _09471_);
  and _17887_ (_09524_, _09470_, word_in[27]);
  or _17888_ (_09060_, _09524_, _09523_);
  not _17889_ (_09525_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _17890_ (_09526_, _09477_, _09525_);
  and _17891_ (_09527_, _09477_, _09277_);
  nor _17892_ (_09528_, _09527_, _09526_);
  nor _17893_ (_09529_, _09528_, _09475_);
  and _17894_ (_09530_, _09475_, word_in[12]);
  or _17895_ (_09531_, _09530_, _09529_);
  and _17896_ (_09532_, _09531_, _09474_);
  and _17897_ (_09533_, _09473_, _09287_);
  or _17898_ (_09534_, _09533_, _09532_);
  and _17899_ (_09535_, _09534_, _09471_);
  and _17900_ (_09536_, _09470_, word_in[28]);
  or _17901_ (_09065_, _09536_, _09535_);
  and _17902_ (_09537_, _09477_, _09297_);
  not _17903_ (_09538_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _17904_ (_09539_, _09477_, _09538_);
  nor _17905_ (_09540_, _09539_, _09537_);
  nor _17906_ (_09541_, _09540_, _09475_);
  and _17907_ (_09542_, _09475_, word_in[13]);
  or _17908_ (_09543_, _09542_, _09541_);
  and _17909_ (_09544_, _09543_, _09474_);
  and _17910_ (_09545_, _09473_, _09305_);
  or _17911_ (_09546_, _09545_, _09544_);
  and _17912_ (_09548_, _09546_, _09471_);
  and _17913_ (_09549_, _09470_, word_in[29]);
  or _17914_ (_09069_, _09549_, _09548_);
  not _17915_ (_09550_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _17916_ (_09552_, _09477_, _09550_);
  and _17917_ (_09553_, _09477_, _09315_);
  or _17918_ (_09554_, _09553_, _09552_);
  or _17919_ (_09555_, _09554_, _09475_);
  not _17920_ (_09556_, word_in[14]);
  nand _17921_ (_09557_, _09475_, _09556_);
  and _17922_ (_09558_, _09557_, _09555_);
  or _17923_ (_09559_, _09558_, _09473_);
  or _17924_ (_09560_, _09474_, _09322_);
  and _17925_ (_09561_, _09560_, _09471_);
  and _17926_ (_09562_, _09561_, _09559_);
  and _17927_ (_09563_, _09470_, word_in[30]);
  or _17928_ (_09074_, _09563_, _09562_);
  nor _17929_ (_09564_, _09477_, _08274_);
  and _17930_ (_09565_, _09477_, _08558_);
  nor _17931_ (_09566_, _09565_, _09564_);
  nor _17932_ (_09567_, _09566_, _09475_);
  and _17933_ (_09568_, _09475_, word_in[15]);
  or _17934_ (_09569_, _09568_, _09567_);
  and _17935_ (_09570_, _09569_, _09474_);
  and _17936_ (_09571_, _09473_, _08566_);
  or _17937_ (_09572_, _09571_, _09570_);
  and _17938_ (_09573_, _09572_, _09471_);
  and _17939_ (_09574_, _09470_, word_in[31]);
  or _17940_ (_09077_, _09574_, _09573_);
  and _17941_ (_09575_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _17942_ (_09576_, _07977_, _06390_);
  and _17943_ (_09577_, _09576_, _06398_);
  or _17944_ (_09578_, _09577_, _09575_);
  and _17945_ (_09087_, _09578_, _06071_);
  and _17946_ (_09579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _17947_ (_09580_, _09579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _17948_ (_09581_, _09580_, _07900_);
  and _17949_ (_09582_, _07904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _17950_ (_09583_, _09582_, _09005_);
  or _17951_ (_09584_, _09583_, _09581_);
  and _17952_ (_09585_, _09005_, _09579_);
  or _17953_ (_09586_, _09585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _17954_ (_09587_, _09586_, _06071_);
  and _17955_ (_09148_, _09587_, _09584_);
  and _17956_ (_09588_, _08546_, _08460_);
  and _17957_ (_09589_, _09588_, _08344_);
  not _17958_ (_09590_, _09589_);
  and _17959_ (_09591_, _08550_, _08621_);
  not _17960_ (_09592_, _09591_);
  not _17961_ (_09593_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _17962_ (_09594_, _08555_, _08318_);
  and _17963_ (_09595_, _09594_, _09049_);
  nor _17964_ (_09596_, _09595_, _09593_);
  and _17965_ (_09597_, _09595_, word_in[0]);
  or _17966_ (_09598_, _09597_, _09596_);
  and _17967_ (_09599_, _09598_, _09592_);
  and _17968_ (_09600_, _09591_, word_in[8]);
  or _17969_ (_09601_, _09600_, _09599_);
  and _17970_ (_09602_, _09601_, _09590_);
  and _17971_ (_09603_, _08539_, _08474_);
  and _17972_ (_09604_, _09603_, _08479_);
  and _17973_ (_09605_, _09604_, _08308_);
  and _17974_ (_09606_, _09589_, _09168_);
  or _17975_ (_09607_, _09606_, _09605_);
  or _17976_ (_09608_, _09607_, _09602_);
  not _17977_ (_09609_, _09605_);
  or _17978_ (_09610_, _09609_, _09043_);
  and _17979_ (_09161_, _09610_, _09608_);
  not _17980_ (_09611_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _17981_ (_09612_, _09595_, _09611_);
  and _17982_ (_09613_, _09595_, word_in[1]);
  or _17983_ (_09614_, _09613_, _09612_);
  and _17984_ (_09615_, _09614_, _09592_);
  and _17985_ (_09616_, _09591_, word_in[9]);
  or _17986_ (_09617_, _09616_, _09615_);
  and _17987_ (_09618_, _09617_, _09590_);
  and _17988_ (_09619_, _09589_, _09194_);
  or _17989_ (_09620_, _09619_, _09605_);
  or _17990_ (_09621_, _09620_, _09618_);
  or _17991_ (_09622_, _09609_, _09075_);
  and _17992_ (_09164_, _09622_, _09621_);
  not _17993_ (_09623_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _17994_ (_09624_, _09595_, _09623_);
  and _17995_ (_09625_, _09595_, word_in[2]);
  or _17996_ (_09626_, _09625_, _09624_);
  and _17997_ (_09627_, _09626_, _09592_);
  and _17998_ (_09628_, _09591_, word_in[10]);
  or _17999_ (_09629_, _09628_, _09627_);
  and _18000_ (_09630_, _09629_, _09590_);
  and _18001_ (_09631_, _09589_, _09217_);
  or _18002_ (_09632_, _09631_, _09605_);
  or _18003_ (_09633_, _09632_, _09630_);
  and _18004_ (_09634_, _08539_, word_in[26]);
  or _18005_ (_09635_, _09609_, _09634_);
  and _18006_ (_14028_, _09635_, _09633_);
  not _18007_ (_09636_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _18008_ (_09637_, _09595_, _09636_);
  and _18009_ (_09638_, _09595_, word_in[3]);
  or _18010_ (_09639_, _09638_, _09637_);
  and _18011_ (_09640_, _09639_, _09592_);
  and _18012_ (_09641_, _09591_, word_in[11]);
  or _18013_ (_09642_, _09641_, _09640_);
  and _18014_ (_09643_, _09642_, _09590_);
  and _18015_ (_09644_, _09589_, _09113_);
  or _18016_ (_09645_, _09644_, _09605_);
  or _18017_ (_09646_, _09645_, _09643_);
  or _18018_ (_09647_, _09609_, _09103_);
  and _18019_ (_14029_, _09647_, _09646_);
  not _18020_ (_09648_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _18021_ (_09649_, _09595_, _09648_);
  and _18022_ (_09650_, _09595_, word_in[4]);
  or _18023_ (_09651_, _09650_, _09649_);
  or _18024_ (_09652_, _09651_, _09591_);
  or _18025_ (_09653_, _09592_, word_in[12]);
  and _18026_ (_09654_, _09653_, _09652_);
  and _18027_ (_09655_, _09654_, _09590_);
  and _18028_ (_09656_, _09589_, _09287_);
  or _18029_ (_09657_, _09656_, _09605_);
  or _18030_ (_09658_, _09657_, _09655_);
  and _18031_ (_09659_, _08539_, word_in[28]);
  or _18032_ (_09660_, _09609_, _09659_);
  and _18033_ (_14030_, _09660_, _09658_);
  not _18034_ (_09661_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _18035_ (_09662_, _09595_, _09661_);
  and _18036_ (_09663_, _09595_, word_in[5]);
  or _18037_ (_09664_, _09663_, _09662_);
  and _18038_ (_09665_, _09664_, _09592_);
  and _18039_ (_09666_, _09591_, word_in[13]);
  or _18040_ (_09667_, _09666_, _09665_);
  and _18041_ (_09668_, _09667_, _09590_);
  and _18042_ (_09669_, _09589_, _09305_);
  or _18043_ (_09670_, _09669_, _09605_);
  or _18044_ (_09671_, _09670_, _09668_);
  or _18045_ (_09672_, _09609_, _09140_);
  and _18046_ (_14031_, _09672_, _09671_);
  not _18047_ (_09673_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _18048_ (_09674_, _09595_, _09673_);
  and _18049_ (_09675_, _09595_, word_in[6]);
  or _18050_ (_09676_, _09675_, _09674_);
  and _18051_ (_09677_, _09676_, _09592_);
  and _18052_ (_09678_, _09591_, word_in[14]);
  or _18053_ (_09679_, _09678_, _09677_);
  and _18054_ (_09680_, _09679_, _09590_);
  and _18055_ (_09681_, _09589_, _09322_);
  or _18056_ (_09682_, _09681_, _09605_);
  or _18057_ (_09683_, _09682_, _09680_);
  and _18058_ (_09684_, _08539_, word_in[30]);
  or _18059_ (_09685_, _09609_, _09684_);
  and _18060_ (_09176_, _09685_, _09683_);
  nor _18061_ (_09686_, _09595_, _08390_);
  and _18062_ (_09687_, _09595_, word_in[7]);
  or _18063_ (_09688_, _09687_, _09686_);
  and _18064_ (_09689_, _09688_, _09592_);
  and _18065_ (_09690_, _09591_, word_in[15]);
  or _18066_ (_09691_, _09690_, _09689_);
  and _18067_ (_09692_, _09691_, _09590_);
  and _18068_ (_09693_, _09589_, _08566_);
  or _18069_ (_09694_, _09693_, _09605_);
  or _18070_ (_09695_, _09694_, _09692_);
  or _18071_ (_09696_, _09609_, _08540_);
  and _18072_ (_09179_, _09696_, _09695_);
  nor _18073_ (_09697_, _06527_, _06146_);
  nor _18074_ (_09698_, _05705_, _05865_);
  and _18075_ (_09699_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _18076_ (_09700_, _09699_, _09698_);
  not _18077_ (_09701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor _18078_ (_09702_, _05696_, _09701_);
  and _18079_ (_09703_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _18080_ (_09704_, _09703_, _09702_);
  and _18081_ (_09705_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _18082_ (_09706_, _05718_, _05862_);
  nor _18083_ (_09707_, _09706_, _09705_);
  and _18084_ (_09708_, _09707_, _09704_);
  and _18085_ (_09709_, _09708_, _09700_);
  and _18086_ (_09710_, _06527_, _05811_);
  not _18087_ (_09711_, _09710_);
  nor _18088_ (_09712_, _09711_, _09709_);
  nor _18089_ (_09713_, _09712_, _09697_);
  nor _18090_ (_09186_, _09713_, rst);
  and _18091_ (_09714_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _18092_ (_09715_, _06993_, _06400_);
  and _18093_ (_09716_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _18094_ (_09717_, _09716_, _09345_);
  or _18095_ (_09718_, _09717_, _09715_);
  or _18096_ (_09719_, _09718_, _09714_);
  and _18097_ (_09193_, _09719_, _06071_);
  and _18098_ (_09235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06071_);
  and _18099_ (_09720_, _09604_, _08344_);
  not _18100_ (_09721_, _09720_);
  and _18101_ (_09722_, _09588_, _08310_);
  not _18102_ (_09723_, _09722_);
  or _18103_ (_09724_, _09723_, _09168_);
  and _18104_ (_09725_, _09173_, _08346_);
  not _18105_ (_09726_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _18106_ (_09727_, _09594_, _09177_);
  nor _18107_ (_09728_, _09727_, _09726_);
  and _18108_ (_09729_, _09727_, _09056_);
  or _18109_ (_09730_, _09729_, _09728_);
  or _18110_ (_09731_, _09730_, _09725_);
  not _18111_ (_09732_, _09725_);
  or _18112_ (_09733_, _09732_, word_in[8]);
  and _18113_ (_09734_, _09733_, _09731_);
  or _18114_ (_09735_, _09734_, _09722_);
  and _18115_ (_09736_, _09735_, _09724_);
  and _18116_ (_09737_, _09736_, _09721_);
  and _18117_ (_09738_, _09720_, word_in[24]);
  or _18118_ (_09253_, _09738_, _09737_);
  or _18119_ (_09739_, _09723_, _09194_);
  not _18120_ (_09740_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _18121_ (_09741_, _09727_, _09740_);
  and _18122_ (_09742_, _09727_, _09080_);
  or _18123_ (_09743_, _09742_, _09741_);
  or _18124_ (_09744_, _09743_, _09725_);
  or _18125_ (_09745_, _09732_, word_in[9]);
  and _18126_ (_09746_, _09745_, _09744_);
  or _18127_ (_09747_, _09746_, _09722_);
  and _18128_ (_09748_, _09747_, _09739_);
  or _18129_ (_09749_, _09748_, _09720_);
  or _18130_ (_09750_, _09721_, word_in[25]);
  and _18131_ (_09257_, _09750_, _09749_);
  and _18132_ (_09751_, _09727_, _09210_);
  not _18133_ (_09752_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _18134_ (_09753_, _09727_, _09752_);
  nor _18135_ (_09754_, _09753_, _09751_);
  nor _18136_ (_09755_, _09754_, _09725_);
  and _18137_ (_09756_, _09725_, word_in[10]);
  or _18138_ (_09757_, _09756_, _09755_);
  and _18139_ (_09758_, _09757_, _09723_);
  and _18140_ (_09759_, _09722_, _09217_);
  or _18141_ (_09760_, _09759_, _09720_);
  or _18142_ (_09761_, _09760_, _09758_);
  or _18143_ (_09762_, _09721_, word_in[26]);
  and _18144_ (_09261_, _09762_, _09761_);
  or _18145_ (_09763_, _09723_, _09113_);
  not _18146_ (_09764_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _18147_ (_09765_, _09727_, _09764_);
  and _18148_ (_09766_, _09727_, _09260_);
  or _18149_ (_09767_, _09766_, _09765_);
  or _18150_ (_09768_, _09767_, _09725_);
  or _18151_ (_09769_, _09732_, word_in[11]);
  and _18152_ (_09770_, _09769_, _09768_);
  or _18153_ (_09771_, _09770_, _09722_);
  and _18154_ (_09772_, _09771_, _09763_);
  or _18155_ (_09773_, _09772_, _09720_);
  or _18156_ (_09774_, _09721_, word_in[27]);
  and _18157_ (_09266_, _09774_, _09773_);
  and _18158_ (_09775_, _09727_, _09277_);
  not _18159_ (_09776_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _18160_ (_09777_, _09727_, _09776_);
  nor _18161_ (_09778_, _09777_, _09775_);
  nor _18162_ (_09779_, _09778_, _09725_);
  and _18163_ (_09780_, _09725_, word_in[12]);
  or _18164_ (_09781_, _09780_, _09779_);
  and _18165_ (_09782_, _09781_, _09723_);
  and _18166_ (_09783_, _09722_, _09287_);
  or _18167_ (_09784_, _09783_, _09782_);
  and _18168_ (_09785_, _09784_, _09721_);
  and _18169_ (_09786_, _09720_, word_in[28]);
  or _18170_ (_09270_, _09786_, _09785_);
  not _18171_ (_09787_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _18172_ (_09788_, _09727_, _09787_);
  and _18173_ (_09789_, _09727_, _09297_);
  or _18174_ (_09790_, _09789_, _09788_);
  or _18175_ (_09791_, _09790_, _09725_);
  or _18176_ (_09792_, _09732_, word_in[13]);
  and _18177_ (_09793_, _09792_, _09791_);
  or _18178_ (_09794_, _09793_, _09722_);
  or _18179_ (_09795_, _09723_, _09305_);
  and _18180_ (_09796_, _09795_, _09794_);
  or _18181_ (_09797_, _09796_, _09720_);
  or _18182_ (_09798_, _09721_, word_in[29]);
  and _18183_ (_09274_, _09798_, _09797_);
  or _18184_ (_09799_, _09723_, _09322_);
  not _18185_ (_09800_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _18186_ (_09801_, _09727_, _09800_);
  and _18187_ (_09802_, _09727_, _09315_);
  or _18188_ (_09803_, _09802_, _09801_);
  or _18189_ (_09804_, _09803_, _09725_);
  nand _18190_ (_09805_, _09725_, _09556_);
  and _18191_ (_09806_, _09805_, _09804_);
  or _18192_ (_09807_, _09806_, _09722_);
  and _18193_ (_09808_, _09807_, _09799_);
  or _18194_ (_09809_, _09808_, _09720_);
  or _18195_ (_09810_, _09721_, word_in[30]);
  and _18196_ (_09278_, _09810_, _09809_);
  or _18197_ (_09811_, _09723_, _08566_);
  nor _18198_ (_09812_, _09727_, _08262_);
  and _18199_ (_09813_, _09727_, _08558_);
  or _18200_ (_09814_, _09813_, _09812_);
  or _18201_ (_09815_, _09814_, _09725_);
  or _18202_ (_09816_, _09732_, word_in[15]);
  and _18203_ (_09817_, _09816_, _09815_);
  or _18204_ (_09818_, _09817_, _09722_);
  and _18205_ (_09819_, _09818_, _09811_);
  or _18206_ (_09820_, _09819_, _09720_);
  or _18207_ (_09821_, _09721_, word_in[31]);
  and _18208_ (_09281_, _09821_, _09820_);
  and _18209_ (_09822_, _09588_, _08328_);
  not _18210_ (_09823_, _09822_);
  and _18211_ (_09824_, _09361_, _08346_);
  not _18212_ (_09825_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _18213_ (_09826_, _09365_, _08318_);
  nor _18214_ (_09827_, _09826_, _09825_);
  and _18215_ (_09828_, _09826_, _09056_);
  nor _18216_ (_09829_, _09828_, _09827_);
  nor _18217_ (_09830_, _09829_, _09824_);
  and _18218_ (_09831_, _09824_, word_in[8]);
  or _18219_ (_09832_, _09831_, _09830_);
  and _18220_ (_09833_, _09832_, _09823_);
  and _18221_ (_09834_, _09604_, _08310_);
  and _18222_ (_09835_, _09822_, _09168_);
  or _18223_ (_09836_, _09835_, _09834_);
  or _18224_ (_09837_, _09836_, _09833_);
  not _18225_ (_09838_, _09834_);
  or _18226_ (_09839_, _09838_, word_in[24]);
  and _18227_ (_09356_, _09839_, _09837_);
  or _18228_ (_09840_, _09823_, _09194_);
  not _18229_ (_09841_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _18230_ (_09842_, _09826_, _09841_);
  and _18231_ (_09843_, _09826_, _09080_);
  or _18232_ (_09844_, _09843_, _09842_);
  or _18233_ (_09845_, _09844_, _09824_);
  not _18234_ (_09846_, _09824_);
  or _18235_ (_09847_, _09846_, word_in[9]);
  and _18236_ (_09848_, _09847_, _09845_);
  or _18237_ (_09849_, _09848_, _09822_);
  and _18238_ (_09850_, _09849_, _09840_);
  or _18239_ (_09851_, _09850_, _09834_);
  or _18240_ (_09852_, _09838_, word_in[25]);
  and _18241_ (_09360_, _09852_, _09851_);
  not _18242_ (_09853_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _18243_ (_09854_, _09826_, _09853_);
  and _18244_ (_09855_, _09826_, _09210_);
  or _18245_ (_09856_, _09855_, _09854_);
  or _18246_ (_09857_, _09856_, _09824_);
  or _18247_ (_09858_, _09846_, word_in[10]);
  and _18248_ (_09859_, _09858_, _09857_);
  or _18249_ (_09860_, _09859_, _09822_);
  or _18250_ (_09861_, _09823_, _09217_);
  and _18251_ (_09862_, _09861_, _09860_);
  or _18252_ (_09863_, _09862_, _09834_);
  or _18253_ (_09864_, _09838_, word_in[26]);
  and _18254_ (_09363_, _09864_, _09863_);
  not _18255_ (_09865_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _18256_ (_09866_, _09826_, _09865_);
  and _18257_ (_09867_, _09826_, _09260_);
  or _18258_ (_09868_, _09867_, _09866_);
  or _18259_ (_09869_, _09868_, _09824_);
  or _18260_ (_09870_, _09846_, word_in[11]);
  and _18261_ (_09871_, _09870_, _09869_);
  or _18262_ (_09872_, _09871_, _09822_);
  or _18263_ (_09873_, _09823_, _09113_);
  and _18264_ (_09874_, _09873_, _09872_);
  or _18265_ (_09875_, _09874_, _09834_);
  or _18266_ (_09876_, _09838_, word_in[27]);
  and _18267_ (_09366_, _09876_, _09875_);
  and _18268_ (_09877_, _09826_, _09277_);
  not _18269_ (_09878_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _18270_ (_09879_, _09826_, _09878_);
  nor _18271_ (_09880_, _09879_, _09877_);
  nor _18272_ (_09881_, _09880_, _09824_);
  and _18273_ (_09882_, _09824_, word_in[12]);
  or _18274_ (_09883_, _09882_, _09881_);
  and _18275_ (_09884_, _09883_, _09823_);
  and _18276_ (_09886_, _09822_, _09287_);
  or _18277_ (_09887_, _09886_, _09834_);
  or _18278_ (_09888_, _09887_, _09884_);
  or _18279_ (_09890_, _09838_, word_in[28]);
  and _18280_ (_09371_, _09890_, _09888_);
  not _18281_ (_09891_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _18282_ (_09893_, _09826_, _09891_);
  and _18283_ (_09894_, _09826_, _09297_);
  or _18284_ (_09896_, _09894_, _09893_);
  or _18285_ (_09897_, _09896_, _09824_);
  or _18286_ (_09899_, _09846_, word_in[13]);
  and _18287_ (_09900_, _09899_, _09897_);
  or _18288_ (_09901_, _09900_, _09822_);
  or _18289_ (_09903_, _09823_, _09305_);
  and _18290_ (_09904_, _09903_, _09901_);
  or _18291_ (_09906_, _09904_, _09834_);
  or _18292_ (_09908_, _09838_, word_in[29]);
  and _18293_ (_09373_, _09908_, _09906_);
  and _18294_ (_09909_, _09826_, _09315_);
  not _18295_ (_09910_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _18296_ (_09911_, _09826_, _09910_);
  nor _18297_ (_09912_, _09911_, _09909_);
  nor _18298_ (_09913_, _09912_, _09824_);
  and _18299_ (_09914_, _09824_, word_in[14]);
  or _18300_ (_09915_, _09914_, _09913_);
  and _18301_ (_09916_, _09915_, _09823_);
  and _18302_ (_09917_, _09822_, _09322_);
  or _18303_ (_09918_, _09917_, _09834_);
  or _18304_ (_09919_, _09918_, _09916_);
  or _18305_ (_09920_, _09838_, word_in[30]);
  and _18306_ (_09376_, _09920_, _09919_);
  nor _18307_ (_09921_, _09826_, _08384_);
  and _18308_ (_09922_, _09826_, _08558_);
  nor _18309_ (_09923_, _09922_, _09921_);
  nor _18310_ (_09924_, _09923_, _09824_);
  and _18311_ (_09925_, _09824_, word_in[15]);
  or _18312_ (_09926_, _09925_, _09924_);
  and _18313_ (_09927_, _09926_, _09823_);
  and _18314_ (_09928_, _09822_, _08566_);
  or _18315_ (_09929_, _09928_, _09834_);
  or _18316_ (_09930_, _09929_, _09927_);
  or _18317_ (_09931_, _09838_, word_in[31]);
  and _18318_ (_09379_, _09931_, _09930_);
  and _18319_ (_09932_, _09588_, _08308_);
  and _18320_ (_09933_, _08551_, _08346_);
  and _18321_ (_09934_, _09594_, _08554_);
  and _18322_ (_09935_, _09934_, _09056_);
  not _18323_ (_09936_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _18324_ (_09937_, _09934_, _09936_);
  nor _18325_ (_09938_, _09937_, _09935_);
  nor _18326_ (_09939_, _09938_, _09933_);
  and _18327_ (_09940_, _09933_, word_in[8]);
  or _18328_ (_09941_, _09940_, _09939_);
  or _18329_ (_09942_, _09941_, _09932_);
  and _18330_ (_09943_, _08539_, _08644_);
  not _18331_ (_09944_, _09943_);
  not _18332_ (_09945_, _09932_);
  or _18333_ (_09946_, _09945_, _09168_);
  and _18334_ (_09947_, _09946_, _09944_);
  and _18335_ (_09948_, _09947_, _09942_);
  and _18336_ (_09949_, _09043_, _08644_);
  or _18337_ (_14032_, _09949_, _09948_);
  not _18338_ (_09950_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _18339_ (_09951_, _09934_, _09950_);
  and _18340_ (_09952_, _09934_, _09080_);
  or _18341_ (_09953_, _09952_, _09951_);
  or _18342_ (_09954_, _09953_, _09933_);
  not _18343_ (_09955_, _09933_);
  or _18344_ (_09956_, _09955_, word_in[9]);
  and _18345_ (_09957_, _09956_, _09954_);
  or _18346_ (_09958_, _09957_, _09932_);
  or _18347_ (_09959_, _09945_, _09194_);
  and _18348_ (_09960_, _09959_, _09958_);
  or _18349_ (_09961_, _09960_, _09943_);
  or _18350_ (_09962_, _09944_, word_in[25]);
  and _18351_ (_14033_, _09962_, _09961_);
  and _18352_ (_09963_, _09634_, _08644_);
  and _18353_ (_09964_, _09934_, _09210_);
  not _18354_ (_09965_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _18355_ (_09966_, _09934_, _09965_);
  nor _18356_ (_09967_, _09966_, _09964_);
  nor _18357_ (_09968_, _09967_, _09933_);
  and _18358_ (_09969_, _09933_, word_in[10]);
  or _18359_ (_09970_, _09969_, _09968_);
  and _18360_ (_09971_, _09970_, _09945_);
  and _18361_ (_09972_, _09932_, _09217_);
  or _18362_ (_09973_, _09972_, _09971_);
  and _18363_ (_09974_, _09973_, _09944_);
  or _18364_ (_14034_, _09974_, _09963_);
  and _18365_ (_09975_, _09103_, _08644_);
  not _18366_ (_09976_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _18367_ (_09977_, _09934_, _09976_);
  and _18368_ (_09978_, _09934_, _09260_);
  or _18369_ (_09979_, _09978_, _09977_);
  or _18370_ (_09980_, _09979_, _09933_);
  or _18371_ (_09981_, _09955_, word_in[11]);
  and _18372_ (_09982_, _09981_, _09980_);
  or _18373_ (_09984_, _09982_, _09932_);
  or _18374_ (_09986_, _09945_, _09113_);
  and _18375_ (_09987_, _09986_, _09944_);
  and _18376_ (_09988_, _09987_, _09984_);
  or _18377_ (_14035_, _09988_, _09975_);
  and _18378_ (_09990_, _09943_, word_in[28]);
  not _18379_ (_09991_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _18380_ (_09992_, _09934_, _09991_);
  and _18381_ (_09993_, _09934_, _09277_);
  or _18382_ (_09995_, _09993_, _09992_);
  or _18383_ (_09997_, _09995_, _09933_);
  or _18384_ (_09998_, _09955_, word_in[12]);
  and _18385_ (_09999_, _09998_, _09997_);
  or _18386_ (_10000_, _09999_, _09932_);
  or _18387_ (_10002_, _09945_, _09287_);
  and _18388_ (_10003_, _10002_, _09944_);
  and _18389_ (_10004_, _10003_, _10000_);
  or _18390_ (_14036_, _10004_, _09990_);
  and _18391_ (_10006_, _09140_, _08644_);
  and _18392_ (_10007_, _09934_, _09297_);
  not _18393_ (_10008_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _18394_ (_10010_, _09934_, _10008_);
  nor _18395_ (_10011_, _10010_, _10007_);
  nor _18396_ (_10012_, _10011_, _09933_);
  and _18397_ (_10013_, _09933_, word_in[13]);
  or _18398_ (_10014_, _10013_, _10012_);
  and _18399_ (_10015_, _10014_, _09945_);
  and _18400_ (_10016_, _09932_, _09305_);
  or _18401_ (_10017_, _10016_, _10015_);
  and _18402_ (_10018_, _10017_, _09944_);
  or _18403_ (_14037_, _10018_, _10006_);
  not _18404_ (_10019_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _18405_ (_10020_, _09934_, _10019_);
  and _18406_ (_10021_, _09934_, _09315_);
  or _18407_ (_10022_, _10021_, _10020_);
  or _18408_ (_10023_, _10022_, _09933_);
  nand _18409_ (_10024_, _09933_, _09556_);
  and _18410_ (_10025_, _10024_, _10023_);
  or _18411_ (_10026_, _10025_, _09932_);
  or _18412_ (_10027_, _09945_, _09322_);
  and _18413_ (_10028_, _10027_, _09944_);
  and _18414_ (_10029_, _10028_, _10026_);
  and _18415_ (_10030_, _09943_, word_in[30]);
  or _18416_ (_14038_, _10030_, _10029_);
  and _18417_ (_10031_, _09934_, _08558_);
  nor _18418_ (_10033_, _09934_, _08268_);
  nor _18419_ (_10034_, _10033_, _10031_);
  nor _18420_ (_10035_, _10034_, _09933_);
  and _18421_ (_10036_, _09933_, word_in[15]);
  or _18422_ (_10037_, _10036_, _10035_);
  and _18423_ (_10038_, _10037_, _09945_);
  and _18424_ (_10039_, _09932_, _08566_);
  or _18425_ (_10040_, _10039_, _10038_);
  and _18426_ (_10041_, _10040_, _09944_);
  and _18427_ (_10042_, _09943_, word_in[31]);
  or _18428_ (_14039_, _10042_, _10041_);
  and _18429_ (_10043_, _08539_, _08482_);
  and _18430_ (_10044_, _10043_, _08308_);
  not _18431_ (_10045_, _10044_);
  and _18432_ (_10046_, _08545_, _08428_);
  not _18433_ (_10047_, _10046_);
  or _18434_ (_10048_, _10047_, word_in[16]);
  and _18435_ (_10049_, _08550_, _08319_);
  not _18436_ (_10050_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18437_ (_10051_, _08317_, _08184_);
  and _18438_ (_10052_, _08555_, _10051_);
  and _18439_ (_10053_, _10052_, _09049_);
  nor _18440_ (_10054_, _10053_, _10050_);
  and _18441_ (_10055_, _10053_, _09056_);
  or _18442_ (_10056_, _10055_, _10054_);
  or _18443_ (_10057_, _10056_, _10049_);
  not _18444_ (_10058_, _10049_);
  or _18445_ (_10059_, _10058_, word_in[8]);
  and _18446_ (_10060_, _10059_, _10057_);
  or _18447_ (_10061_, _10060_, _10046_);
  and _18448_ (_10062_, _10061_, _10048_);
  and _18449_ (_10063_, _10062_, _10045_);
  and _18450_ (_10064_, _10044_, word_in[24]);
  or _18451_ (_09547_, _10064_, _10063_);
  and _18452_ (_10065_, _10046_, word_in[17]);
  not _18453_ (_10066_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _18454_ (_10067_, _10053_, _10066_);
  and _18455_ (_10068_, _10053_, word_in[1]);
  or _18456_ (_10069_, _10068_, _10067_);
  and _18457_ (_10070_, _10069_, _10058_);
  and _18458_ (_10071_, _10049_, word_in[9]);
  or _18459_ (_10072_, _10071_, _10070_);
  and _18460_ (_10073_, _10072_, _10047_);
  or _18461_ (_10074_, _10073_, _10065_);
  and _18462_ (_10075_, _10074_, _10045_);
  and _18463_ (_10076_, _10044_, word_in[25]);
  or _18464_ (_09551_, _10076_, _10075_);
  and _18465_ (_10078_, _10046_, word_in[18]);
  not _18466_ (_10079_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _18467_ (_10080_, _10053_, _10079_);
  and _18468_ (_10082_, _10053_, word_in[2]);
  or _18469_ (_10083_, _10082_, _10080_);
  and _18470_ (_10084_, _10083_, _10058_);
  and _18471_ (_10085_, _10049_, word_in[10]);
  or _18472_ (_10087_, _10085_, _10084_);
  and _18473_ (_10088_, _10087_, _10047_);
  or _18474_ (_10089_, _10088_, _10078_);
  and _18475_ (_10090_, _10089_, _10045_);
  and _18476_ (_10092_, _10044_, word_in[26]);
  or _18477_ (_14040_, _10092_, _10090_);
  and _18478_ (_10093_, _10046_, word_in[19]);
  not _18479_ (_10095_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _18480_ (_10096_, _10053_, _10095_);
  and _18481_ (_10097_, _10053_, word_in[3]);
  or _18482_ (_10098_, _10097_, _10096_);
  and _18483_ (_10100_, _10098_, _10058_);
  and _18484_ (_10101_, _10049_, word_in[11]);
  or _18485_ (_10102_, _10101_, _10100_);
  and _18486_ (_10103_, _10102_, _10047_);
  or _18487_ (_10105_, _10103_, _10093_);
  and _18488_ (_10107_, _10105_, _10045_);
  and _18489_ (_10108_, _10044_, word_in[27]);
  or _18490_ (_14041_, _10108_, _10107_);
  and _18491_ (_10109_, _10046_, word_in[20]);
  not _18492_ (_10110_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _18493_ (_10111_, _10053_, _10110_);
  and _18494_ (_10112_, _10053_, word_in[4]);
  or _18495_ (_10113_, _10112_, _10111_);
  and _18496_ (_10114_, _10113_, _10058_);
  and _18497_ (_10115_, _10049_, word_in[12]);
  or _18498_ (_10116_, _10115_, _10114_);
  and _18499_ (_10117_, _10116_, _10047_);
  or _18500_ (_10118_, _10117_, _10109_);
  and _18501_ (_10119_, _10118_, _10045_);
  and _18502_ (_10120_, _10044_, word_in[28]);
  or _18503_ (_14042_, _10120_, _10119_);
  not _18504_ (_10121_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _18505_ (_10122_, _10053_, _10121_);
  and _18506_ (_10123_, _10053_, word_in[5]);
  or _18507_ (_10124_, _10123_, _10122_);
  and _18508_ (_10125_, _10124_, _10058_);
  and _18509_ (_10126_, _10049_, word_in[13]);
  or _18510_ (_10127_, _10126_, _10125_);
  and _18511_ (_10128_, _10127_, _10047_);
  and _18512_ (_10129_, _10046_, word_in[21]);
  or _18513_ (_10130_, _10129_, _10128_);
  and _18514_ (_10131_, _10130_, _10045_);
  and _18515_ (_10132_, _10044_, word_in[29]);
  or _18516_ (_14043_, _10132_, _10131_);
  and _18517_ (_10133_, _10046_, word_in[22]);
  not _18518_ (_10134_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _18519_ (_10135_, _10053_, _10134_);
  and _18520_ (_10136_, _10053_, word_in[6]);
  or _18521_ (_10137_, _10136_, _10135_);
  and _18522_ (_10138_, _10137_, _10058_);
  and _18523_ (_10139_, _10049_, word_in[14]);
  or _18524_ (_10140_, _10139_, _10138_);
  and _18525_ (_10141_, _10140_, _10047_);
  or _18526_ (_10142_, _10141_, _10133_);
  and _18527_ (_10143_, _10142_, _10045_);
  and _18528_ (_10144_, _10044_, word_in[30]);
  or _18529_ (_14044_, _10144_, _10143_);
  and _18530_ (_10145_, _10046_, word_in[23]);
  nor _18531_ (_10146_, _10053_, _08365_);
  and _18532_ (_10147_, _10053_, word_in[7]);
  or _18533_ (_10148_, _10147_, _10146_);
  and _18534_ (_10149_, _10148_, _10058_);
  and _18535_ (_10150_, _10049_, word_in[15]);
  or _18536_ (_10151_, _10150_, _10149_);
  and _18537_ (_10152_, _10151_, _10047_);
  or _18538_ (_10153_, _10152_, _10145_);
  and _18539_ (_10154_, _10153_, _10045_);
  and _18540_ (_10155_, _10044_, word_in[31]);
  or _18541_ (_14045_, _10155_, _10154_);
  and _18542_ (_10156_, _09169_, _08420_);
  not _18543_ (_10157_, _10156_);
  and _18544_ (_10158_, _09173_, _08323_);
  and _18545_ (_10159_, _10052_, _09177_);
  and _18546_ (_10160_, _10159_, _09056_);
  not _18547_ (_10161_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _18548_ (_10162_, _10159_, _10161_);
  nor _18549_ (_10163_, _10162_, _10160_);
  nor _18550_ (_10164_, _10163_, _10158_);
  and _18551_ (_10165_, _10158_, word_in[8]);
  or _18552_ (_10166_, _10165_, _10164_);
  and _18553_ (_10167_, _10166_, _10157_);
  and _18554_ (_10168_, _10043_, _08344_);
  and _18555_ (_10169_, _10156_, _09168_);
  or _18556_ (_10171_, _10169_, _10168_);
  or _18557_ (_10172_, _10171_, _10167_);
  not _18558_ (_10173_, _10168_);
  or _18559_ (_10175_, _10173_, _09043_);
  and _18560_ (_14046_, _10175_, _10172_);
  not _18561_ (_10177_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _18562_ (_10179_, _10159_, _10177_);
  and _18563_ (_10181_, _10159_, _09080_);
  or _18564_ (_10182_, _10181_, _10179_);
  or _18565_ (_10183_, _10182_, _10158_);
  not _18566_ (_10185_, _10158_);
  or _18567_ (_10186_, _10185_, word_in[9]);
  and _18568_ (_10188_, _10186_, _10183_);
  or _18569_ (_10189_, _10188_, _10156_);
  or _18570_ (_10191_, _10157_, _09194_);
  and _18571_ (_10192_, _10191_, _10173_);
  and _18572_ (_10193_, _10192_, _10189_);
  and _18573_ (_10194_, _10168_, _09075_);
  or _18574_ (_14047_, _10194_, _10193_);
  not _18575_ (_10195_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _18576_ (_10196_, _10159_, _10195_);
  and _18577_ (_10197_, _10159_, _09210_);
  or _18578_ (_10198_, _10197_, _10196_);
  or _18579_ (_10199_, _10198_, _10158_);
  or _18580_ (_10200_, _10185_, word_in[10]);
  and _18581_ (_10201_, _10200_, _10199_);
  or _18582_ (_10202_, _10201_, _10156_);
  or _18583_ (_10203_, _10157_, _09217_);
  and _18584_ (_10204_, _10203_, _10173_);
  and _18585_ (_10205_, _10204_, _10202_);
  and _18586_ (_10206_, _10168_, _09634_);
  or _18587_ (_14048_, _10206_, _10205_);
  and _18588_ (_10207_, _10159_, _09260_);
  not _18589_ (_10208_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _18590_ (_10209_, _10159_, _10208_);
  nor _18591_ (_10210_, _10209_, _10207_);
  nor _18592_ (_10211_, _10210_, _10158_);
  and _18593_ (_10212_, _10158_, word_in[11]);
  or _18594_ (_10213_, _10212_, _10211_);
  and _18595_ (_10214_, _10213_, _10157_);
  and _18596_ (_10215_, _10156_, _09113_);
  or _18597_ (_10216_, _10215_, _10168_);
  or _18598_ (_10217_, _10216_, _10214_);
  or _18599_ (_10218_, _10173_, _09103_);
  and _18600_ (_14049_, _10218_, _10217_);
  and _18601_ (_10219_, _10159_, _09277_);
  not _18602_ (_10220_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _18603_ (_10221_, _10159_, _10220_);
  nor _18604_ (_10222_, _10221_, _10219_);
  nor _18605_ (_10223_, _10222_, _10158_);
  and _18606_ (_10224_, _10158_, word_in[12]);
  or _18607_ (_10225_, _10224_, _10223_);
  and _18608_ (_10226_, _10225_, _10157_);
  and _18609_ (_10227_, _10156_, _09287_);
  or _18610_ (_10228_, _10227_, _10168_);
  or _18611_ (_10229_, _10228_, _10226_);
  or _18612_ (_10230_, _10173_, _09659_);
  and _18613_ (_14050_, _10230_, _10229_);
  and _18614_ (_10231_, _10159_, _09297_);
  not _18615_ (_10232_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _18616_ (_10233_, _10159_, _10232_);
  nor _18617_ (_10234_, _10233_, _10231_);
  nor _18618_ (_10235_, _10234_, _10158_);
  and _18619_ (_10236_, _10158_, word_in[13]);
  or _18620_ (_10237_, _10236_, _10235_);
  and _18621_ (_10238_, _10237_, _10157_);
  and _18622_ (_10239_, _10156_, _09305_);
  or _18623_ (_10240_, _10239_, _10168_);
  or _18624_ (_10241_, _10240_, _10238_);
  or _18625_ (_10242_, _10173_, _09140_);
  and _18626_ (_14051_, _10242_, _10241_);
  and _18627_ (_10243_, _10159_, _09315_);
  not _18628_ (_10244_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _18629_ (_10245_, _10159_, _10244_);
  nor _18630_ (_10246_, _10245_, _10243_);
  nor _18631_ (_10247_, _10246_, _10158_);
  and _18632_ (_10248_, _10158_, word_in[14]);
  or _18633_ (_10249_, _10248_, _10247_);
  and _18634_ (_10250_, _10249_, _10157_);
  and _18635_ (_10251_, _10156_, _09322_);
  or _18636_ (_10252_, _10251_, _10168_);
  or _18637_ (_10253_, _10252_, _10250_);
  or _18638_ (_10254_, _10173_, _09684_);
  and _18639_ (_14052_, _10254_, _10253_);
  and _18640_ (_10255_, _10159_, _08558_);
  nor _18641_ (_10256_, _10159_, _08282_);
  nor _18642_ (_10257_, _10256_, _10255_);
  nor _18643_ (_10258_, _10257_, _10158_);
  and _18644_ (_10259_, _10158_, word_in[15]);
  or _18645_ (_10260_, _10259_, _10258_);
  and _18646_ (_10261_, _10260_, _10157_);
  and _18647_ (_10262_, _10156_, _08566_);
  or _18648_ (_10263_, _10262_, _10168_);
  or _18649_ (_10264_, _10263_, _10261_);
  or _18650_ (_10265_, _10173_, _08540_);
  and _18651_ (_14053_, _10265_, _10264_);
  and _18652_ (_10266_, _10043_, _08310_);
  and _18653_ (_10267_, _09357_, _08420_);
  and _18654_ (_10268_, _09361_, _08323_);
  not _18655_ (_10269_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18656_ (_10270_, _10052_, _09365_);
  nor _18657_ (_10271_, _10270_, _10269_);
  and _18658_ (_10272_, _10270_, _09056_);
  or _18659_ (_10273_, _10272_, _10271_);
  or _18660_ (_10274_, _10273_, _10268_);
  not _18661_ (_10275_, _10268_);
  or _18662_ (_10276_, _10275_, word_in[8]);
  and _18663_ (_10277_, _10276_, _10274_);
  or _18664_ (_10278_, _10277_, _10267_);
  not _18665_ (_10279_, _10267_);
  or _18666_ (_10280_, _10279_, _09168_);
  and _18667_ (_10281_, _10280_, _10278_);
  or _18668_ (_10282_, _10281_, _10266_);
  not _18669_ (_10283_, _10266_);
  or _18670_ (_10284_, _10283_, word_in[24]);
  and _18671_ (_14008_, _10284_, _10282_);
  not _18672_ (_10285_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _18673_ (_10286_, _10270_, _10285_);
  and _18674_ (_10287_, _10270_, _09080_);
  or _18675_ (_10288_, _10287_, _10286_);
  or _18676_ (_10289_, _10288_, _10268_);
  or _18677_ (_10290_, _10275_, word_in[9]);
  and _18678_ (_10291_, _10290_, _10289_);
  or _18679_ (_10292_, _10291_, _10267_);
  or _18680_ (_10293_, _10279_, _09194_);
  and _18681_ (_10294_, _10293_, _10283_);
  and _18682_ (_10295_, _10294_, _10292_);
  and _18683_ (_10296_, _10266_, word_in[25]);
  or _18684_ (_14009_, _10296_, _10295_);
  and _18685_ (_10297_, _10270_, _09210_);
  not _18686_ (_10298_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _18687_ (_10299_, _10270_, _10298_);
  nor _18688_ (_10300_, _10299_, _10297_);
  nor _18689_ (_10301_, _10300_, _10268_);
  and _18690_ (_10302_, _10268_, word_in[10]);
  or _18691_ (_10303_, _10302_, _10301_);
  and _18692_ (_10304_, _10303_, _10279_);
  and _18693_ (_10305_, _10267_, _09217_);
  or _18694_ (_10306_, _10305_, _10266_);
  or _18695_ (_10307_, _10306_, _10304_);
  or _18696_ (_10308_, _10283_, word_in[26]);
  and _18697_ (_14010_, _10308_, _10307_);
  and _18698_ (_10309_, _10270_, _09260_);
  not _18699_ (_10310_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _18700_ (_10311_, _10270_, _10310_);
  nor _18701_ (_10312_, _10311_, _10309_);
  nor _18702_ (_10313_, _10312_, _10268_);
  and _18703_ (_10314_, _10268_, word_in[11]);
  or _18704_ (_10315_, _10314_, _10313_);
  and _18705_ (_10316_, _10315_, _10279_);
  and _18706_ (_10317_, _10267_, _09113_);
  or _18707_ (_10318_, _10317_, _10266_);
  or _18708_ (_10319_, _10318_, _10316_);
  or _18709_ (_10320_, _10283_, word_in[27]);
  and _18710_ (_14011_, _10320_, _10319_);
  and _18711_ (_10321_, _10267_, _09287_);
  and _18712_ (_10322_, _10270_, _09277_);
  not _18713_ (_10323_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _18714_ (_10324_, _10270_, _10323_);
  nor _18715_ (_10325_, _10324_, _10322_);
  nor _18716_ (_10326_, _10325_, _10268_);
  and _18717_ (_10327_, _10268_, word_in[12]);
  or _18718_ (_10328_, _10327_, _10326_);
  and _18719_ (_10329_, _10328_, _10279_);
  or _18720_ (_10330_, _10329_, _10321_);
  and _18721_ (_10331_, _10330_, _10283_);
  and _18722_ (_10332_, _10266_, word_in[28]);
  or _18723_ (_14012_, _10332_, _10331_);
  and _18724_ (_10333_, _10270_, _09297_);
  not _18725_ (_10334_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _18726_ (_10335_, _10270_, _10334_);
  nor _18727_ (_10336_, _10335_, _10333_);
  nor _18728_ (_10337_, _10336_, _10268_);
  and _18729_ (_10338_, _10268_, word_in[13]);
  or _18730_ (_10339_, _10338_, _10337_);
  and _18731_ (_10340_, _10339_, _10279_);
  and _18732_ (_10341_, _10267_, _09305_);
  or _18733_ (_10342_, _10341_, _10266_);
  or _18734_ (_10343_, _10342_, _10340_);
  or _18735_ (_10344_, _10283_, word_in[29]);
  and _18736_ (_14013_, _10344_, _10343_);
  and _18737_ (_10345_, _10270_, _09315_);
  not _18738_ (_10346_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _18739_ (_10347_, _10270_, _10346_);
  nor _18740_ (_10348_, _10347_, _10345_);
  nor _18741_ (_10349_, _10348_, _10268_);
  and _18742_ (_10350_, _10268_, word_in[14]);
  or _18743_ (_10351_, _10350_, _10349_);
  and _18744_ (_10352_, _10351_, _10279_);
  and _18745_ (_10353_, _10267_, _09322_);
  or _18746_ (_10354_, _10353_, _10266_);
  or _18747_ (_10355_, _10354_, _10352_);
  or _18748_ (_10356_, _10283_, word_in[30]);
  and _18749_ (_14014_, _10356_, _10355_);
  nor _18750_ (_10357_, _10270_, _08360_);
  and _18751_ (_10358_, _10270_, _08558_);
  or _18752_ (_10359_, _10358_, _10357_);
  or _18753_ (_10360_, _10359_, _10268_);
  or _18754_ (_10361_, _10275_, word_in[15]);
  and _18755_ (_10362_, _10361_, _10360_);
  or _18756_ (_10363_, _10362_, _10267_);
  or _18757_ (_10364_, _10279_, _08566_);
  and _18758_ (_10365_, _10364_, _10363_);
  and _18759_ (_10366_, _10365_, _10283_);
  and _18760_ (_10367_, _10266_, word_in[31]);
  or _18761_ (_14015_, _10367_, _10366_);
  and _18762_ (_10368_, _09472_, _08420_);
  not _18763_ (_10369_, _10368_);
  and _18764_ (_10370_, _08551_, _08323_);
  not _18765_ (_10371_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _18766_ (_10372_, _10052_, _08554_);
  nor _18767_ (_10373_, _10372_, _10371_);
  and _18768_ (_10374_, _10372_, _09056_);
  or _18769_ (_10375_, _10374_, _10373_);
  or _18770_ (_10376_, _10375_, _10370_);
  not _18771_ (_10377_, _10370_);
  or _18772_ (_10378_, _10377_, word_in[8]);
  and _18773_ (_10379_, _10378_, _10376_);
  and _18774_ (_10380_, _10379_, _10369_);
  and _18775_ (_10381_, _10043_, _08328_);
  and _18776_ (_10382_, _10368_, _09168_);
  or _18777_ (_10383_, _10382_, _10381_);
  or _18778_ (_10384_, _10383_, _10380_);
  not _18779_ (_10385_, _10381_);
  or _18780_ (_10386_, _10385_, word_in[24]);
  and _18781_ (_14016_, _10386_, _10384_);
  not _18782_ (_10387_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _18783_ (_10388_, _10372_, _10387_);
  and _18784_ (_10389_, _10372_, _09080_);
  or _18785_ (_10390_, _10389_, _10388_);
  or _18786_ (_10391_, _10390_, _10370_);
  or _18787_ (_10392_, _10377_, word_in[9]);
  and _18788_ (_10393_, _10392_, _10391_);
  or _18789_ (_10394_, _10393_, _10368_);
  or _18790_ (_10395_, _10369_, _09194_);
  and _18791_ (_10396_, _10395_, _10394_);
  or _18792_ (_10397_, _10396_, _10381_);
  or _18793_ (_10398_, _10385_, word_in[25]);
  and _18794_ (_14017_, _10398_, _10397_);
  not _18795_ (_10399_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _18796_ (_10400_, _10372_, _10399_);
  and _18797_ (_10401_, _10372_, _09210_);
  or _18798_ (_10402_, _10401_, _10400_);
  or _18799_ (_10403_, _10402_, _10370_);
  or _18800_ (_10404_, _10377_, word_in[10]);
  and _18801_ (_10405_, _10404_, _10403_);
  or _18802_ (_10406_, _10405_, _10368_);
  or _18803_ (_10407_, _10369_, _09217_);
  and _18804_ (_10408_, _10407_, _10385_);
  and _18805_ (_10409_, _10408_, _10406_);
  and _18806_ (_10410_, _10381_, _09634_);
  or _18807_ (_14018_, _10410_, _10409_);
  and _18808_ (_10411_, _10372_, _09260_);
  not _18809_ (_10412_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _18810_ (_10413_, _10372_, _10412_);
  nor _18811_ (_10414_, _10413_, _10411_);
  nor _18812_ (_10415_, _10414_, _10370_);
  and _18813_ (_10416_, _10370_, word_in[11]);
  or _18814_ (_10417_, _10416_, _10415_);
  and _18815_ (_10418_, _10417_, _10369_);
  and _18816_ (_10420_, _10368_, _09113_);
  or _18817_ (_10421_, _10420_, _10381_);
  or _18818_ (_10422_, _10421_, _10418_);
  or _18819_ (_10423_, _10385_, _09103_);
  and _18820_ (_14019_, _10423_, _10422_);
  not _18821_ (_10425_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _18822_ (_10426_, _10372_, _10425_);
  and _18823_ (_10428_, _10372_, _09277_);
  or _18824_ (_10429_, _10428_, _10426_);
  or _18825_ (_10431_, _10429_, _10370_);
  or _18826_ (_10432_, _10377_, word_in[12]);
  and _18827_ (_10434_, _10432_, _10431_);
  or _18828_ (_10435_, _10434_, _10368_);
  or _18829_ (_10436_, _10369_, _09287_);
  and _18830_ (_10437_, _10436_, _10385_);
  and _18831_ (_10438_, _10437_, _10435_);
  and _18832_ (_10439_, _10381_, _09659_);
  or _18833_ (_14020_, _10439_, _10438_);
  and _18834_ (_10440_, _10372_, _09297_);
  not _18835_ (_10441_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _18836_ (_10442_, _10372_, _10441_);
  nor _18837_ (_10443_, _10442_, _10440_);
  nor _18838_ (_10444_, _10443_, _10370_);
  and _18839_ (_10445_, _10370_, word_in[13]);
  or _18840_ (_10446_, _10445_, _10444_);
  and _18841_ (_10447_, _10446_, _10369_);
  and _18842_ (_10448_, _10368_, _09305_);
  or _18843_ (_10450_, _10448_, _10381_);
  or _18844_ (_10451_, _10450_, _10447_);
  or _18845_ (_10452_, _10385_, _09140_);
  and _18846_ (_14021_, _10452_, _10451_);
  and _18847_ (_10453_, _10372_, _09315_);
  not _18848_ (_10454_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _18849_ (_10455_, _10372_, _10454_);
  nor _18850_ (_10456_, _10455_, _10453_);
  nor _18851_ (_10457_, _10456_, _10370_);
  and _18852_ (_10458_, _10370_, word_in[14]);
  or _18853_ (_10460_, _10458_, _10457_);
  and _18854_ (_10461_, _10460_, _10369_);
  and _18855_ (_10462_, _10368_, _09322_);
  or _18856_ (_10463_, _10462_, _10381_);
  or _18857_ (_10464_, _10463_, _10461_);
  or _18858_ (_10465_, _10385_, _09684_);
  and _18859_ (_14022_, _10465_, _10464_);
  nor _18860_ (_10466_, _10372_, _08299_);
  and _18861_ (_10467_, _10372_, _08558_);
  or _18862_ (_10468_, _10467_, _10466_);
  or _18863_ (_10469_, _10468_, _10370_);
  or _18864_ (_10470_, _10377_, word_in[15]);
  and _18865_ (_10471_, _10470_, _10469_);
  or _18866_ (_10472_, _10471_, _10368_);
  or _18867_ (_10473_, _10369_, _08566_);
  and _18868_ (_10474_, _10473_, _10385_);
  and _18869_ (_10475_, _10474_, _10472_);
  and _18870_ (_10476_, _10381_, _08540_);
  or _18871_ (_14023_, _10476_, _10475_);
  and _18872_ (_10477_, _08547_, _08344_);
  not _18873_ (_10478_, _10477_);
  and _18874_ (_10479_, _08522_, _08310_);
  and _18875_ (_10481_, _08550_, _10479_);
  not _18876_ (_10483_, _10481_);
  not _18877_ (_10484_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _18878_ (_10485_, _09049_, _08556_);
  nor _18879_ (_10486_, _10485_, _10484_);
  and _18880_ (_10487_, _10485_, word_in[0]);
  or _18881_ (_10488_, _10487_, _10486_);
  and _18882_ (_10489_, _10488_, _10483_);
  and _18883_ (_10490_, _10481_, word_in[8]);
  or _18884_ (_10491_, _10490_, _10489_);
  and _18885_ (_10492_, _10491_, _10478_);
  not _18886_ (_10493_, _08479_);
  and _18887_ (_10494_, _09603_, _10493_);
  and _18888_ (_10495_, _10494_, _08308_);
  and _18889_ (_10496_, _10477_, _09168_);
  or _18890_ (_10497_, _10496_, _10495_);
  or _18891_ (_10498_, _10497_, _10492_);
  not _18892_ (_10499_, _10495_);
  or _18893_ (_10500_, _10499_, _09043_);
  and _18894_ (_09885_, _10500_, _10498_);
  not _18895_ (_10501_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _18896_ (_10502_, _10485_, _10501_);
  and _18897_ (_10503_, _10485_, word_in[1]);
  or _18898_ (_10504_, _10503_, _10502_);
  and _18899_ (_10505_, _10504_, _10483_);
  and _18900_ (_10506_, _10481_, word_in[9]);
  or _18901_ (_10507_, _10506_, _10505_);
  and _18902_ (_10508_, _10507_, _10478_);
  and _18903_ (_10509_, _10477_, _09194_);
  or _18904_ (_10510_, _10509_, _10495_);
  or _18905_ (_10511_, _10510_, _10508_);
  or _18906_ (_10512_, _10499_, _09075_);
  and _18907_ (_09889_, _10512_, _10511_);
  not _18908_ (_10513_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _18909_ (_10514_, _10485_, _10513_);
  and _18910_ (_10515_, _10485_, word_in[2]);
  or _18911_ (_10516_, _10515_, _10514_);
  and _18912_ (_10517_, _10516_, _10483_);
  and _18913_ (_10518_, _10481_, word_in[10]);
  or _18914_ (_10519_, _10518_, _10517_);
  and _18915_ (_10520_, _10519_, _10478_);
  and _18916_ (_10521_, _10477_, _09217_);
  or _18917_ (_10522_, _10521_, _10495_);
  or _18918_ (_10523_, _10522_, _10520_);
  or _18919_ (_10524_, _10499_, _09634_);
  and _18920_ (_09892_, _10524_, _10523_);
  not _18921_ (_10525_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _18922_ (_10526_, _10485_, _10525_);
  and _18923_ (_10527_, _10485_, word_in[3]);
  or _18924_ (_10528_, _10527_, _10526_);
  and _18925_ (_10529_, _10528_, _10483_);
  and _18926_ (_10530_, _10481_, word_in[11]);
  or _18927_ (_10531_, _10530_, _10529_);
  and _18928_ (_10532_, _10531_, _10478_);
  and _18929_ (_10533_, _10477_, _09113_);
  or _18930_ (_10534_, _10533_, _10495_);
  or _18931_ (_10535_, _10534_, _10532_);
  or _18932_ (_10536_, _10499_, _09103_);
  and _18933_ (_09895_, _10536_, _10535_);
  not _18934_ (_10537_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _18935_ (_10538_, _10485_, _10537_);
  and _18936_ (_10539_, _10485_, word_in[4]);
  or _18937_ (_10540_, _10539_, _10538_);
  and _18938_ (_10541_, _10540_, _10483_);
  and _18939_ (_10542_, _10481_, word_in[12]);
  or _18940_ (_10543_, _10542_, _10541_);
  and _18941_ (_10544_, _10543_, _10478_);
  and _18942_ (_10545_, _10477_, _09287_);
  or _18943_ (_10546_, _10545_, _10495_);
  or _18944_ (_10547_, _10546_, _10544_);
  or _18945_ (_10548_, _10499_, _09659_);
  and _18946_ (_09898_, _10548_, _10547_);
  not _18947_ (_10549_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _18948_ (_10550_, _10485_, _10549_);
  and _18949_ (_10551_, _10485_, word_in[5]);
  or _18950_ (_10552_, _10551_, _10550_);
  and _18951_ (_10553_, _10552_, _10483_);
  and _18952_ (_10554_, _10481_, word_in[13]);
  or _18953_ (_10555_, _10554_, _10553_);
  and _18954_ (_10556_, _10555_, _10478_);
  and _18955_ (_10557_, _10477_, _09305_);
  or _18956_ (_10558_, _10557_, _10495_);
  or _18957_ (_10559_, _10558_, _10556_);
  or _18958_ (_10560_, _10499_, _09140_);
  and _18959_ (_09902_, _10560_, _10559_);
  not _18960_ (_10561_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _18961_ (_10562_, _10485_, _10561_);
  and _18962_ (_10563_, _10485_, word_in[6]);
  or _18963_ (_10564_, _10563_, _10562_);
  and _18964_ (_10565_, _10564_, _10483_);
  and _18965_ (_10566_, _10481_, word_in[14]);
  or _18966_ (_10567_, _10566_, _10565_);
  and _18967_ (_10568_, _10567_, _10478_);
  and _18968_ (_10569_, _10477_, _09322_);
  or _18969_ (_10570_, _10569_, _10495_);
  or _18970_ (_10571_, _10570_, _10568_);
  or _18971_ (_10572_, _10499_, _09684_);
  and _18972_ (_09905_, _10572_, _10571_);
  nor _18973_ (_10573_, _10485_, _08402_);
  and _18974_ (_10574_, _10485_, word_in[7]);
  or _18975_ (_10575_, _10574_, _10573_);
  and _18976_ (_10576_, _10575_, _10483_);
  and _18977_ (_10577_, _10481_, word_in[15]);
  or _18978_ (_10578_, _10577_, _10576_);
  and _18979_ (_10579_, _10578_, _10478_);
  and _18980_ (_10580_, _10477_, _08566_);
  or _18981_ (_10581_, _10580_, _10495_);
  or _18982_ (_10582_, _10581_, _10579_);
  or _18983_ (_10583_, _10499_, _08540_);
  and _18984_ (_09907_, _10583_, _10582_);
  and _18985_ (_10584_, _08547_, _08310_);
  not _18986_ (_10585_, _10584_);
  and _18987_ (_10586_, _09173_, _08350_);
  and _18988_ (_10587_, _09177_, _08556_);
  and _18989_ (_10588_, _10587_, _09056_);
  not _18990_ (_10589_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _18991_ (_10590_, _10587_, _10589_);
  nor _18992_ (_10591_, _10590_, _10588_);
  nor _18993_ (_10592_, _10591_, _10586_);
  and _18994_ (_10593_, _10586_, word_in[8]);
  or _18995_ (_10594_, _10593_, _10592_);
  and _18996_ (_10595_, _10594_, _10585_);
  and _18997_ (_10596_, _10494_, _08344_);
  and _18998_ (_10597_, _10584_, _09168_);
  or _18999_ (_10598_, _10597_, _10596_);
  or _19000_ (_10599_, _10598_, _10595_);
  not _19001_ (_10600_, _10596_);
  or _19002_ (_10601_, _10600_, word_in[24]);
  and _19003_ (_14024_, _10601_, _10599_);
  nor _19004_ (_10602_, _09341_, _08865_);
  and _19005_ (_10603_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _19006_ (_10604_, _10603_, _10602_);
  and _19007_ (_09983_, _10604_, _06071_);
  or _19008_ (_10605_, _10585_, _09194_);
  not _19009_ (_10606_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _19010_ (_10607_, _10587_, _10606_);
  and _19011_ (_10608_, _10587_, _09080_);
  or _19012_ (_10609_, _10608_, _10607_);
  or _19013_ (_10610_, _10609_, _10586_);
  not _19014_ (_10611_, _10586_);
  or _19015_ (_10612_, _10611_, word_in[9]);
  and _19016_ (_10613_, _10612_, _10610_);
  or _19017_ (_10614_, _10613_, _10584_);
  and _19018_ (_10615_, _10614_, _10605_);
  and _19019_ (_10616_, _10615_, _10600_);
  and _19020_ (_10617_, _10596_, word_in[25]);
  or _19021_ (_09985_, _10617_, _10616_);
  or _19022_ (_10618_, _10611_, word_in[10]);
  not _19023_ (_10619_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _19024_ (_10620_, _10587_, _10619_);
  and _19025_ (_10621_, _10587_, _09210_);
  or _19026_ (_10622_, _10621_, _10620_);
  or _19027_ (_10623_, _10622_, _10586_);
  and _19028_ (_10624_, _10623_, _10585_);
  and _19029_ (_10625_, _10624_, _10618_);
  and _19030_ (_10626_, _10584_, _09217_);
  or _19031_ (_10627_, _10626_, _10596_);
  or _19032_ (_10628_, _10627_, _10625_);
  or _19033_ (_10629_, _10600_, word_in[26]);
  and _19034_ (_09989_, _10629_, _10628_);
  and _19035_ (_10630_, _10587_, _09260_);
  not _19036_ (_10631_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _19037_ (_10632_, _10587_, _10631_);
  nor _19038_ (_10633_, _10632_, _10630_);
  nor _19039_ (_10634_, _10633_, _10586_);
  and _19040_ (_10635_, _10586_, word_in[11]);
  or _19041_ (_10636_, _10635_, _10634_);
  and _19042_ (_10637_, _10636_, _10585_);
  and _19043_ (_10638_, _10584_, _09113_);
  or _19044_ (_10639_, _10638_, _10596_);
  or _19045_ (_10640_, _10639_, _10637_);
  or _19046_ (_10641_, _10600_, word_in[27]);
  and _19047_ (_09994_, _10641_, _10640_);
  and _19048_ (_10642_, _10587_, _09277_);
  not _19049_ (_10643_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _19050_ (_10644_, _10587_, _10643_);
  nor _19051_ (_10645_, _10644_, _10642_);
  nor _19052_ (_10646_, _10645_, _10586_);
  and _19053_ (_10647_, _10586_, word_in[12]);
  or _19054_ (_10648_, _10647_, _10646_);
  and _19055_ (_10649_, _10648_, _10585_);
  and _19056_ (_10650_, _10584_, _09287_);
  or _19057_ (_10651_, _10650_, _10596_);
  or _19058_ (_10652_, _10651_, _10649_);
  or _19059_ (_10653_, _10600_, word_in[28]);
  and _19060_ (_09996_, _10653_, _10652_);
  not _19061_ (_10654_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _19062_ (_10655_, _10587_, _10654_);
  and _19063_ (_10656_, _10587_, _09297_);
  or _19064_ (_10657_, _10656_, _10655_);
  or _19065_ (_10658_, _10657_, _10586_);
  or _19066_ (_10659_, _10611_, word_in[13]);
  and _19067_ (_10660_, _10659_, _10658_);
  or _19068_ (_10661_, _10660_, _10584_);
  or _19069_ (_10662_, _10585_, _09305_);
  and _19070_ (_10663_, _10662_, _10661_);
  or _19071_ (_10664_, _10663_, _10596_);
  or _19072_ (_10665_, _10600_, word_in[29]);
  and _19073_ (_10001_, _10665_, _10664_);
  or _19074_ (_10666_, _10585_, _09322_);
  not _19075_ (_10667_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _19076_ (_10668_, _10587_, _10667_);
  and _19077_ (_10669_, _10587_, _09315_);
  or _19078_ (_10670_, _10669_, _10668_);
  or _19079_ (_10671_, _10670_, _10586_);
  nand _19080_ (_10672_, _10586_, _09556_);
  and _19081_ (_10673_, _10672_, _10671_);
  or _19082_ (_10674_, _10673_, _10584_);
  and _19083_ (_10675_, _10674_, _10666_);
  or _19084_ (_10676_, _10675_, _10596_);
  or _19085_ (_10677_, _10600_, word_in[30]);
  and _19086_ (_10005_, _10677_, _10676_);
  and _19087_ (_10678_, _10587_, _08558_);
  nor _19088_ (_10679_, _10587_, _08288_);
  nor _19089_ (_10680_, _10679_, _10678_);
  nor _19090_ (_10681_, _10680_, _10586_);
  and _19091_ (_10682_, _10586_, word_in[15]);
  or _19092_ (_10683_, _10682_, _10681_);
  and _19093_ (_10684_, _10683_, _10585_);
  and _19094_ (_10685_, _10584_, _08566_);
  or _19095_ (_10686_, _10685_, _10596_);
  or _19096_ (_10687_, _10686_, _10684_);
  or _19097_ (_10688_, _10600_, word_in[31]);
  and _19098_ (_10009_, _10688_, _10687_);
  or _19099_ (_10689_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not _19100_ (_10690_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _19101_ (_10691_, _06530_, _10690_);
  and _19102_ (_10692_, _10691_, _06071_);
  and _19103_ (_10032_, _10692_, _10689_);
  and _19104_ (_10693_, _10494_, _08310_);
  not _19105_ (_10694_, _10693_);
  and _19106_ (_10695_, _08547_, _08328_);
  not _19107_ (_10696_, _10695_);
  and _19108_ (_10697_, _09361_, _08350_);
  and _19109_ (_10698_, _09365_, _08532_);
  and _19110_ (_10699_, _10698_, _09056_);
  not _19111_ (_10700_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _19112_ (_10701_, _10698_, _10700_);
  nor _19113_ (_10702_, _10701_, _10699_);
  nor _19114_ (_10703_, _10702_, _10697_);
  and _19115_ (_10704_, _10697_, word_in[8]);
  or _19116_ (_10705_, _10704_, _10703_);
  and _19117_ (_10706_, _10705_, _10696_);
  and _19118_ (_10707_, _10695_, _09168_);
  or _19119_ (_10708_, _10707_, _10706_);
  and _19120_ (_10709_, _10708_, _10694_);
  and _19121_ (_10710_, _10693_, word_in[24]);
  or _19122_ (_10077_, _10710_, _10709_);
  and _19123_ (_10711_, _10698_, _09080_);
  not _19124_ (_10712_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _19125_ (_10713_, _10698_, _10712_);
  nor _19126_ (_10714_, _10713_, _10711_);
  nor _19127_ (_10715_, _10714_, _10697_);
  and _19128_ (_10716_, _10697_, word_in[9]);
  or _19129_ (_10717_, _10716_, _10715_);
  and _19130_ (_10718_, _10717_, _10696_);
  and _19131_ (_10719_, _10695_, _09194_);
  or _19132_ (_10720_, _10719_, _10693_);
  or _19133_ (_10721_, _10720_, _10718_);
  or _19134_ (_10722_, _10694_, word_in[25]);
  and _19135_ (_10081_, _10722_, _10721_);
  and _19136_ (_10723_, _10698_, _09210_);
  not _19137_ (_10724_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _19138_ (_10725_, _10698_, _10724_);
  nor _19139_ (_10726_, _10725_, _10723_);
  nor _19140_ (_10727_, _10726_, _10697_);
  and _19141_ (_10728_, _10697_, word_in[10]);
  or _19142_ (_10729_, _10728_, _10727_);
  and _19143_ (_10730_, _10729_, _10696_);
  and _19144_ (_10731_, _10695_, _09217_);
  or _19145_ (_10732_, _10731_, _10693_);
  or _19146_ (_10733_, _10732_, _10730_);
  or _19147_ (_10734_, _10694_, word_in[26]);
  and _19148_ (_10086_, _10734_, _10733_);
  and _19149_ (_10735_, _10698_, _09260_);
  not _19150_ (_10736_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _19151_ (_10737_, _10698_, _10736_);
  nor _19152_ (_10738_, _10737_, _10735_);
  nor _19153_ (_10739_, _10738_, _10697_);
  and _19154_ (_10740_, _10697_, word_in[11]);
  or _19155_ (_10741_, _10740_, _10739_);
  and _19156_ (_10742_, _10741_, _10696_);
  and _19157_ (_10743_, _10695_, _09113_);
  or _19158_ (_10744_, _10743_, _10693_);
  or _19159_ (_10745_, _10744_, _10742_);
  or _19160_ (_10746_, _10694_, word_in[27]);
  and _19161_ (_10091_, _10746_, _10745_);
  not _19162_ (_10747_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _19163_ (_10748_, _10698_, _10747_);
  and _19164_ (_10749_, _10698_, _09277_);
  or _19165_ (_10750_, _10749_, _10748_);
  or _19166_ (_10751_, _10750_, _10697_);
  not _19167_ (_10752_, _10697_);
  or _19168_ (_10753_, _10752_, word_in[12]);
  and _19169_ (_10754_, _10753_, _10751_);
  or _19170_ (_10755_, _10754_, _10695_);
  or _19171_ (_10756_, _10696_, _09287_);
  and _19172_ (_10757_, _10756_, _10755_);
  or _19173_ (_10758_, _10757_, _10693_);
  or _19174_ (_10759_, _10694_, word_in[28]);
  and _19175_ (_10094_, _10759_, _10758_);
  and _19176_ (_10760_, _10698_, _09297_);
  not _19177_ (_10761_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _19178_ (_10762_, _10698_, _10761_);
  nor _19179_ (_10763_, _10762_, _10760_);
  nor _19180_ (_10764_, _10763_, _10697_);
  and _19181_ (_10765_, _10697_, word_in[13]);
  or _19182_ (_10766_, _10765_, _10764_);
  and _19183_ (_10767_, _10766_, _10696_);
  and _19184_ (_10768_, _10695_, _09305_);
  or _19185_ (_10769_, _10768_, _10693_);
  or _19186_ (_10770_, _10769_, _10767_);
  or _19187_ (_10771_, _10694_, word_in[29]);
  and _19188_ (_10099_, _10771_, _10770_);
  and _19189_ (_10772_, _10698_, _09315_);
  not _19190_ (_10773_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _19191_ (_10774_, _10698_, _10773_);
  nor _19192_ (_10775_, _10774_, _10772_);
  nor _19193_ (_10776_, _10775_, _10697_);
  and _19194_ (_10777_, _10697_, word_in[14]);
  or _19195_ (_10778_, _10777_, _10776_);
  and _19196_ (_10779_, _10778_, _10696_);
  and _19197_ (_10780_, _10695_, _09322_);
  or _19198_ (_10781_, _10780_, _10693_);
  or _19199_ (_10782_, _10781_, _10779_);
  or _19200_ (_10783_, _10694_, word_in[30]);
  and _19201_ (_10104_, _10783_, _10782_);
  and _19202_ (_10784_, _10698_, _08558_);
  nor _19203_ (_10785_, _10698_, _08397_);
  nor _19204_ (_10786_, _10785_, _10784_);
  nor _19205_ (_10787_, _10786_, _10697_);
  and _19206_ (_10788_, _10697_, word_in[15]);
  or _19207_ (_10789_, _10788_, _10787_);
  and _19208_ (_10790_, _10789_, _10696_);
  and _19209_ (_10791_, _10695_, _08566_);
  or _19210_ (_10792_, _10791_, _10693_);
  or _19211_ (_10793_, _10792_, _10790_);
  or _19212_ (_10794_, _10694_, word_in[31]);
  and _19213_ (_10106_, _10794_, _10793_);
  not _19214_ (_10795_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _19215_ (_10796_, _08557_, _10795_);
  and _19216_ (_10797_, _09056_, _08557_);
  or _19217_ (_10798_, _10797_, _10796_);
  or _19218_ (_10799_, _10798_, _08552_);
  not _19219_ (_10800_, _08552_);
  or _19220_ (_10801_, _10800_, word_in[8]);
  and _19221_ (_10802_, _10801_, _10799_);
  or _19222_ (_10803_, _10802_, _08548_);
  or _19223_ (_10804_, _09168_, _08549_);
  and _19224_ (_10805_, _10804_, _08544_);
  and _19225_ (_10806_, _10805_, _10803_);
  and _19226_ (_10807_, _08542_, word_in[24]);
  or _19227_ (_10170_, _10807_, _10806_);
  and _19228_ (_10808_, _08542_, word_in[25]);
  not _19229_ (_10809_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _19230_ (_10810_, _08557_, _10809_);
  and _19231_ (_10811_, _09080_, _08557_);
  or _19232_ (_10812_, _10811_, _10810_);
  or _19233_ (_10813_, _10812_, _08552_);
  or _19234_ (_10814_, _10800_, word_in[9]);
  and _19235_ (_10815_, _10814_, _10813_);
  or _19236_ (_10816_, _10815_, _08548_);
  or _19237_ (_10817_, _09194_, _08549_);
  and _19238_ (_10818_, _10817_, _08544_);
  and _19239_ (_10819_, _10818_, _10816_);
  or _19240_ (_10174_, _10819_, _10808_);
  not _19241_ (_10820_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _19242_ (_10821_, _08557_, _10820_);
  and _19243_ (_10822_, _09210_, _08557_);
  or _19244_ (_10823_, _10822_, _10821_);
  or _19245_ (_10824_, _10823_, _08552_);
  or _19246_ (_10825_, _10800_, word_in[10]);
  and _19247_ (_10826_, _10825_, _10824_);
  or _19248_ (_10827_, _10826_, _08548_);
  or _19249_ (_10828_, _09217_, _08549_);
  and _19250_ (_10829_, _10828_, _08544_);
  and _19251_ (_10830_, _10829_, _10827_);
  and _19252_ (_10831_, _08542_, word_in[26]);
  or _19253_ (_10176_, _10831_, _10830_);
  and _19254_ (_10832_, _07979_, _06360_);
  and _19255_ (_10833_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _19256_ (_10834_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _19257_ (_10835_, _10834_, _07983_);
  or _19258_ (_10836_, _10835_, _10833_);
  or _19259_ (_10837_, _10836_, _10832_);
  and _19260_ (_10178_, _10837_, _06071_);
  not _19261_ (_10838_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _19262_ (_10839_, _08557_, _10838_);
  and _19263_ (_10840_, _09260_, _08557_);
  or _19264_ (_10841_, _10840_, _10839_);
  or _19265_ (_10842_, _10841_, _08552_);
  or _19266_ (_10843_, _10800_, word_in[11]);
  and _19267_ (_10844_, _10843_, _10842_);
  or _19268_ (_10845_, _10844_, _08548_);
  or _19269_ (_10846_, _09113_, _08549_);
  and _19270_ (_10847_, _10846_, _08544_);
  and _19271_ (_10848_, _10847_, _10845_);
  and _19272_ (_10849_, _08542_, word_in[27]);
  or _19273_ (_10180_, _10849_, _10848_);
  not _19274_ (_10850_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _19275_ (_10851_, _08557_, _10850_);
  and _19276_ (_10852_, _09277_, _08557_);
  or _19277_ (_10853_, _10852_, _10851_);
  or _19278_ (_10854_, _10853_, _08552_);
  or _19279_ (_10855_, _10800_, word_in[12]);
  and _19280_ (_10856_, _10855_, _10854_);
  or _19281_ (_10857_, _10856_, _08548_);
  or _19282_ (_10858_, _09287_, _08549_);
  and _19283_ (_10859_, _10858_, _08544_);
  and _19284_ (_10860_, _10859_, _10857_);
  and _19285_ (_10861_, _08542_, word_in[28]);
  or _19286_ (_10184_, _10861_, _10860_);
  not _19287_ (_10862_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _19288_ (_10863_, _08557_, _10862_);
  and _19289_ (_10864_, _09297_, _08557_);
  or _19290_ (_10865_, _10864_, _10863_);
  or _19291_ (_10866_, _10865_, _08552_);
  or _19292_ (_10867_, _10800_, word_in[13]);
  and _19293_ (_10868_, _10867_, _10866_);
  or _19294_ (_10869_, _10868_, _08548_);
  or _19295_ (_10870_, _09305_, _08549_);
  and _19296_ (_10871_, _10870_, _08544_);
  and _19297_ (_10872_, _10871_, _10869_);
  and _19298_ (_10873_, _08542_, word_in[29]);
  or _19299_ (_10187_, _10873_, _10872_);
  not _19300_ (_10874_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _19301_ (_10875_, _08557_, _10874_);
  and _19302_ (_10876_, _09315_, _08557_);
  or _19303_ (_10878_, _10876_, _10875_);
  or _19304_ (_10879_, _10878_, _08552_);
  nand _19305_ (_10880_, _08552_, _09556_);
  and _19306_ (_10881_, _10880_, _10879_);
  or _19307_ (_10882_, _10881_, _08548_);
  or _19308_ (_10883_, _09322_, _08549_);
  and _19309_ (_10884_, _10883_, _08544_);
  and _19310_ (_10885_, _10884_, _10882_);
  and _19311_ (_10886_, _08542_, word_in[30]);
  or _19312_ (_10190_, _10886_, _10885_);
  not _19313_ (_10887_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _19314_ (_10888_, _09028_, _07105_);
  nand _19315_ (_10889_, _10888_, _10887_);
  and _19316_ (_10890_, _10889_, _08989_);
  or _19317_ (_10891_, _10888_, _08799_);
  and _19318_ (_10892_, _10891_, _10890_);
  nor _19319_ (_10893_, _08989_, _07945_);
  or _19320_ (_10894_, _10893_, _10892_);
  and _19321_ (_10419_, _10894_, _06071_);
  and _19322_ (_10895_, _09026_, _06815_);
  and _19323_ (_10896_, _10895_, _06809_);
  not _19324_ (_10897_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _19325_ (_10898_, _08801_, _10897_);
  nand _19326_ (_10899_, _10898_, _10896_);
  or _19327_ (_10900_, _10899_, _08802_);
  nand _19328_ (_10902_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and _19329_ (_10903_, _06735_, _06715_);
  and _19330_ (_10904_, _06706_, _06615_);
  nor _19331_ (_10905_, _10904_, _10903_);
  nor _19332_ (_10906_, _10905_, _10902_);
  or _19333_ (_10907_, _10902_, _06349_);
  and _19334_ (_10908_, _10907_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _19335_ (_10910_, _10908_, _10896_);
  or _19336_ (_10911_, _10910_, _10906_);
  and _19337_ (_10912_, _10911_, _08985_);
  nor _19338_ (_10913_, _09341_, _08985_);
  or _19339_ (_10914_, _10913_, _10912_);
  and _19340_ (_10915_, _10914_, _06071_);
  and _19341_ (_10424_, _10915_, _10900_);
  not _19342_ (_10916_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _19343_ (_10917_, _09028_, _06032_);
  nand _19344_ (_10918_, _10917_, _10916_);
  and _19345_ (_10919_, _10918_, _08989_);
  or _19346_ (_10920_, _10917_, _08799_);
  and _19347_ (_10921_, _10920_, _10919_);
  nor _19348_ (_10922_, _08989_, _06609_);
  or _19349_ (_10923_, _10922_, _10921_);
  and _19350_ (_10427_, _10923_, _06071_);
  and _19351_ (_10924_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _19352_ (_10925_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06071_);
  and _19353_ (_10926_, _10925_, _07011_);
  or _19354_ (_10430_, _10926_, _10924_);
  not _19355_ (_10927_, _06006_);
  nor _19356_ (_10928_, _06803_, _10927_);
  not _19357_ (_10929_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _19358_ (_10930_, _06005_, _05982_);
  nor _19359_ (_10931_, _10930_, _10929_);
  or _19360_ (_10932_, _10931_, _10928_);
  and _19361_ (_10933_, _10896_, _06071_);
  and _19362_ (_10934_, _10933_, _10932_);
  not _19363_ (_10935_, _10896_);
  and _19364_ (_10936_, _10930_, _10927_);
  or _19365_ (_10937_, _10936_, _10935_);
  and _19366_ (_10938_, _10937_, _08157_);
  or _19367_ (_10433_, _10938_, _10934_);
  and _19368_ (_10939_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _19369_ (_10940_, _10939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _19370_ (_10449_, _10940_, _06071_);
  and _19371_ (_10941_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _19372_ (_10942_, _10941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _19373_ (_10459_, _10942_, _06071_);
  and _19374_ (_10943_, _05954_, _07767_);
  and _19375_ (_10944_, _06378_, _05923_);
  not _19376_ (_10945_, _06815_);
  nor _19377_ (_10946_, _10945_, _05967_);
  and _19378_ (_10947_, _10946_, _10944_);
  and _19379_ (_10948_, _10947_, _10943_);
  and _19380_ (_10949_, _10948_, _06805_);
  or _19381_ (_10950_, _10949_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _19382_ (_10951_, _07768_, _06820_);
  and _19383_ (_10952_, _10951_, _09248_);
  not _19384_ (_10953_, _10952_);
  and _19385_ (_10954_, _10953_, _10950_);
  nand _19386_ (_10955_, _10949_, _06803_);
  and _19387_ (_10956_, _10955_, _10954_);
  nor _19388_ (_10957_, _10953_, _06359_);
  or _19389_ (_10958_, _10957_, _10956_);
  and _19390_ (_10480_, _10958_, _06071_);
  and _19391_ (_10959_, _10947_, _06806_);
  nand _19392_ (_10960_, _10959_, _06004_);
  and _19393_ (_10961_, _10960_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _19394_ (_10962_, _10961_, _09249_);
  or _19395_ (_10963_, _07753_, _06005_);
  and _19396_ (_10964_, _10963_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _19397_ (_10965_, _10964_, _08802_);
  and _19398_ (_10966_, _10965_, _10959_);
  or _19399_ (_10967_, _10966_, _10962_);
  nand _19400_ (_10968_, _09341_, _09249_);
  and _19401_ (_10969_, _10968_, _06071_);
  and _19402_ (_10482_, _10969_, _10967_);
  and _19403_ (_10970_, _09584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and _19404_ (_10971_, _09580_, _07891_);
  and _19405_ (_10972_, _09005_, _10971_);
  or _19406_ (_10973_, _10972_, _10970_);
  and _19407_ (_10877_, _10973_, _06071_);
  and _19408_ (_10974_, _07010_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _19409_ (_10976_, _10974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _19410_ (_10901_, _10976_, _06071_);
  nor _19411_ (_10977_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _19412_ (_10978_, _10977_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _19413_ (_10979_, _10978_, _08110_);
  or _19414_ (_10980_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _19415_ (_10981_, _10980_, _06071_);
  and _19416_ (_10909_, _10981_, _10979_);
  not _19417_ (_10982_, _08660_);
  and _19418_ (_10984_, _10982_, _08619_);
  or _19419_ (_10985_, _08018_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _19420_ (_03483_, _10985_, _06071_);
  and _19421_ (_10987_, _03483_, _08021_);
  and _19422_ (_10975_, _10987_, _10984_);
  and _19423_ (_10988_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  not _19424_ (_10989_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor _19425_ (_10990_, _06530_, _10989_);
  or _19426_ (_10992_, _10990_, _10988_);
  and _19427_ (_10983_, _10992_, _06071_);
  and _19428_ (_10994_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  not _19429_ (_10995_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor _19430_ (_10997_, _06530_, _10995_);
  or _19431_ (_10998_, _10997_, _10994_);
  and _19432_ (_10986_, _10998_, _06071_);
  and _19433_ (_11000_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _19434_ (_11001_, _06530_, _09022_);
  or _19435_ (_11002_, _11001_, _11000_);
  and _19436_ (_10991_, _11002_, _06071_);
  and _19437_ (_11003_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not _19438_ (_11005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor _19439_ (_11006_, _06530_, _11005_);
  or _19440_ (_11007_, _11006_, _11003_);
  and _19441_ (_10993_, _11007_, _06071_);
  and _19442_ (_11008_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _19443_ (_11009_, _06530_, _05815_);
  or _19444_ (_11010_, _11009_, _11008_);
  and _19445_ (_10996_, _11010_, _06071_);
  and _19446_ (_11011_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _19447_ (_11012_, _06530_, _05760_);
  or _19448_ (_11013_, _11012_, _11011_);
  and _19449_ (_10999_, _11013_, _06071_);
  and _19450_ (_11014_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _19451_ (_11015_, _06530_, _05865_);
  or _19452_ (_11016_, _11015_, _11014_);
  and _19453_ (_11004_, _11016_, _06071_);
  and _19454_ (_11017_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _19455_ (_11018_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _06071_);
  and _19456_ (_11019_, _11018_, _07011_);
  or _19457_ (_11033_, _11019_, _11017_);
  and _19458_ (_11020_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _19459_ (_11021_, _11020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _19460_ (_11034_, _11021_, _06071_);
  and _19461_ (_11022_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  not _19462_ (_11023_, _09037_);
  and _19463_ (_11024_, _11023_, _06399_);
  and _19464_ (_11025_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _19465_ (_11026_, _11025_, _09345_);
  or _19466_ (_11027_, _11026_, _11024_);
  or _19467_ (_11028_, _11027_, _11022_);
  and _19468_ (_11072_, _11028_, _06071_);
  not _19469_ (_11029_, _10978_);
  or _19470_ (_11030_, _11029_, _07564_);
  or _19471_ (_11031_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _19472_ (_11032_, _11031_, _06071_);
  and _19473_ (_11159_, _11032_, _11030_);
  and _19474_ (_11175_, _07239_, _06071_);
  not _19475_ (_11035_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _19476_ (_11036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _19477_ (_11037_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _19478_ (_11038_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _19479_ (_11039_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _19480_ (_11040_, _11039_, _11037_);
  and _19481_ (_11041_, _11040_, _11038_);
  nor _19482_ (_11042_, _11041_, _11037_);
  nor _19483_ (_11043_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _19484_ (_11044_, _11043_, _11036_);
  not _19485_ (_11045_, _11044_);
  nor _19486_ (_11046_, _11045_, _11042_);
  nor _19487_ (_11047_, _11046_, _11036_);
  not _19488_ (_11048_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _19489_ (_11049_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _19490_ (_11050_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _19491_ (_11051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _19492_ (_11052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _19493_ (_11053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _19494_ (_11054_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _19495_ (_11055_, _11054_, _11053_);
  and _19496_ (_11056_, _11055_, _11052_);
  and _19497_ (_11057_, _11056_, _11051_);
  and _19498_ (_11058_, _11057_, _11050_);
  and _19499_ (_11059_, _11058_, _11049_);
  and _19500_ (_11060_, _11059_, _11048_);
  and _19501_ (_11061_, _11060_, _11047_);
  nor _19502_ (_11062_, _11061_, _11035_);
  and _19503_ (_11063_, _11061_, _11035_);
  nor _19504_ (_11064_, _11063_, _11062_);
  not _19505_ (_11065_, _11064_);
  and _19506_ (_11066_, _11059_, _11047_);
  nor _19507_ (_11067_, _11066_, _11048_);
  nor _19508_ (_11068_, _11067_, _11061_);
  not _19509_ (_11069_, _11068_);
  and _19510_ (_11070_, _11047_, _11058_);
  nor _19511_ (_11071_, _11070_, _11049_);
  or _19512_ (_11073_, _11071_, _11066_);
  not _19513_ (_11074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _19514_ (_11075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _19515_ (_11076_, _11047_, _11057_);
  and _19516_ (_11077_, _11076_, _11075_);
  nor _19517_ (_11078_, _11077_, _11074_);
  or _19518_ (_11079_, _11078_, _11070_);
  and _19519_ (_11080_, _11047_, _11055_);
  and _19520_ (_11081_, _11080_, _11052_);
  nor _19521_ (_11082_, _11081_, _11051_);
  nor _19522_ (_11083_, _11082_, _11076_);
  not _19523_ (_11084_, _11083_);
  nor _19524_ (_11085_, _11080_, _11052_);
  nor _19525_ (_11086_, _11085_, _11081_);
  not _19526_ (_11087_, _11086_);
  and _19527_ (_11088_, _11047_, _11054_);
  nor _19528_ (_11089_, _11088_, _11053_);
  nor _19529_ (_11090_, _11089_, _11080_);
  not _19530_ (_11091_, _11090_);
  nor _19531_ (_11092_, _11047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _19532_ (_11093_, _11047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _19533_ (_11094_, _11093_, _11092_);
  not _19534_ (_11095_, _11094_);
  and _19535_ (_11096_, _05769_, _05726_);
  and _19536_ (_11097_, _11096_, _05880_);
  and _19537_ (_11098_, _11097_, _05861_);
  not _19538_ (_11099_, _11098_);
  nor _19539_ (_11100_, _05810_, _05788_);
  and _19540_ (_11101_, _11100_, _05848_);
  and _19541_ (_11102_, _11101_, _05854_);
  nor _19542_ (_11103_, _05880_, _05726_);
  and _19543_ (_11104_, _05880_, _05726_);
  nor _19544_ (_11105_, _11104_, _11103_);
  and _19545_ (_11106_, _11105_, _11102_);
  and _19546_ (_11107_, _05860_, _05788_);
  and _19547_ (_11108_, _05768_, _05747_);
  and _19548_ (_11109_, _11108_, _05727_);
  and _19549_ (_11110_, _11109_, _05880_);
  and _19550_ (_11111_, _11110_, _11107_);
  nor _19551_ (_11112_, _11111_, _11106_);
  and _19552_ (_11113_, _11112_, _11099_);
  nor _19553_ (_11114_, _05860_, _05853_);
  nor _19554_ (_11115_, _05768_, _05748_);
  and _19555_ (_11116_, _11115_, _11103_);
  and _19556_ (_11117_, _11108_, _05726_);
  and _19557_ (_11118_, _11117_, _05880_);
  and _19558_ (_11119_, _11107_, _11118_);
  nor _19559_ (_11120_, _11119_, _11116_);
  nor _19560_ (_11121_, _11120_, _11114_);
  and _19561_ (_11122_, _11103_, _05769_);
  and _19562_ (_11123_, _11101_, _11122_);
  and _19563_ (_11124_, _11110_, _05847_);
  or _19564_ (_11125_, _11124_, _11123_);
  nor _19565_ (_11126_, _05880_, _05727_);
  and _19566_ (_11127_, _11108_, _11126_);
  and _19567_ (_11128_, _11107_, _11127_);
  and _19568_ (_11129_, _05853_, _11122_);
  or _19569_ (_11130_, _11129_, _11128_);
  or _19570_ (_11131_, _11130_, _11125_);
  nor _19571_ (_11132_, _11131_, _11121_);
  nand _19572_ (_11133_, _11132_, _11113_);
  and _19573_ (_11134_, _11102_, _11104_);
  and _19574_ (_11135_, _11116_, _11101_);
  nor _19575_ (_11136_, _11135_, _11134_);
  and _19576_ (_11137_, _11126_, _05769_);
  and _19577_ (_11138_, _11115_, _05726_);
  and _19578_ (_11139_, _11138_, _05880_);
  nor _19579_ (_11140_, _11139_, _11137_);
  nor _19580_ (_11141_, _11140_, _05857_);
  and _19581_ (_11142_, _05880_, _05727_);
  and _19582_ (_11143_, _11142_, _05769_);
  or _19583_ (_11144_, _11139_, _11143_);
  and _19584_ (_11145_, _11144_, _05861_);
  nor _19585_ (_11146_, _11145_, _11141_);
  and _19586_ (_11147_, _05861_, _05855_);
  and _19587_ (_11148_, _11107_, _05854_);
  nor _19588_ (_11149_, _11148_, _11147_);
  and _19589_ (_11150_, _11149_, _11146_);
  and _19590_ (_11151_, _11115_, _11126_);
  nor _19591_ (_11152_, _05860_, _05849_);
  not _19592_ (_11153_, _11152_);
  and _19593_ (_11154_, _11153_, _11151_);
  not _19594_ (_11155_, _05853_);
  nor _19595_ (_11156_, _11110_, _11139_);
  nor _19596_ (_11157_, _11156_, _11155_);
  nor _19597_ (_11158_, _11157_, _11154_);
  not _19598_ (_11160_, _11107_);
  and _19599_ (_11161_, _11108_, _11103_);
  nor _19600_ (_11162_, _11161_, _11143_);
  nor _19601_ (_11163_, _11162_, _11160_);
  nor _19602_ (_11164_, _11161_, _11097_);
  nor _19603_ (_11165_, _11164_, _11155_);
  nor _19604_ (_11166_, _11165_, _11163_);
  and _19605_ (_11167_, _11166_, _11158_);
  and _19606_ (_11168_, _11167_, _11150_);
  nand _19607_ (_11169_, _11168_, _11136_);
  and _19608_ (_11170_, _11097_, _11107_);
  and _19609_ (_11171_, _11115_, _11142_);
  and _19610_ (_11172_, _11171_, _05850_);
  nor _19611_ (_11173_, _11172_, _11170_);
  nor _19612_ (_11174_, _11139_, _11122_);
  nor _19613_ (_11176_, _11174_, _11160_);
  and _19614_ (_11177_, _05854_, _05727_);
  and _19615_ (_11178_, _11177_, _05853_);
  nor _19616_ (_11179_, _11178_, _11176_);
  nand _19617_ (_11180_, _11179_, _11173_);
  not _19618_ (_11182_, _11171_);
  nor _19619_ (_11183_, _11114_, _11182_);
  and _19620_ (_11185_, _11116_, _05850_);
  and _19621_ (_11186_, _11101_, _11143_);
  nor _19622_ (_11187_, _11186_, _11185_);
  not _19623_ (_11189_, _11187_);
  or _19624_ (_11190_, _11189_, _11183_);
  or _19625_ (_11191_, _11190_, _11180_);
  and _19626_ (_11192_, _05880_, _05857_);
  and _19627_ (_11193_, _05829_, _05810_);
  and _19628_ (_11194_, _11193_, _11192_);
  or _19629_ (_11195_, _11194_, _11101_);
  and _19630_ (_11196_, _11195_, _11138_);
  and _19631_ (_11197_, _11194_, _11096_);
  nand _19632_ (_11198_, _05847_, _05769_);
  nor _19633_ (_11199_, _11198_, _11105_);
  or _19634_ (_11200_, _11199_, _11197_);
  and _19635_ (_11201_, _05858_, _05788_);
  and _19636_ (_11202_, _11201_, _05848_);
  and _19637_ (_11203_, _05882_, _05857_);
  and _19638_ (_11204_, _11203_, _11193_);
  or _19639_ (_11206_, _11204_, _11202_);
  or _19640_ (_11207_, _11206_, _11200_);
  or _19641_ (_11208_, _11207_, _11196_);
  and _19642_ (_11209_, _05853_, _05769_);
  and _19643_ (_11210_, _11209_, _11105_);
  or _19644_ (_11211_, _11109_, _11171_);
  or _19645_ (_11212_, _11211_, _11097_);
  or _19646_ (_11213_, _11212_, _11137_);
  and _19647_ (_11214_, _11213_, _11101_);
  or _19648_ (_11215_, _11214_, _11210_);
  or _19649_ (_11216_, _11215_, _11208_);
  or _19650_ (_11217_, _11216_, _11191_);
  or _19651_ (_11218_, _11217_, _11169_);
  nor _19652_ (_11219_, _11218_, _11133_);
  nor _19653_ (_11221_, _11040_, _11038_);
  nor _19654_ (_11222_, _11221_, _11041_);
  not _19655_ (_11224_, _11222_);
  nor _19656_ (_11225_, _11224_, _11219_);
  and _19657_ (_11226_, _11151_, _05850_);
  nor _19658_ (_11227_, _11226_, _11134_);
  and _19659_ (_11228_, _11227_, _11187_);
  and _19660_ (_11229_, _11228_, _11113_);
  and _19661_ (_11230_, _11097_, _05847_);
  nor _19662_ (_11231_, _11230_, _11197_);
  and _19663_ (_11232_, _11231_, _11173_);
  and _19664_ (_11233_, _11232_, _11179_);
  and _19665_ (_11234_, _11233_, _11229_);
  not _19666_ (_11235_, _11234_);
  nor _19667_ (_11236_, _11235_, _11219_);
  not _19668_ (_11237_, _11236_);
  nor _19669_ (_11238_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _19670_ (_11239_, _11238_, _11038_);
  and _19671_ (_11240_, _11239_, _11237_);
  and _19672_ (_11241_, _11224_, _11219_);
  nor _19673_ (_11242_, _11241_, _11225_);
  and _19674_ (_11243_, _11242_, _11240_);
  nor _19675_ (_11244_, _11243_, _11225_);
  not _19676_ (_11245_, _11244_);
  and _19677_ (_11246_, _11045_, _11042_);
  nor _19678_ (_11247_, _11246_, _11046_);
  and _19679_ (_11248_, _11247_, _11245_);
  and _19680_ (_11249_, _11248_, _11095_);
  and _19681_ (_11250_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _19682_ (_11251_, _11250_, _11054_);
  nand _19683_ (_11252_, _11251_, _11092_);
  or _19684_ (_11253_, _11251_, _11092_);
  and _19685_ (_11254_, _11253_, _11252_);
  and _19686_ (_11255_, _11254_, _11249_);
  and _19687_ (_11256_, _11255_, _11091_);
  and _19688_ (_11257_, _11256_, _11087_);
  and _19689_ (_11258_, _11257_, _11084_);
  nor _19690_ (_11259_, _11076_, _11075_);
  or _19691_ (_11260_, _11259_, _11077_);
  and _19692_ (_11261_, _11260_, _11258_);
  and _19693_ (_11262_, _11261_, _11079_);
  and _19694_ (_11263_, _11262_, _11073_);
  and _19695_ (_11264_, _11263_, _11069_);
  and _19696_ (_11265_, _11264_, _11065_);
  nor _19697_ (_11266_, _11264_, _11065_);
  nor _19698_ (_11267_, _11266_, _11265_);
  or _19699_ (_11268_, _11267_, _09711_);
  or _19700_ (_11269_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _19701_ (_11270_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _19702_ (_11271_, _11270_, _11269_);
  and _19703_ (_11272_, _11271_, _11268_);
  and _19704_ (_11273_, _06071_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _19705_ (_11274_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _19706_ (_11181_, _11274_, _11272_);
  and _19707_ (_11275_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not _19708_ (_11276_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor _19709_ (_11277_, _06530_, _11276_);
  or _19710_ (_11278_, _11277_, _11275_);
  and _19711_ (_11184_, _11278_, _06071_);
  and _19712_ (_11279_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _19713_ (_11280_, _06530_, _09701_);
  or _19714_ (_11281_, _11280_, _11279_);
  and _19715_ (_11188_, _11281_, _06071_);
  and _19716_ (_11282_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _19717_ (_11283_, _06530_, _05833_);
  or _19718_ (_11284_, _11283_, _11282_);
  and _19719_ (_11205_, _11284_, _06071_);
  not _19720_ (_11286_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _19721_ (_11287_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _19722_ (_11288_, _11063_, _11287_);
  nor _19723_ (_11289_, _11288_, _11286_);
  and _19724_ (_11290_, _11288_, _11286_);
  nor _19725_ (_11292_, _11290_, _11289_);
  not _19726_ (_11293_, _11292_);
  nor _19727_ (_11294_, _11063_, _11287_);
  or _19728_ (_11295_, _11294_, _11288_);
  and _19729_ (_11296_, _11295_, _11265_);
  and _19730_ (_11297_, _11296_, _11293_);
  nor _19731_ (_11298_, _11296_, _11293_);
  nor _19732_ (_11299_, _11298_, _11297_);
  or _19733_ (_11300_, _11299_, _09711_);
  or _19734_ (_11301_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _19735_ (_11302_, _11301_, _11270_);
  and _19736_ (_11304_, _11302_, _11300_);
  and _19737_ (_11305_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _19738_ (_11220_, _11305_, _11304_);
  nor _19739_ (_11307_, _11295_, _11265_);
  nor _19740_ (_11308_, _11307_, _11296_);
  or _19741_ (_11309_, _11308_, _09711_);
  or _19742_ (_11310_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _19743_ (_11311_, _11310_, _11270_);
  and _19744_ (_11312_, _11311_, _11309_);
  and _19745_ (_11313_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _19746_ (_11223_, _11313_, _11312_);
  or _19747_ (_11314_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _19748_ (_11315_, _06530_, _05737_);
  and _19749_ (_11316_, _11315_, _06071_);
  and _19750_ (_11285_, _11316_, _11314_);
  nor _19751_ (_11317_, _11263_, _11069_);
  nor _19752_ (_11318_, _11317_, _11264_);
  or _19753_ (_11319_, _11318_, _09711_);
  or _19754_ (_11320_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _19755_ (_11321_, _11320_, _11270_);
  and _19756_ (_11322_, _11321_, _11319_);
  and _19757_ (_11323_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _19758_ (_11291_, _11323_, _11322_);
  and _19759_ (_11324_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _19760_ (_11325_, _06530_, _06958_);
  or _19761_ (_11326_, _11325_, _11324_);
  and _19762_ (_11303_, _11326_, _06071_);
  and _19763_ (_11327_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _19764_ (_11328_, _06530_, _05862_);
  or _19765_ (_11329_, _11328_, _11327_);
  and _19766_ (_11306_, _11329_, _06071_);
  and _19767_ (_11330_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _19768_ (_11331_, _06530_, _05693_);
  or _19769_ (_11332_, _11331_, _11330_);
  and _19770_ (_11339_, _11332_, _06071_);
  nor _19771_ (_11333_, _06527_, _06231_);
  or _19772_ (_11334_, _05811_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor _19773_ (_11335_, _05718_, _10690_);
  nor _19774_ (_11336_, _05696_, _10989_);
  or _19775_ (_11337_, _11336_, _11335_);
  and _19776_ (_11338_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _19777_ (_11340_, _05711_, _05817_);
  nor _19778_ (_11341_, _05705_, _05815_);
  or _19779_ (_11342_, _11341_, _11340_);
  or _19780_ (_11343_, _11342_, _11338_);
  or _19781_ (_11344_, _11343_, _11337_);
  and _19782_ (_11345_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _19783_ (_11346_, _11345_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _19784_ (_11347_, _11346_, _11344_);
  and _19785_ (_11348_, _11347_, _06527_);
  and _19786_ (_11349_, _11348_, _11334_);
  nor _19787_ (_11350_, _11349_, _11333_);
  nor _19788_ (_11373_, _11350_, rst);
  nor _19789_ (_11351_, _06527_, _06224_);
  nor _19790_ (_11352_, _05705_, _05789_);
  nor _19791_ (_11353_, _05711_, _05791_);
  nor _19792_ (_11354_, _11353_, _11352_);
  and _19793_ (_11355_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _19794_ (_11356_, _05700_, _05793_);
  nor _19795_ (_11357_, _11356_, _11355_);
  and _19796_ (_11358_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _19797_ (_11359_, _05718_);
  and _19798_ (_11360_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _19799_ (_11361_, _11360_, _11358_);
  and _19800_ (_11362_, _11361_, _11357_);
  and _19801_ (_11363_, _11362_, _11354_);
  nor _19802_ (_11364_, _11363_, _09711_);
  nor _19803_ (_11365_, _11364_, _11351_);
  nor _19804_ (_11389_, _11365_, rst);
  nor _19805_ (_11366_, _11236_, _05709_);
  nor _19806_ (_11367_, _11219_, _05698_);
  and _19807_ (_11368_, _11219_, _05698_);
  nor _19808_ (_11369_, _11368_, _11367_);
  and _19809_ (_11370_, _11369_, _11366_);
  nor _19810_ (_11371_, _11369_, _11366_);
  nor _19811_ (_11372_, _11371_, _11370_);
  or _19812_ (_11374_, _11372_, _06528_);
  or _19813_ (_11375_, _06527_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _19814_ (_11376_, _11375_, _11270_);
  and _19815_ (_11393_, _11376_, _11374_);
  and _19816_ (_11377_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _19817_ (_11378_, _11262_, _11073_);
  nor _19818_ (_11379_, _11378_, _11263_);
  or _19819_ (_11380_, _11379_, _09711_);
  or _19820_ (_11381_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _19821_ (_11382_, _11381_, _11270_);
  and _19822_ (_11383_, _11382_, _11380_);
  or _19823_ (_11402_, _11383_, _11377_);
  and _19824_ (_11384_, \oc8051_top_1.oc8051_decoder1.state [1], _05686_);
  and _19825_ (_11385_, _11384_, _05685_);
  and _19826_ (_11386_, _08740_, _08737_);
  nor _19827_ (_11387_, _08746_, _11386_);
  and _19828_ (_11388_, _11387_, _08736_);
  and _19829_ (_11390_, _08714_, _08712_);
  and _19830_ (_11391_, _08732_, _11390_);
  and _19831_ (_11392_, _08710_, _08707_);
  and _19832_ (_11394_, _08715_, _11392_);
  and _19833_ (_11395_, _11394_, _08725_);
  and _19834_ (_11396_, _11395_, _08732_);
  or _19835_ (_11397_, _11396_, _11391_);
  nand _19836_ (_11398_, _11397_, _11388_);
  not _19837_ (_11399_, _08736_);
  and _19838_ (_11400_, _08758_, _11399_);
  and _19839_ (_11401_, _11400_, _08732_);
  and _19840_ (_11403_, _11401_, _08728_);
  and _19841_ (_11404_, _11387_, _11399_);
  and _19842_ (_11405_, _11404_, _08728_);
  nor _19843_ (_11406_, _11405_, _11403_);
  and _19844_ (_11407_, _08746_, _11386_);
  and _19845_ (_11408_, _11407_, _08736_);
  and _19846_ (_11410_, _11408_, _08732_);
  and _19847_ (_11411_, _08726_, _08753_);
  and _19848_ (_11412_, _11411_, _11394_);
  and _19849_ (_11413_, _11412_, _11410_);
  and _19850_ (_11414_, _11388_, _08732_);
  and _19851_ (_11415_, _11394_, _08726_);
  and _19852_ (_11416_, _11415_, _11414_);
  nor _19853_ (_11417_, _11416_, _11413_);
  and _19854_ (_11418_, _11417_, _11406_);
  nand _19855_ (_11419_, _11418_, _11398_);
  nand _19856_ (_11420_, _11419_, _11385_);
  or _19857_ (_11421_, _06526_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19858_ (_11422_, _08756_, _08721_);
  and _19859_ (_11423_, _11422_, _11400_);
  and _19860_ (_11424_, _11423_, _11421_);
  not _19861_ (_11425_, _11424_);
  and _19862_ (_11426_, _11384_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19863_ (_11427_, _11422_, _11404_);
  nand _19864_ (_11428_, _11427_, _11426_);
  nand _19865_ (_11429_, _11421_, _11405_);
  and _19866_ (_11430_, _11429_, _11428_);
  and _19867_ (_11431_, _11430_, _11425_);
  nand _19868_ (_11433_, _11431_, _11420_);
  nor _19869_ (_11434_, _06527_, _06080_);
  and _19870_ (_11435_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _19871_ (_11436_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor _19872_ (_11438_, _05700_, _05754_);
  nor _19873_ (_11439_, _11438_, _11436_);
  nor _19874_ (_11441_, _05705_, _05749_);
  and _19875_ (_11442_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _19876_ (_11444_, _11442_, _11441_);
  nor _19877_ (_11445_, _05718_, _10995_);
  nor _19878_ (_11446_, _05711_, _05760_);
  nor _19879_ (_11447_, _11446_, _11445_);
  and _19880_ (_11448_, _11447_, _11444_);
  and _19881_ (_11449_, _11448_, _11439_);
  nor _19882_ (_11450_, _11449_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19883_ (_11451_, _11450_, _11435_);
  nor _19884_ (_11452_, _11451_, _06528_);
  nor _19885_ (_11453_, _11452_, _11434_);
  and _19886_ (_11454_, _11453_, _11433_);
  and _19887_ (_11455_, _11431_, _11420_);
  nor _19888_ (_11456_, _06527_, _06075_);
  nor _19889_ (_11457_, _05705_, _05760_);
  nor _19890_ (_11458_, _05711_, _05754_);
  nor _19891_ (_11459_, _11458_, _11457_);
  nor _19892_ (_11460_, _05696_, _10995_);
  nor _19893_ (_11461_, _05700_, _05756_);
  nor _19894_ (_11462_, _11461_, _11460_);
  and _19895_ (_11463_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _19896_ (_11464_, _05718_, _05749_);
  nor _19897_ (_11465_, _11464_, _11463_);
  and _19898_ (_11466_, _11465_, _11462_);
  and _19899_ (_11467_, _11466_, _11459_);
  nor _19900_ (_11468_, _11467_, _09711_);
  nor _19901_ (_11469_, _11468_, _11456_);
  and _19902_ (_11470_, _11469_, _11455_);
  nor _19903_ (_11471_, _11470_, _11454_);
  not _19904_ (_11472_, _11471_);
  and _19905_ (_11473_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _19906_ (_11474_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _19907_ (_11475_, _11474_);
  nor _19908_ (_11476_, _06527_, _06258_);
  and _19909_ (_11477_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19910_ (_11478_, _05696_, _06850_);
  and _19911_ (_11479_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _19912_ (_11480_, _11479_, _11478_);
  nor _19913_ (_11481_, _05705_, _05737_);
  and _19914_ (_11482_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _19915_ (_11483_, _11482_, _11481_);
  and _19916_ (_11484_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _19917_ (_11485_, _05711_, _05739_);
  nor _19918_ (_11486_, _11485_, _11484_);
  and _19919_ (_11487_, _11486_, _11483_);
  and _19920_ (_11488_, _11487_, _11480_);
  nor _19921_ (_11490_, _11488_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19922_ (_11491_, _11490_, _11477_);
  nor _19923_ (_11492_, _11491_, _06528_);
  nor _19924_ (_11493_, _11492_, _11476_);
  and _19925_ (_11495_, _11493_, _11433_);
  nor _19926_ (_11496_, _06527_, _06256_);
  nor _19927_ (_11497_, _05705_, _05739_);
  and _19928_ (_11498_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _19929_ (_11500_, _11498_, _11497_);
  and _19930_ (_11501_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor _19931_ (_11503_, _05700_, _05732_);
  nor _19932_ (_11504_, _11503_, _11501_);
  and _19933_ (_11505_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _19934_ (_11506_, _05718_, _05737_);
  nor _19935_ (_11507_, _11506_, _11505_);
  and _19936_ (_11508_, _11507_, _11504_);
  and _19937_ (_11509_, _11508_, _11500_);
  nor _19938_ (_11510_, _11509_, _09711_);
  nor _19939_ (_11511_, _11510_, _11496_);
  and _19940_ (_11512_, _11511_, _11455_);
  nor _19941_ (_11513_, _11512_, _11495_);
  nand _19942_ (_11514_, _11513_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _19943_ (_11515_, _11513_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _19944_ (_11516_, _11515_, _11514_);
  nor _19945_ (_11517_, _06527_, _06277_);
  and _19946_ (_11518_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19947_ (_11519_, _05696_, _06532_);
  and _19948_ (_11520_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _19949_ (_11521_, _11520_, _11519_);
  nor _19950_ (_11522_, _05705_, _05693_);
  and _19951_ (_11523_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _19952_ (_11524_, _11523_, _11522_);
  and _19953_ (_11525_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _19954_ (_11526_, _05711_, _05716_);
  nor _19955_ (_11527_, _11526_, _11525_);
  and _19956_ (_11528_, _11527_, _11524_);
  and _19957_ (_11529_, _11528_, _11521_);
  nor _19958_ (_11530_, _11529_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19959_ (_11531_, _11530_, _11518_);
  nor _19960_ (_11532_, _11531_, _06528_);
  nor _19961_ (_11533_, _11532_, _11517_);
  and _19962_ (_11534_, _11533_, _11433_);
  nor _19963_ (_11535_, _06527_, _06279_);
  nor _19964_ (_11536_, _05705_, _05716_);
  and _19965_ (_11537_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _19966_ (_11538_, _11537_, _11536_);
  and _19967_ (_11539_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _19968_ (_11540_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _19969_ (_11541_, _11540_, _11539_);
  nor _19970_ (_11542_, _05718_, _05693_);
  nor _19971_ (_11543_, _05700_, _05708_);
  nor _19972_ (_11545_, _11543_, _11542_);
  and _19973_ (_11546_, _11545_, _11541_);
  and _19974_ (_11547_, _11546_, _11538_);
  nor _19975_ (_11548_, _11547_, _09711_);
  nor _19976_ (_11549_, _11548_, _11535_);
  and _19977_ (_11550_, _11549_, _11455_);
  nor _19978_ (_11551_, _11550_, _11534_);
  nor _19979_ (_11552_, _11551_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _19980_ (_11553_, _11551_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _19981_ (_11554_, _06527_, _06148_);
  or _19982_ (_11555_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05811_);
  nor _19983_ (_11556_, _05718_, _09701_);
  nor _19984_ (_11557_, _05696_, _06958_);
  or _19985_ (_11558_, _11557_, _11556_);
  and _19986_ (_11559_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _19987_ (_11560_, _05705_, _05862_);
  nor _19988_ (_11561_, _05711_, _05865_);
  or _19989_ (_11562_, _11561_, _11560_);
  or _19990_ (_11563_, _11562_, _11559_);
  or _19991_ (_11564_, _11563_, _11558_);
  and _19992_ (_11565_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _19993_ (_11566_, _11565_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _19994_ (_11567_, _11566_, _11564_);
  and _19995_ (_11568_, _11567_, _06527_);
  and _19996_ (_11569_, _11568_, _11555_);
  nor _19997_ (_11570_, _11569_, _11554_);
  and _19998_ (_11571_, _11570_, _11433_);
  and _19999_ (_11572_, _11455_, _09713_);
  nor _20000_ (_11573_, _11572_, _11571_);
  nand _20001_ (_11574_, _11573_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _20002_ (_11575_, _06527_, _06167_);
  and _20003_ (_11576_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20004_ (_11577_, _05696_, _11276_);
  and _20005_ (_11578_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _20006_ (_11579_, _11578_, _11577_);
  nor _20007_ (_11580_, _05705_, _05833_);
  and _20008_ (_11581_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _20009_ (_11582_, _11581_, _11580_);
  nor _20010_ (_11583_, _05718_, _09022_);
  nor _20011_ (_11584_, _05711_, _05835_);
  nor _20012_ (_11585_, _11584_, _11583_);
  and _20013_ (_11586_, _11585_, _11582_);
  and _20014_ (_11587_, _11586_, _11579_);
  nor _20015_ (_11588_, _11587_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20016_ (_11589_, _11588_, _11576_);
  nor _20017_ (_11590_, _11589_, _06528_);
  nor _20018_ (_11591_, _11590_, _11575_);
  and _20019_ (_11592_, _11591_, _11433_);
  nor _20020_ (_11593_, _06527_, _06169_);
  nor _20021_ (_11594_, _05705_, _05835_);
  and _20022_ (_11595_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _20023_ (_11596_, _11595_, _11594_);
  nor _20024_ (_11597_, _05696_, _09022_);
  and _20025_ (_11598_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _20026_ (_11600_, _11598_, _11597_);
  nor _20027_ (_11601_, _05718_, _05833_);
  and _20028_ (_11602_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _20029_ (_11603_, _11602_, _11601_);
  and _20030_ (_11604_, _11603_, _11600_);
  and _20031_ (_11605_, _11604_, _11596_);
  nor _20032_ (_11606_, _11605_, _09711_);
  nor _20033_ (_11607_, _11606_, _11593_);
  and _20034_ (_11608_, _11607_, _11455_);
  nor _20035_ (_11609_, _11608_, _11592_);
  nor _20036_ (_11610_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20037_ (_11611_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _20038_ (_11612_, _11350_);
  or _20039_ (_11613_, _11455_, _11612_);
  nor _20040_ (_11614_, _06527_, _06233_);
  nor _20041_ (_11615_, _05705_, _05817_);
  and _20042_ (_11616_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _20043_ (_11617_, _11616_, _11615_);
  nor _20044_ (_11618_, _05696_, _10690_);
  and _20045_ (_11619_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _20046_ (_11620_, _11619_, _11618_);
  and _20047_ (_11621_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _20048_ (_11622_, _05718_, _05815_);
  nor _20049_ (_11623_, _11622_, _11621_);
  and _20050_ (_11624_, _11623_, _11620_);
  and _20051_ (_11625_, _11624_, _11617_);
  nor _20052_ (_11626_, _11625_, _09711_);
  nor _20053_ (_11627_, _11626_, _11614_);
  not _20054_ (_11628_, _11627_);
  or _20055_ (_11629_, _11628_, _11433_);
  nand _20056_ (_11630_, _11629_, _11613_);
  or _20057_ (_11631_, _11630_, _06241_);
  nor _20058_ (_11632_, _06527_, _06214_);
  and _20059_ (_11633_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20060_ (_11634_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor _20061_ (_11635_, _05700_, _05791_);
  nor _20062_ (_11636_, _11635_, _11634_);
  and _20063_ (_11637_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _20064_ (_11638_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _20065_ (_11639_, _11638_, _11637_);
  and _20066_ (_11640_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor _20067_ (_11641_, _05711_, _05789_);
  nor _20068_ (_11642_, _11641_, _11640_);
  and _20069_ (_11643_, _11642_, _11639_);
  and _20070_ (_11644_, _11643_, _11636_);
  nor _20071_ (_11645_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20072_ (_11646_, _11645_, _11633_);
  nor _20073_ (_11647_, _11646_, _06528_);
  nor _20074_ (_11648_, _11647_, _11632_);
  not _20075_ (_11649_, _11648_);
  or _20076_ (_11650_, _11649_, _11455_);
  not _20077_ (_11651_, _11365_);
  or _20078_ (_11652_, _11433_, _11651_);
  and _20079_ (_11653_, _11652_, _11650_);
  nand _20080_ (_11654_, _11653_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _20081_ (_11655_, _06527_, _06190_);
  and _20082_ (_11656_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20083_ (_11657_, _05696_, _06962_);
  and _20084_ (_11658_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20085_ (_11659_, _11658_, _11657_);
  nor _20086_ (_11660_, _05705_, _05782_);
  and _20087_ (_11661_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20088_ (_11662_, _11661_, _11660_);
  nor _20089_ (_11663_, _05718_, _11005_);
  nor _20090_ (_11664_, _05711_, _05773_);
  nor _20091_ (_11665_, _11664_, _11663_);
  and _20092_ (_11666_, _11665_, _11662_);
  and _20093_ (_11667_, _11666_, _11659_);
  nor _20094_ (_11668_, _11667_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20095_ (_11669_, _11668_, _11656_);
  nor _20096_ (_11670_, _11669_, _06528_);
  nor _20097_ (_11671_, _11670_, _11655_);
  not _20098_ (_11672_, _11671_);
  or _20099_ (_11673_, _11672_, _11455_);
  nor _20100_ (_11674_, _06527_, _06188_);
  nor _20101_ (_11675_, _05705_, _05773_);
  and _20102_ (_11676_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20103_ (_11678_, _11676_, _11675_);
  nor _20104_ (_11679_, _05696_, _11005_);
  and _20105_ (_11680_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20106_ (_11681_, _11680_, _11679_);
  and _20107_ (_11682_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _20108_ (_11683_, _05718_, _05782_);
  nor _20109_ (_11684_, _11683_, _11682_);
  and _20110_ (_11685_, _11684_, _11681_);
  and _20111_ (_11686_, _11685_, _11678_);
  nor _20112_ (_11687_, _11686_, _09711_);
  nor _20113_ (_11688_, _11687_, _11674_);
  not _20114_ (_11689_, _11688_);
  or _20115_ (_11690_, _11689_, _11433_);
  and _20116_ (_11691_, _11690_, _11673_);
  and _20117_ (_11693_, _11691_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _20118_ (_11694_, _11653_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20119_ (_11695_, _11694_, _11654_);
  and _20120_ (_11696_, _11695_, _11693_);
  not _20121_ (_11697_, _11696_);
  nand _20122_ (_11698_, _11697_, _11654_);
  nand _20123_ (_11699_, _11630_, _06241_);
  and _20124_ (_11700_, _11699_, _11631_);
  and _20125_ (_11701_, _11700_, _11698_);
  not _20126_ (_11702_, _11701_);
  nand _20127_ (_11703_, _11702_, _11631_);
  nor _20128_ (_11704_, _11703_, _11611_);
  nor _20129_ (_11705_, _11704_, _11610_);
  or _20130_ (_11706_, _11573_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20131_ (_11707_, _11706_, _11574_);
  nand _20132_ (_11708_, _11707_, _11705_);
  nand _20133_ (_11709_, _11708_, _11574_);
  nor _20134_ (_11710_, _11709_, _11553_);
  nor _20135_ (_11711_, _11710_, _11552_);
  nand _20136_ (_11713_, _11711_, _11516_);
  nand _20137_ (_11714_, _11713_, _11514_);
  and _20138_ (_11715_, _11714_, _11475_);
  or _20139_ (_11716_, _11715_, _11473_);
  or _20140_ (_11717_, _11716_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _20141_ (_11718_, _11717_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _20142_ (_11719_, _11718_, _06243_);
  or _20143_ (_11721_, _11719_, _11472_);
  and _20144_ (_11722_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _20145_ (_11723_, _11722_, _11716_);
  and _20146_ (_11724_, _11723_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand _20147_ (_11725_, _11724_, _11472_);
  and _20148_ (_11726_, _11725_, _11721_);
  nand _20149_ (_11727_, _11726_, _06172_);
  or _20150_ (_11728_, _11726_, _06172_);
  and _20151_ (_11729_, _11429_, _11420_);
  not _20152_ (_11730_, _11385_);
  nor _20153_ (_11731_, _08741_, _08736_);
  and _20154_ (_11732_, _11731_, _08728_);
  and _20155_ (_11733_, _08760_, _08764_);
  and _20156_ (_11734_, _11733_, _08728_);
  or _20157_ (_11735_, _11734_, _11732_);
  and _20158_ (_11736_, _08748_, _11399_);
  and _20159_ (_11737_, _11736_, _08732_);
  and _20160_ (_11738_, _11737_, _08757_);
  and _20161_ (_11739_, _11410_, _11390_);
  or _20162_ (_11740_, _11739_, _11738_);
  nor _20163_ (_11741_, _11740_, _11735_);
  or _20164_ (_11742_, _11741_, _11730_);
  and _20165_ (_11743_, _11742_, _11729_);
  not _20166_ (_11744_, _11421_);
  and _20167_ (_11745_, _11411_, _08717_);
  nor _20168_ (_11746_, _11745_, _11423_);
  nor _20169_ (_11747_, _11746_, _11744_);
  and _20170_ (_11748_, _11738_, _11385_);
  nor _20171_ (_11749_, _11748_, _11747_);
  nor _20172_ (_11750_, _11749_, _11433_);
  nor _20173_ (_11751_, _11750_, _11743_);
  and _20174_ (_11752_, _11751_, _11728_);
  and _20175_ (_11753_, _11752_, _11727_);
  not _20176_ (_11754_, _07108_);
  or _20177_ (_11755_, _07324_, _07297_);
  and _20178_ (_11756_, _07323_, _07320_);
  nor _20179_ (_11757_, _11756_, _11755_);
  and _20180_ (_11758_, _11756_, _11755_);
  nor _20181_ (_11759_, _11758_, _11757_);
  nor _20182_ (_11760_, _11759_, _07531_);
  not _20183_ (_11761_, _07296_);
  and _20184_ (_11762_, _07531_, _11761_);
  or _20185_ (_11763_, _11762_, _11760_);
  or _20186_ (_11764_, _11763_, _11754_);
  not _20187_ (_11765_, _07344_);
  or _20188_ (_11766_, _07751_, _11765_);
  and _20189_ (_11768_, _06731_, _06725_);
  or _20190_ (_11769_, _11768_, _06716_);
  nor _20191_ (_11770_, _11769_, _06732_);
  not _20192_ (_11771_, _11770_);
  and _20193_ (_11772_, _06699_, _06685_);
  nor _20194_ (_11773_, _11772_, _06700_);
  nor _20195_ (_11774_, _11773_, _06616_);
  not _20196_ (_11775_, _11774_);
  or _20197_ (_11776_, _07411_, _06166_);
  and _20198_ (_11777_, _06352_, _06251_);
  and _20199_ (_11778_, _06349_, _06305_);
  nor _20200_ (_11779_, _11778_, _11777_);
  and _20201_ (_11780_, _11779_, _11776_);
  and _20202_ (_11781_, _11780_, _07940_);
  nor _20203_ (_11782_, _06252_, _10897_);
  or _20204_ (_11783_, _11782_, _06305_);
  nand _20205_ (_11784_, _11783_, _07696_);
  and _20206_ (_11785_, _11784_, _07937_);
  and _20207_ (_11786_, _11785_, _07934_);
  and _20208_ (_11787_, _11786_, _11781_);
  and _20209_ (_11788_, _11787_, _11775_);
  and _20210_ (_11789_, _11788_, _11771_);
  and _20211_ (_11790_, _11789_, _11766_);
  and _20212_ (_11791_, _11790_, _11764_);
  nor _20213_ (_11792_, _11791_, _11428_);
  and _20214_ (_11793_, _11732_, _11385_);
  not _20215_ (_11794_, _11793_);
  and _20216_ (_11795_, \oc8051_top_1.oc8051_decoder1.state [0], _05686_);
  not _20217_ (_11796_, _11406_);
  and _20218_ (_11797_, _11793_, _08746_);
  nor _20219_ (_11798_, _11797_, _11796_);
  nor _20220_ (_11799_, _11798_, _11795_);
  and _20221_ (_11800_, _11799_, _11794_);
  and _20222_ (_11801_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _20223_ (_11802_, _11388_, _08764_);
  and _20224_ (_11803_, _11802_, _08757_);
  nor _20225_ (_11804_, _11803_, _11738_);
  and _20226_ (_11805_, _08760_, _08732_);
  and _20227_ (_11806_, _11805_, _08757_);
  not _20228_ (_11807_, _11806_);
  and _20229_ (_11808_, _11807_, _11804_);
  and _20230_ (_11810_, _11394_, _08727_);
  and _20231_ (_11811_, _11802_, _11810_);
  and _20232_ (_11812_, _11733_, _11810_);
  nor _20233_ (_11813_, _11812_, _11811_);
  and _20234_ (_11814_, _11813_, _11808_);
  nor _20235_ (_11815_, _11814_, _11744_);
  not _20236_ (_11816_, _11815_);
  and _20237_ (_11817_, _11811_, _05686_);
  and _20238_ (_11818_, _11812_, _05686_);
  nor _20239_ (_11819_, _11818_, _11817_);
  nor _20240_ (_11821_, _11819_, _06526_);
  nor _20241_ (_11822_, _11821_, _11793_);
  and _20242_ (_11823_, _11822_, _11816_);
  nor _20243_ (_11824_, _11823_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _20244_ (_11825_, _11824_, _11801_);
  and _20245_ (_11826_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _20246_ (_11827_, _11428_);
  and _20247_ (_11828_, _11737_, _11422_);
  not _20248_ (_11829_, _11828_);
  and _20249_ (_11830_, _11731_, _08746_);
  and _20250_ (_11831_, _11830_, _08764_);
  and _20251_ (_11833_, _11831_, _08757_);
  and _20252_ (_11834_, _11831_, _11422_);
  nor _20253_ (_11835_, _11834_, _11833_);
  and _20254_ (_11836_, _11835_, _11829_);
  and _20255_ (_11837_, _11414_, _08728_);
  not _20256_ (_11838_, _11837_);
  and _20257_ (_11839_, _11422_, _11414_);
  and _20258_ (_11840_, _11408_, _08764_);
  and _20259_ (_11841_, _11840_, _11422_);
  nor _20260_ (_11842_, _11841_, _11839_);
  nand _20261_ (_11843_, _11842_, _11838_);
  and _20262_ (_11844_, _11831_, _11412_);
  and _20263_ (_11845_, _11802_, _08728_);
  nor _20264_ (_11846_, _11845_, _11844_);
  and _20265_ (_11847_, _11412_, _11401_);
  nor _20266_ (_11848_, _11847_, _11413_);
  nand _20267_ (_11849_, _11848_, _11846_);
  nor _20268_ (_11850_, _11849_, _11843_);
  and _20269_ (_11851_, _11850_, _11836_);
  and _20270_ (_11852_, _11736_, _08764_);
  and _20271_ (_11853_, _11852_, _08757_);
  and _20272_ (_11854_, _11852_, _11422_);
  nor _20273_ (_11855_, _11854_, _11853_);
  and _20274_ (_11856_, _11414_, _11412_);
  and _20275_ (_11857_, _11733_, _11412_);
  nor _20276_ (_11858_, _11857_, _11856_);
  and _20277_ (_11859_, _11840_, _11412_);
  and _20278_ (_11860_, _11408_, _08728_);
  nor _20279_ (_11861_, _11860_, _11859_);
  and _20280_ (_11862_, _11861_, _11858_);
  and _20281_ (_11863_, _11862_, _11855_);
  and _20282_ (_11864_, _11852_, _11412_);
  and _20283_ (_11865_, _11422_, _11410_);
  nor _20284_ (_11866_, _11865_, _11864_);
  and _20285_ (_11867_, _11830_, _08732_);
  and _20286_ (_11868_, _11867_, _08756_);
  and _20287_ (_11869_, _11733_, _11422_);
  nor _20288_ (_11870_, _11869_, _11868_);
  and _20289_ (_11872_, _11870_, _11866_);
  and _20290_ (_11873_, _11872_, _11863_);
  and _20291_ (_11874_, _11395_, _08764_);
  and _20292_ (_11875_, _11874_, _11388_);
  and _20293_ (_11876_, _11802_, _11422_);
  nor _20294_ (_11877_, _11876_, _11875_);
  nor _20295_ (_11878_, _11867_, _11404_);
  not _20296_ (_11879_, _11878_);
  and _20297_ (_11880_, _11879_, _11412_);
  and _20298_ (_11881_, _11805_, _11422_);
  nor _20299_ (_11882_, _11881_, _11880_);
  and _20300_ (_11883_, _11882_, _11877_);
  and _20301_ (_11884_, _11400_, _08764_);
  and _20302_ (_11885_, _11884_, _11412_);
  and _20303_ (_11887_, _11412_, _08765_);
  nor _20304_ (_11888_, _11887_, _11885_);
  nor _20305_ (_11889_, _08732_, _08715_);
  and _20306_ (_11890_, _11889_, _11388_);
  and _20307_ (_11891_, _11805_, _11412_);
  nor _20308_ (_11893_, _11891_, _11890_);
  and _20309_ (_11894_, _11893_, _11888_);
  not _20310_ (_11895_, _11427_);
  and _20311_ (_11896_, _11895_, _11406_);
  and _20312_ (_11897_, _11896_, _11894_);
  and _20313_ (_11899_, _11897_, _11883_);
  and _20314_ (_11900_, _11899_, _11873_);
  and _20315_ (_11901_, _11900_, _11851_);
  nor _20316_ (_11902_, _11901_, _11744_);
  nor _20317_ (_11903_, _11902_, _11827_);
  and _20318_ (_11904_, _11903_, _11794_);
  nor _20319_ (_11905_, _11904_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _20320_ (_11906_, _11905_, _11826_);
  and _20321_ (_11907_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _20322_ (_11908_, _11408_, _11395_);
  and _20323_ (_11909_, _11805_, _11395_);
  nor _20324_ (_11910_, _11909_, _11908_);
  or _20325_ (_11911_, _11414_, _11400_);
  and _20326_ (_11912_, _11911_, _11395_);
  nor _20327_ (_11913_, _11912_, _11427_);
  and _20328_ (_11914_, _11913_, _11910_);
  or _20329_ (_11915_, _11879_, _11831_);
  and _20330_ (_11916_, _11915_, _11395_);
  and _20331_ (_11917_, _11733_, _11395_);
  and _20332_ (_11918_, _11852_, _11395_);
  or _20333_ (_11919_, _11918_, _11917_);
  and _20334_ (_11920_, _11410_, _08728_);
  and _20335_ (_11921_, _11395_, _08765_);
  or _20336_ (_11922_, _11921_, _11920_);
  or _20337_ (_11923_, _11922_, _11919_);
  nor _20338_ (_11924_, _11923_, _11916_);
  and _20339_ (_11925_, _11924_, _11914_);
  and _20340_ (_11926_, _11925_, _11808_);
  nor _20341_ (_11927_, _11926_, _11744_);
  nor _20342_ (_11928_, _11799_, _11794_);
  nor _20343_ (_11929_, _11928_, _11827_);
  not _20344_ (_11930_, _11929_);
  nor _20345_ (_11931_, _11930_, _11927_);
  nor _20346_ (_11932_, _11931_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _20347_ (_11933_, _11932_, _11907_);
  nor _20348_ (_11934_, _11933_, _11906_);
  and _20349_ (_11935_, _11934_, _11825_);
  and _20350_ (_11936_, _06363_, _06012_);
  and _20351_ (_11937_, _11936_, _06840_);
  not _20352_ (_11938_, _11937_);
  nor _20353_ (_11939_, _11938_, _07945_);
  and _20354_ (_11940_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _20355_ (_11942_, _11940_, _11939_);
  and _20356_ (_11943_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _20357_ (_11944_, _11938_, _06434_);
  nor _20358_ (_11945_, _11944_, _11943_);
  and _20359_ (_11946_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _20360_ (_11947_, _11938_, _09037_);
  nor _20361_ (_11948_, _11947_, _11946_);
  nor _20362_ (_11949_, _11937_, _05997_);
  and _20363_ (_11950_, _11937_, _07978_);
  nor _20364_ (_11951_, _11950_, _11949_);
  and _20365_ (_11952_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _20366_ (_11953_, _11952_, _11948_);
  and _20367_ (_11954_, _11953_, _11945_);
  and _20368_ (_11955_, _11954_, _11942_);
  nor _20369_ (_11956_, _11954_, _11942_);
  or _20370_ (_11957_, _11956_, _11955_);
  and _20371_ (_11958_, _11957_, _05899_);
  or _20372_ (_11959_, _11958_, _06017_);
  and _20373_ (_11960_, _11959_, _11938_);
  or _20374_ (_11961_, _11960_, _11939_);
  and _20375_ (_11962_, _11961_, _11935_);
  not _20376_ (_11963_, _11962_);
  and _20377_ (_11964_, _08985_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _20378_ (_11965_, _11964_, _10893_);
  not _20379_ (_11966_, _11965_);
  and _20380_ (_11967_, _11933_, _11825_);
  and _20381_ (_11968_, _11967_, _11906_);
  and _20382_ (_11969_, _11968_, _11966_);
  not _20383_ (_11970_, _11933_);
  and _20384_ (_11971_, _11970_, _11906_);
  and _20385_ (_11972_, _11971_, _11825_);
  and _20386_ (_11973_, _05923_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _20387_ (_11974_, _08991_, _06364_);
  nor _20388_ (_11975_, _11974_, _11973_);
  and _20389_ (_11976_, _11965_, _06378_);
  not _20390_ (_11977_, _11976_);
  nor _20391_ (_11978_, _11965_, _06378_);
  not _20392_ (_11979_, _11978_);
  and _20393_ (_11980_, _08721_, _06030_);
  and _20394_ (_11981_, _08753_, _06004_);
  or _20395_ (_11982_, _11981_, _11980_);
  nor _20396_ (_11983_, _11982_, _09348_);
  and _20397_ (_11984_, _11983_, _11979_);
  and _20398_ (_11985_, _11984_, _11977_);
  and _20399_ (_11986_, _11985_, _11975_);
  not _20400_ (_11987_, _08991_);
  nor _20401_ (_11989_, _11965_, _08721_);
  and _20402_ (_11990_, _11989_, _11987_);
  and _20403_ (_11991_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _20404_ (_11992_, _11965_, _08721_);
  and _20405_ (_11993_, _11992_, _08991_);
  and _20406_ (_11994_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _20407_ (_11995_, _11994_, _11991_);
  nor _20408_ (_11996_, _11965_, _08753_);
  and _20409_ (_11997_, _11996_, _08991_);
  and _20410_ (_11998_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _20411_ (_11999_, _11965_, _08753_);
  and _20412_ (_12000_, _11999_, _11987_);
  and _20413_ (_12001_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _20414_ (_12002_, _12001_, _11998_);
  and _20415_ (_12003_, _12002_, _11995_);
  and _20416_ (_12004_, _11992_, _11987_);
  and _20417_ (_12005_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _20418_ (_12006_, _11999_, _08991_);
  and _20419_ (_12007_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _20420_ (_12008_, _12007_, _12005_);
  and _20421_ (_12009_, _11996_, _11987_);
  and _20422_ (_12010_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _20423_ (_12011_, _11989_, _08991_);
  and _20424_ (_12013_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _20425_ (_12014_, _12013_, _12010_);
  and _20426_ (_12015_, _12014_, _12008_);
  and _20427_ (_12016_, _12015_, _12003_);
  nor _20428_ (_12017_, _12016_, _11986_);
  not _20429_ (_12019_, _07945_);
  and _20430_ (_12020_, _11986_, _12019_);
  nor _20431_ (_12021_, _12020_, _12017_);
  not _20432_ (_12022_, _12021_);
  and _20433_ (_12023_, _12022_, _11972_);
  not _20434_ (_12024_, _11607_);
  nor _20435_ (_12025_, _11970_, _11906_);
  and _20436_ (_12026_, _12025_, _11825_);
  and _20437_ (_12027_, _12026_, _12024_);
  or _20438_ (_12028_, _12027_, _12023_);
  nor _20439_ (_12029_, _12028_, _11969_);
  and _20440_ (_12030_, _12029_, _11963_);
  nor _20441_ (_12031_, _12030_, _06378_);
  and _20442_ (_12032_, _12030_, _06378_);
  nor _20443_ (_12033_, _12032_, _12031_);
  and _20444_ (_12034_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _20445_ (_12035_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _20446_ (_12036_, _12035_, _12034_);
  and _20447_ (_12037_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _20448_ (_12038_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _20449_ (_12039_, _12038_, _12037_);
  and _20450_ (_12040_, _12039_, _12036_);
  and _20451_ (_12041_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _20452_ (_12042_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _20453_ (_12043_, _12042_, _12041_);
  and _20454_ (_12044_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _20455_ (_12045_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _20456_ (_12046_, _12045_, _12044_);
  and _20457_ (_12047_, _12046_, _12043_);
  and _20458_ (_12049_, _12047_, _12040_);
  nor _20459_ (_12050_, _12049_, _11986_);
  and _20460_ (_12051_, _11986_, _06360_);
  nor _20461_ (_12052_, _12051_, _12050_);
  not _20462_ (_12053_, _12052_);
  and _20463_ (_12054_, _12053_, _11972_);
  not _20464_ (_12055_, _12054_);
  nor _20465_ (_12056_, _11938_, _06359_);
  nor _20466_ (_12057_, _11938_, _06993_);
  and _20467_ (_12058_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _20468_ (_12059_, _12058_, _12057_);
  and _20469_ (_12060_, _12059_, _11955_);
  nor _20470_ (_12061_, _11938_, _06609_);
  and _20471_ (_12062_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _20472_ (_12063_, _12062_, _12061_);
  and _20473_ (_12064_, _12063_, _12060_);
  nor _20474_ (_12065_, _11938_, _09341_);
  and _20475_ (_12066_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _20476_ (_12067_, _12066_, _12065_);
  and _20477_ (_12068_, _12067_, _12064_);
  nor _20478_ (_12069_, _11937_, _05955_);
  nor _20479_ (_12070_, _12069_, _12068_);
  and _20480_ (_12071_, _12069_, _12068_);
  or _20481_ (_12072_, _12071_, _12070_);
  nor _20482_ (_12073_, _12072_, _05898_);
  or _20483_ (_12074_, _12073_, _05959_);
  and _20484_ (_12075_, _12074_, _11938_);
  or _20485_ (_12076_, _12075_, _12056_);
  and _20486_ (_12077_, _12076_, _11934_);
  not _20487_ (_12078_, _12077_);
  not _20488_ (_12079_, _11825_);
  not _20489_ (_12080_, _11469_);
  and _20490_ (_12081_, _12025_, _12080_);
  nor _20491_ (_12082_, _12081_, _12079_);
  and _20492_ (_12083_, _12082_, _12078_);
  and _20493_ (_12084_, _12083_, _12055_);
  nor _20494_ (_12085_, _12084_, _06807_);
  and _20495_ (_12086_, _12084_, _06807_);
  nor _20496_ (_12087_, _12086_, _12085_);
  nor _20497_ (_12088_, _11971_, _11825_);
  not _20498_ (_12090_, _11511_);
  and _20499_ (_12091_, _12026_, _12090_);
  nor _20500_ (_12092_, _12091_, _12088_);
  nor _20501_ (_12093_, _12067_, _12064_);
  nor _20502_ (_12094_, _12093_, _12068_);
  nor _20503_ (_12095_, _12094_, _05898_);
  nor _20504_ (_12096_, _12095_, _05944_);
  nor _20505_ (_12097_, _12096_, _11937_);
  nor _20506_ (_12098_, _12097_, _12065_);
  not _20507_ (_12100_, _12098_);
  and _20508_ (_12102_, _12100_, _11935_);
  and _20509_ (_12103_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _20510_ (_12104_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _20511_ (_12105_, _12104_, _12103_);
  and _20512_ (_12106_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _20513_ (_12107_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _20514_ (_12108_, _12107_, _12106_);
  and _20515_ (_12109_, _12108_, _12105_);
  and _20516_ (_12110_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _20517_ (_12112_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _20518_ (_12113_, _12112_, _12110_);
  and _20519_ (_12114_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _20520_ (_12115_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor _20521_ (_12116_, _12115_, _12114_);
  and _20522_ (_12117_, _12116_, _12113_);
  and _20523_ (_12118_, _12117_, _12109_);
  nor _20524_ (_12119_, _12118_, _11986_);
  not _20525_ (_12120_, _09341_);
  and _20526_ (_12121_, _11986_, _12120_);
  nor _20527_ (_12122_, _12121_, _12119_);
  not _20528_ (_12123_, _12122_);
  and _20529_ (_12124_, _12123_, _11972_);
  nor _20530_ (_12125_, _12124_, _12102_);
  and _20531_ (_12126_, _12125_, _12092_);
  nor _20532_ (_12127_, _12126_, _06819_);
  and _20533_ (_12128_, _12126_, _06819_);
  nor _20534_ (_12129_, _12128_, _12127_);
  and _20535_ (_12130_, _12129_, _12087_);
  not _20536_ (_12131_, _11549_);
  and _20537_ (_12132_, _12026_, _12131_);
  not _20538_ (_12133_, _12025_);
  and _20539_ (_12134_, _12088_, _12133_);
  nor _20540_ (_12135_, _12134_, _12132_);
  nor _20541_ (_12136_, _12063_, _12060_);
  nor _20542_ (_12137_, _12136_, _12064_);
  nor _20543_ (_12138_, _12137_, _05898_);
  nor _20544_ (_12139_, _12138_, _05928_);
  nor _20545_ (_12140_, _12139_, _11937_);
  nor _20546_ (_12142_, _12140_, _12061_);
  not _20547_ (_12143_, _12142_);
  and _20548_ (_12144_, _12143_, _11935_);
  and _20549_ (_12145_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _20550_ (_12146_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _20551_ (_12147_, _12146_, _12145_);
  and _20552_ (_12148_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _20553_ (_12149_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _20554_ (_12150_, _12149_, _12148_);
  and _20555_ (_12151_, _12150_, _12147_);
  and _20556_ (_12152_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _20557_ (_12153_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _20558_ (_12154_, _12153_, _12152_);
  and _20559_ (_12155_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _20560_ (_12156_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _20561_ (_12157_, _12156_, _12155_);
  and _20562_ (_12158_, _12157_, _12154_);
  and _20563_ (_12159_, _12158_, _12151_);
  nor _20564_ (_12160_, _12159_, _11986_);
  not _20565_ (_12161_, _06609_);
  and _20566_ (_12162_, _11986_, _12161_);
  nor _20567_ (_12163_, _12162_, _12160_);
  not _20568_ (_12164_, _12163_);
  and _20569_ (_12165_, _12164_, _11972_);
  nor _20570_ (_12166_, _12165_, _12144_);
  and _20571_ (_12167_, _12166_, _12135_);
  nor _20572_ (_12168_, _12167_, _07767_);
  and _20573_ (_12169_, _12167_, _07767_);
  nor _20574_ (_12171_, _12169_, _12168_);
  not _20575_ (_12172_, _09713_);
  and _20576_ (_12173_, _12026_, _12172_);
  and _20577_ (_12174_, _11968_, _11987_);
  nor _20578_ (_12176_, _12174_, _12173_);
  and _20579_ (_12177_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _20580_ (_12178_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _20581_ (_12180_, _12178_, _12177_);
  and _20582_ (_12182_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _20583_ (_12183_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _20584_ (_12184_, _12183_, _12182_);
  and _20585_ (_12185_, _12184_, _12180_);
  and _20586_ (_12186_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _20587_ (_12187_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _20588_ (_12188_, _12187_, _12186_);
  and _20589_ (_12189_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _20590_ (_12191_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _20591_ (_12192_, _12191_, _12189_);
  and _20592_ (_12194_, _12192_, _12188_);
  and _20593_ (_12195_, _12194_, _12185_);
  nor _20594_ (_12196_, _12195_, _11986_);
  not _20595_ (_12197_, _06993_);
  and _20596_ (_12198_, _11986_, _12197_);
  nor _20597_ (_12199_, _12198_, _12196_);
  not _20598_ (_12201_, _12199_);
  and _20599_ (_12202_, _12201_, _11972_);
  not _20600_ (_12204_, _12202_);
  nor _20601_ (_12205_, _12059_, _11955_);
  nor _20602_ (_12207_, _12205_, _12060_);
  nor _20603_ (_12208_, _12207_, _05898_);
  nor _20604_ (_12209_, _12208_, _05902_);
  nor _20605_ (_12210_, _12209_, _11937_);
  nor _20606_ (_12212_, _12210_, _12057_);
  not _20607_ (_12213_, _12212_);
  and _20608_ (_12215_, _12213_, _11935_);
  and _20609_ (_12216_, _11933_, _12079_);
  nor _20610_ (_12218_, _12216_, _12215_);
  and _20611_ (_12219_, _12218_, _12204_);
  and _20612_ (_12221_, _12219_, _12176_);
  nor _20613_ (_12222_, _12221_, _06364_);
  and _20614_ (_12223_, _12221_, _06364_);
  nor _20615_ (_12224_, _12223_, _12222_);
  and _20616_ (_12225_, _12224_, _12171_);
  and _20617_ (_12227_, _12225_, _12130_);
  and _20618_ (_12228_, _12227_, _12033_);
  nor _20619_ (_12230_, _06805_, _06013_);
  and _20620_ (_12231_, _12230_, _12228_);
  and _20621_ (_12233_, _12231_, _11800_);
  not _20622_ (_12234_, _12233_);
  nor _20623_ (_12236_, _11747_, _11827_);
  not _20624_ (_12237_, _12236_);
  not _20625_ (_12238_, _07792_);
  not _20626_ (_12239_, _11799_);
  not _20627_ (_12240_, _07687_);
  nor _20628_ (_12241_, _06689_, _06687_);
  and _20629_ (_12242_, _12241_, _11773_);
  nor _20630_ (_12243_, _11793_, _08039_);
  and _20631_ (_12244_, _12243_, _12242_);
  and _20632_ (_12245_, _12244_, _12240_);
  and _20633_ (_12246_, _12245_, _12239_);
  and _20634_ (_12247_, _12246_, _07612_);
  and _20635_ (_12248_, _12247_, _07368_);
  and _20636_ (_12249_, _12248_, _12238_);
  not _20637_ (_12250_, _12249_);
  nor _20638_ (_12251_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _20639_ (_12252_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _20640_ (_12253_, _12252_, _12251_);
  nor _20641_ (_12255_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _20642_ (_12256_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _20643_ (_12257_, _12256_, _12255_);
  and _20644_ (_12258_, _12257_, _12253_);
  and _20645_ (_12259_, _12258_, _11928_);
  not _20646_ (_12260_, _12259_);
  and _20647_ (_12262_, _11800_, _06118_);
  and _20648_ (_12263_, _11797_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _20649_ (_12264_, _12263_, _12262_);
  and _20650_ (_12266_, _12264_, _12260_);
  and _20651_ (_12267_, _12266_, _12250_);
  and _20652_ (_12268_, _11405_, _08764_);
  or _20653_ (_12269_, _12268_, _11403_);
  and _20654_ (_12270_, _11732_, _08764_);
  nor _20655_ (_12271_, _12270_, _12269_);
  not _20656_ (_12272_, _12271_);
  nor _20657_ (_12273_, _12272_, _12267_);
  and _20658_ (_12274_, _11405_, _08732_);
  nor _20659_ (_12275_, _12274_, _11739_);
  and _20660_ (_12276_, _11732_, _08732_);
  not _20661_ (_12277_, _12276_);
  and _20662_ (_12278_, _12277_, _11417_);
  and _20663_ (_12279_, _12278_, _12275_);
  and _20664_ (_12280_, _12279_, _11398_);
  and _20665_ (_12282_, _12280_, _12267_);
  nor _20666_ (_12283_, _12282_, _12273_);
  nor _20667_ (_12284_, _11738_, _11734_);
  and _20668_ (_12285_, _12284_, _11895_);
  not _20669_ (_12286_, _12285_);
  nor _20670_ (_12288_, _12286_, _12283_);
  nor _20671_ (_12289_, _12288_, _11730_);
  nor _20672_ (_12291_, _12289_, _12237_);
  not _20673_ (_12292_, _08941_);
  and _20674_ (_12294_, _11928_, _12292_);
  nor _20675_ (_12295_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and _20676_ (_12296_, _12295_, _08985_);
  and _20677_ (_12297_, _12296_, _10935_);
  not _20678_ (_12298_, _12297_);
  and _20679_ (_12299_, _12298_, _11797_);
  nor _20680_ (_12301_, _12299_, _12294_);
  not _20681_ (_12302_, _12301_);
  nor _20682_ (_12304_, _12302_, _12291_);
  and _20683_ (_12305_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _20684_ (_12306_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _20685_ (_12307_, _12306_, _12305_);
  and _20686_ (_12308_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _20687_ (_12309_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _20688_ (_12310_, _12309_, _12308_);
  and _20689_ (_12311_, _12310_, _12307_);
  and _20690_ (_12312_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _20691_ (_12313_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _20692_ (_12314_, _12313_, _12312_);
  and _20693_ (_12316_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _20694_ (_12317_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _20695_ (_12318_, _12317_, _12316_);
  and _20696_ (_12319_, _12318_, _12314_);
  and _20697_ (_12320_, _12319_, _12311_);
  nor _20698_ (_12321_, _12320_, _11986_);
  and _20699_ (_12322_, _11986_, _07978_);
  nor _20700_ (_12323_, _12322_, _12321_);
  not _20701_ (_12324_, _12323_);
  and _20702_ (_12325_, _12324_, _11972_);
  and _20703_ (_12326_, _12026_, _11689_);
  nor _20704_ (_12328_, _12326_, _12325_);
  nor _20705_ (_12329_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _20706_ (_12330_, _12329_, _11952_);
  nor _20707_ (_12332_, _12330_, _05898_);
  nor _20708_ (_12333_, _12332_, _05998_);
  nor _20709_ (_12335_, _12333_, _11937_);
  nor _20710_ (_12336_, _12335_, _11950_);
  not _20711_ (_12337_, _12336_);
  and _20712_ (_12338_, _12337_, _11935_);
  and _20713_ (_12339_, _11968_, _08753_);
  nor _20714_ (_12340_, _12339_, _12338_);
  and _20715_ (_12341_, _12340_, _12328_);
  and _20716_ (_12343_, _12341_, _06030_);
  nor _20717_ (_12344_, _12341_, _06030_);
  or _20718_ (_12346_, _12344_, _12343_);
  nor _20719_ (_12347_, _12346_, _06827_);
  and _20720_ (_12348_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _20721_ (_12349_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _20722_ (_12350_, _12349_, _12348_);
  and _20723_ (_12351_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _20724_ (_12352_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _20725_ (_12353_, _12352_, _12351_);
  and _20726_ (_12354_, _12353_, _12350_);
  and _20727_ (_12355_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _20728_ (_12356_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _20729_ (_12357_, _12356_, _12355_);
  and _20730_ (_12359_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _20731_ (_12360_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _20732_ (_12362_, _12360_, _12359_);
  and _20733_ (_12363_, _12362_, _12357_);
  and _20734_ (_12364_, _12363_, _12354_);
  nor _20735_ (_12365_, _12364_, _11986_);
  and _20736_ (_12366_, _11986_, _11023_);
  nor _20737_ (_12368_, _12366_, _12365_);
  not _20738_ (_12369_, _12368_);
  and _20739_ (_12370_, _12369_, _11972_);
  and _20740_ (_12371_, _11971_, _12079_);
  nor _20741_ (_12372_, _11952_, _11948_);
  nor _20742_ (_12374_, _12372_, _11953_);
  nor _20743_ (_12375_, _12374_, _05898_);
  nor _20744_ (_12376_, _12375_, _05985_);
  nor _20745_ (_12377_, _12376_, _11937_);
  nor _20746_ (_12378_, _12377_, _11947_);
  not _20747_ (_12379_, _12378_);
  and _20748_ (_12380_, _12379_, _11935_);
  or _20749_ (_12381_, _12380_, _12371_);
  and _20750_ (_12382_, _12026_, _11651_);
  and _20751_ (_12383_, _11968_, _08725_);
  or _20752_ (_12384_, _12383_, _12382_);
  or _20753_ (_12385_, _12384_, _12381_);
  nor _20754_ (_12386_, _12385_, _12370_);
  nor _20755_ (_12387_, _12386_, _05993_);
  and _20756_ (_12388_, _12386_, _05993_);
  nor _20757_ (_12389_, _12388_, _12387_);
  nor _20758_ (_12390_, _11953_, _11945_);
  nor _20759_ (_12391_, _12390_, _11954_);
  nor _20760_ (_12393_, _12391_, _05898_);
  nor _20761_ (_12394_, _12393_, _05972_);
  nor _20762_ (_12395_, _12394_, _11937_);
  nor _20763_ (_12397_, _12395_, _11944_);
  not _20764_ (_12398_, _12397_);
  and _20765_ (_12399_, _12398_, _11935_);
  not _20766_ (_12400_, _12399_);
  and _20767_ (_12401_, _11968_, _11392_);
  and _20768_ (_12402_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _20769_ (_12403_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _20770_ (_12404_, _12403_, _12402_);
  and _20771_ (_12405_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _20772_ (_12406_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _20773_ (_12407_, _12406_, _12405_);
  and _20774_ (_12408_, _12407_, _12404_);
  and _20775_ (_12409_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _20776_ (_12410_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _20777_ (_12411_, _12410_, _12409_);
  and _20778_ (_12412_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _20779_ (_12413_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _20780_ (_12414_, _12413_, _12412_);
  and _20781_ (_12416_, _12414_, _12411_);
  and _20782_ (_12417_, _12416_, _12408_);
  nor _20783_ (_12418_, _12417_, _11986_);
  and _20784_ (_12419_, _11986_, _06435_);
  nor _20785_ (_12420_, _12419_, _12418_);
  not _20786_ (_12421_, _12420_);
  and _20787_ (_12422_, _12421_, _11972_);
  and _20788_ (_12423_, _12026_, _11628_);
  or _20789_ (_12424_, _12423_, _12422_);
  nor _20790_ (_12425_, _12424_, _12401_);
  and _20791_ (_12426_, _12425_, _12400_);
  nor _20792_ (_12427_, _12426_, _05981_);
  and _20793_ (_12428_, _12426_, _05981_);
  nor _20794_ (_12429_, _12428_, _12427_);
  nor _20795_ (_12430_, _12429_, _12389_);
  and _20796_ (_12431_, _12430_, _12347_);
  and _20797_ (_12432_, _12431_, _12228_);
  nor _20798_ (_12433_, _05967_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _20799_ (_12434_, _12433_, _12432_);
  not _20800_ (_12435_, _12434_);
  and _20801_ (_12436_, _12435_, _12304_);
  and _20802_ (_12437_, _12436_, _12234_);
  not _20803_ (_12438_, _11748_);
  and _20804_ (_12439_, _07494_, _07479_);
  not _20805_ (_12441_, _12439_);
  and _20806_ (_12442_, _07495_, _06715_);
  and _20807_ (_12443_, _12442_, _12441_);
  not _20808_ (_12444_, _12443_);
  and _20809_ (_12445_, _07920_, _07344_);
  not _20810_ (_12446_, _12445_);
  nor _20811_ (_12447_, _07442_, _06302_);
  and _20812_ (_12449_, _07573_, _06660_);
  nor _20813_ (_12450_, _12449_, _06120_);
  nor _20814_ (_12451_, _12450_, _12447_);
  and _20815_ (_12452_, _12451_, _06701_);
  nor _20816_ (_12453_, _12451_, _06701_);
  nor _20817_ (_12454_, _12453_, _12452_);
  and _20818_ (_12455_, _12454_, _06145_);
  and _20819_ (_12456_, _06701_, _06349_);
  nor _20820_ (_12457_, _06187_, _06128_);
  and _20821_ (_12458_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _20822_ (_12459_, _12458_, _12457_);
  or _20823_ (_12460_, _12459_, _06779_);
  nor _20824_ (_12462_, _12460_, _12456_);
  not _20825_ (_12463_, _12462_);
  nor _20826_ (_12464_, _12463_, _12455_);
  and _20827_ (_12465_, _12464_, _12446_);
  and _20828_ (_12466_, _12465_, _12444_);
  nor _20829_ (_12467_, _12466_, _12438_);
  and _20830_ (_12469_, _11750_, _11743_);
  and _20831_ (_12470_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _20832_ (_12472_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20833_ (_12473_, _12472_, _12470_);
  and _20834_ (_12474_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _20835_ (_12475_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _20836_ (_12476_, _12475_, _12474_);
  and _20837_ (_12477_, _12476_, _11722_);
  and _20838_ (_12478_, _12477_, _12473_);
  and _20839_ (_12479_, _12478_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _20840_ (_12480_, _12478_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _20841_ (_12481_, _12480_, _12479_);
  and _20842_ (_12482_, _12481_, _12469_);
  and _20843_ (_12483_, _12024_, _11424_);
  and _20844_ (_12484_, _11749_, _11455_);
  and _20845_ (_12485_, _12484_, _11743_);
  and _20846_ (_12486_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _20847_ (_12487_, _12486_, _12483_);
  or _20848_ (_12488_, _12487_, _12482_);
  nor _20849_ (_12489_, _12488_, _12467_);
  nand _20850_ (_12491_, _12489_, _12437_);
  or _20851_ (_12492_, _12491_, _11792_);
  or _20852_ (_12493_, _12492_, _11753_);
  not _20853_ (_12494_, _06530_);
  and _20854_ (_12495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _20855_ (_12497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _20856_ (_12498_, _12497_, _12495_);
  and _20857_ (_12499_, _12498_, _11250_);
  and _20858_ (_12500_, _12499_, _12494_);
  and _20859_ (_12501_, _12500_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _20860_ (_12502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _20861_ (_12503_, _12502_, _12501_);
  nor _20862_ (_12504_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _20863_ (_12505_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _20864_ (_12506_, _12505_, _12504_);
  or _20865_ (_12507_, _12506_, _12437_);
  and _20866_ (_12508_, _12507_, _06071_);
  and _20867_ (_11409_, _12508_, _12493_);
  nor _20868_ (_11432_, _12368_, rst);
  or _20869_ (_12509_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  nand _20870_ (_12510_, _06530_, _10995_);
  and _20871_ (_12511_, _12510_, _06071_);
  and _20872_ (_11437_, _12511_, _12509_);
  or _20873_ (_12512_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _20874_ (_12513_, _06530_, _05739_);
  and _20875_ (_12514_, _12513_, _06071_);
  and _20876_ (_11440_, _12514_, _12512_);
  and _20877_ (_11443_, _08725_, _06071_);
  nor _20878_ (_12515_, _06993_, _06996_);
  and _20879_ (_12516_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _20880_ (_12517_, _12516_, _06390_);
  or _20881_ (_12518_, _12517_, _12515_);
  or _20882_ (_12519_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _20883_ (_12520_, _12519_, _06071_);
  and _20884_ (_11489_, _12520_, _12518_);
  or _20885_ (_12521_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _20886_ (_12522_, _06530_, _05693_);
  and _20887_ (_12523_, _12522_, _06071_);
  and _20888_ (_11494_, _12523_, _12521_);
  and _20889_ (_12524_, _06071_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _20890_ (_12525_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _20891_ (_12527_, _11874_, _11731_);
  or _20892_ (_12528_, _12527_, _11908_);
  or _20893_ (_12529_, _11879_, _11852_);
  and _20894_ (_12530_, _12529_, _11810_);
  or _20895_ (_12531_, _12530_, _12528_);
  and _20896_ (_12532_, _08761_, _08764_);
  and _20897_ (_12533_, _11831_, _11810_);
  or _20898_ (_12534_, _12533_, _11844_);
  and _20899_ (_12535_, _11805_, _08728_);
  or _20900_ (_12536_, _12535_, _12534_);
  or _20901_ (_12537_, _12536_, _12532_);
  or _20902_ (_12538_, _12537_, _12531_);
  or _20903_ (_12539_, _11864_, _11859_);
  or _20904_ (_12540_, _12539_, _11834_);
  and _20905_ (_12541_, _11889_, _11736_);
  and _20906_ (_12542_, _11889_, _11407_);
  or _20907_ (_12543_, _12542_, _12541_);
  or _20908_ (_12544_, _12543_, _11854_);
  or _20909_ (_12545_, _12544_, _12540_);
  not _20910_ (_12546_, _11398_);
  and _20911_ (_12547_, _11805_, _11810_);
  and _20912_ (_12548_, _11810_, _11414_);
  and _20913_ (_12549_, _11810_, _08765_);
  or _20914_ (_12550_, _12549_, _12548_);
  or _20915_ (_12551_, _12550_, _12547_);
  or _20916_ (_12552_, _12551_, _12546_);
  or _20917_ (_12553_, _12552_, _12545_);
  or _20918_ (_12555_, _12553_, _12538_);
  and _20919_ (_12556_, _12555_, _08775_);
  or _20920_ (_11499_, _12556_, _12525_);
  and _20921_ (_12558_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _06071_);
  and _20922_ (_11502_, _12558_, _05811_);
  and _20923_ (_12559_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor _20924_ (_12561_, _08865_, _06609_);
  or _20925_ (_12562_, _12561_, _12559_);
  and _20926_ (_11544_, _12562_, _06071_);
  and _20927_ (_12563_, _08254_, word_in[0]);
  nand _20928_ (_12564_, _08174_, _09175_);
  or _20929_ (_12565_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _20930_ (_12566_, _12565_, _12564_);
  and _20931_ (_12567_, _12566_, _08196_);
  or _20932_ (_12568_, _12567_, _08184_);
  nand _20933_ (_12569_, _08174_, _09726_);
  or _20934_ (_12570_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _20935_ (_12571_, _12570_, _12569_);
  and _20936_ (_12572_, _12571_, _08221_);
  nand _20937_ (_12573_, _08174_, _09936_);
  or _20938_ (_12574_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _20939_ (_12575_, _12574_, _12573_);
  and _20940_ (_12576_, _12575_, _08200_);
  nand _20941_ (_12577_, _08174_, _09476_);
  or _20942_ (_12578_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _20943_ (_12579_, _12578_, _12577_);
  and _20944_ (_12580_, _12579_, _08208_);
  or _20945_ (_12581_, _12580_, _12576_);
  or _20946_ (_12582_, _12581_, _12572_);
  or _20947_ (_12583_, _12582_, _12568_);
  nand _20948_ (_12584_, _08174_, _10161_);
  or _20949_ (_12585_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _20950_ (_12586_, _12585_, _12584_);
  and _20951_ (_12587_, _12586_, _08196_);
  or _20952_ (_12588_, _12587_, _08281_);
  nand _20953_ (_12589_, _08174_, _10589_);
  or _20954_ (_12590_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _20955_ (_12591_, _12590_, _12589_);
  and _20956_ (_12592_, _12591_, _08221_);
  nand _20957_ (_12593_, _08174_, _10795_);
  or _20958_ (_12594_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _20959_ (_12595_, _12594_, _12593_);
  and _20960_ (_12596_, _12595_, _08200_);
  nand _20961_ (_12597_, _08174_, _10371_);
  or _20962_ (_12598_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _20963_ (_12599_, _12598_, _12597_);
  and _20964_ (_12601_, _12599_, _08208_);
  or _20965_ (_12602_, _12601_, _12596_);
  or _20966_ (_12603_, _12602_, _12592_);
  or _20967_ (_12604_, _12603_, _12588_);
  and _20968_ (_12605_, _12604_, _12583_);
  and _20969_ (_12606_, _12605_, _08253_);
  or _20970_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12606_, _12563_);
  and _20971_ (_12607_, _08254_, word_in[1]);
  nand _20972_ (_12608_, _08174_, _09490_);
  or _20973_ (_12609_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _20974_ (_12610_, _12609_, _12608_);
  and _20975_ (_12611_, _12610_, _08208_);
  or _20976_ (_12612_, _12611_, _08184_);
  nand _20977_ (_12613_, _08174_, _09740_);
  or _20978_ (_12614_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _20979_ (_12615_, _12614_, _12613_);
  and _20980_ (_12616_, _12615_, _08221_);
  nand _20981_ (_12617_, _08174_, _09950_);
  or _20982_ (_12618_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _20983_ (_12619_, _12618_, _12617_);
  and _20984_ (_12620_, _12619_, _08200_);
  nand _20985_ (_12621_, _08174_, _09197_);
  or _20986_ (_12622_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _20987_ (_12623_, _12622_, _12621_);
  and _20988_ (_12625_, _12623_, _08196_);
  or _20989_ (_12626_, _12625_, _12620_);
  or _20990_ (_12627_, _12626_, _12616_);
  or _20991_ (_12628_, _12627_, _12612_);
  nand _20992_ (_12629_, _08174_, _10387_);
  or _20993_ (_12630_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _20994_ (_12631_, _12630_, _12629_);
  and _20995_ (_12632_, _12631_, _08208_);
  or _20996_ (_12633_, _12632_, _08281_);
  nand _20997_ (_12634_, _08174_, _10809_);
  or _20998_ (_12635_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _20999_ (_12636_, _12635_, _12634_);
  and _21000_ (_12637_, _12636_, _08200_);
  nand _21001_ (_12638_, _08174_, _10606_);
  or _21002_ (_12639_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _21003_ (_12640_, _12639_, _12638_);
  and _21004_ (_12641_, _12640_, _08221_);
  or _21005_ (_12642_, _12641_, _12637_);
  nand _21006_ (_12643_, _08174_, _10177_);
  or _21007_ (_12644_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _21008_ (_12645_, _12644_, _12643_);
  and _21009_ (_12646_, _12645_, _08196_);
  or _21010_ (_12647_, _12646_, _12642_);
  or _21011_ (_12648_, _12647_, _12633_);
  and _21012_ (_12649_, _12648_, _12628_);
  and _21013_ (_12650_, _12649_, _08253_);
  or _21014_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12650_, _12607_);
  and _21015_ (_12651_, _08254_, word_in[2]);
  nand _21016_ (_12652_, _08174_, _09502_);
  or _21017_ (_12653_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _21018_ (_12654_, _12653_, _12652_);
  and _21019_ (_12655_, _12654_, _08208_);
  or _21020_ (_12656_, _12655_, _08184_);
  nand _21021_ (_12657_, _08174_, _09752_);
  or _21022_ (_12658_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _21023_ (_12659_, _12658_, _12657_);
  and _21024_ (_12660_, _12659_, _08221_);
  nand _21025_ (_12661_, _08174_, _09965_);
  or _21026_ (_12662_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _21027_ (_12663_, _12662_, _12661_);
  and _21028_ (_12664_, _12663_, _08200_);
  nand _21029_ (_12665_, _08174_, _09208_);
  or _21030_ (_12666_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _21031_ (_12667_, _12666_, _12665_);
  and _21032_ (_12668_, _12667_, _08196_);
  or _21033_ (_12669_, _12668_, _12664_);
  or _21034_ (_12670_, _12669_, _12660_);
  or _21035_ (_12671_, _12670_, _12656_);
  nand _21036_ (_12672_, _08174_, _10399_);
  or _21037_ (_12673_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _21038_ (_12674_, _12673_, _12672_);
  and _21039_ (_12675_, _12674_, _08208_);
  or _21040_ (_12676_, _12675_, _08281_);
  nand _21041_ (_12677_, _08174_, _10820_);
  or _21042_ (_12678_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _21043_ (_12679_, _12678_, _12677_);
  and _21044_ (_12680_, _12679_, _08200_);
  nand _21045_ (_12681_, _08174_, _10619_);
  or _21046_ (_12682_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _21047_ (_12683_, _12682_, _12681_);
  and _21048_ (_12684_, _12683_, _08221_);
  or _21049_ (_12685_, _12684_, _12680_);
  nand _21050_ (_12686_, _08174_, _10195_);
  or _21051_ (_12687_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _21052_ (_12688_, _12687_, _12686_);
  and _21053_ (_12689_, _12688_, _08196_);
  or _21054_ (_12690_, _12689_, _12685_);
  or _21055_ (_12691_, _12690_, _12676_);
  and _21056_ (_12692_, _12691_, _12671_);
  and _21057_ (_12693_, _12692_, _08253_);
  or _21058_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12693_, _12651_);
  and _21059_ (_12695_, _08254_, word_in[3]);
  nand _21060_ (_12696_, _08174_, _09513_);
  or _21061_ (_12697_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _21062_ (_12698_, _12697_, _12696_);
  and _21063_ (_12699_, _12698_, _08208_);
  or _21064_ (_12700_, _12699_, _08184_);
  nand _21065_ (_12701_, _08174_, _09764_);
  or _21066_ (_12702_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _21067_ (_12703_, _12702_, _12701_);
  and _21068_ (_12704_, _12703_, _08221_);
  nand _21069_ (_12705_, _08174_, _09976_);
  or _21070_ (_12706_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _21071_ (_12707_, _12706_, _12705_);
  and _21072_ (_12708_, _12707_, _08200_);
  nand _21073_ (_12709_, _08174_, _09258_);
  or _21074_ (_12710_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _21075_ (_12711_, _12710_, _12709_);
  and _21076_ (_12712_, _12711_, _08196_);
  or _21077_ (_12713_, _12712_, _12708_);
  or _21078_ (_12714_, _12713_, _12704_);
  or _21079_ (_12715_, _12714_, _12700_);
  nand _21080_ (_12716_, _08174_, _10412_);
  or _21081_ (_12717_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _21082_ (_12718_, _12717_, _12716_);
  and _21083_ (_12719_, _12718_, _08208_);
  or _21084_ (_12720_, _12719_, _08281_);
  nand _21085_ (_12721_, _08174_, _10838_);
  or _21086_ (_12722_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _21087_ (_12723_, _12722_, _12721_);
  and _21088_ (_12724_, _12723_, _08200_);
  nand _21089_ (_12725_, _08174_, _10631_);
  or _21090_ (_12726_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _21091_ (_12727_, _12726_, _12725_);
  and _21092_ (_12728_, _12727_, _08221_);
  or _21093_ (_12729_, _12728_, _12724_);
  nand _21094_ (_12730_, _08174_, _10208_);
  or _21095_ (_12731_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _21096_ (_12732_, _12731_, _12730_);
  and _21097_ (_12733_, _12732_, _08196_);
  or _21098_ (_12734_, _12733_, _12729_);
  or _21099_ (_12735_, _12734_, _12720_);
  and _21100_ (_12736_, _12735_, _12715_);
  and _21101_ (_12737_, _12736_, _08253_);
  or _21102_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _12737_, _12695_);
  and _21103_ (_12738_, _08254_, word_in[4]);
  nand _21104_ (_12739_, _08174_, _09275_);
  or _21105_ (_12740_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _21106_ (_12741_, _12740_, _12739_);
  and _21107_ (_12742_, _12741_, _08196_);
  or _21108_ (_12743_, _12742_, _08184_);
  nand _21109_ (_12744_, _08174_, _09776_);
  or _21110_ (_12745_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _21111_ (_12746_, _12745_, _12744_);
  and _21112_ (_12747_, _12746_, _08221_);
  nand _21113_ (_12748_, _08174_, _09991_);
  or _21114_ (_12749_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _21115_ (_12750_, _12749_, _12748_);
  and _21116_ (_12751_, _12750_, _08200_);
  nand _21117_ (_12752_, _08174_, _09525_);
  or _21118_ (_12753_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _21119_ (_12754_, _12753_, _12752_);
  and _21120_ (_12755_, _12754_, _08208_);
  or _21121_ (_12756_, _12755_, _12751_);
  or _21122_ (_12757_, _12756_, _12747_);
  or _21123_ (_12758_, _12757_, _12743_);
  nand _21124_ (_12759_, _08174_, _10220_);
  or _21125_ (_12760_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _21126_ (_12761_, _12760_, _12759_);
  and _21127_ (_12762_, _12761_, _08196_);
  or _21128_ (_12763_, _12762_, _08281_);
  nand _21129_ (_12764_, _08174_, _10643_);
  or _21130_ (_12765_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _21131_ (_12766_, _12765_, _12764_);
  and _21132_ (_12767_, _12766_, _08221_);
  nand _21133_ (_12768_, _08174_, _10850_);
  or _21134_ (_12769_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _21135_ (_12770_, _12769_, _12768_);
  and _21136_ (_12771_, _12770_, _08200_);
  nand _21137_ (_12772_, _08174_, _10425_);
  or _21138_ (_12773_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _21139_ (_12774_, _12773_, _12772_);
  and _21140_ (_12775_, _12774_, _08208_);
  or _21141_ (_12776_, _12775_, _12771_);
  or _21142_ (_12777_, _12776_, _12767_);
  or _21143_ (_12778_, _12777_, _12763_);
  and _21144_ (_12779_, _12778_, _12758_);
  and _21145_ (_12780_, _12779_, _08253_);
  or _21146_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _12780_, _12738_);
  and _21147_ (_12781_, _08254_, word_in[5]);
  nand _21148_ (_12782_, _08174_, _09295_);
  or _21149_ (_12783_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _21150_ (_12784_, _12783_, _12782_);
  and _21151_ (_12785_, _12784_, _08196_);
  or _21152_ (_12786_, _12785_, _08184_);
  nand _21153_ (_12787_, _08174_, _09787_);
  or _21154_ (_12788_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _21155_ (_12789_, _12788_, _12787_);
  and _21156_ (_12790_, _12789_, _08221_);
  nand _21157_ (_12791_, _08174_, _10008_);
  or _21158_ (_12792_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _21159_ (_12793_, _12792_, _12791_);
  and _21160_ (_12794_, _12793_, _08200_);
  nand _21161_ (_12795_, _08174_, _09538_);
  or _21162_ (_12796_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _21163_ (_12797_, _12796_, _12795_);
  and _21164_ (_12798_, _12797_, _08208_);
  or _21165_ (_12799_, _12798_, _12794_);
  or _21166_ (_12800_, _12799_, _12790_);
  or _21167_ (_12801_, _12800_, _12786_);
  nand _21168_ (_12802_, _08174_, _10232_);
  or _21169_ (_12803_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _21170_ (_12804_, _12803_, _12802_);
  and _21171_ (_12805_, _12804_, _08196_);
  or _21172_ (_12806_, _12805_, _08281_);
  nand _21173_ (_12807_, _08174_, _10654_);
  or _21174_ (_12808_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _21175_ (_12809_, _12808_, _12807_);
  and _21176_ (_12810_, _12809_, _08221_);
  nand _21177_ (_12811_, _08174_, _10862_);
  or _21178_ (_12812_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _21179_ (_12813_, _12812_, _12811_);
  and _21180_ (_12814_, _12813_, _08200_);
  nand _21181_ (_12815_, _08174_, _10441_);
  or _21182_ (_12816_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _21183_ (_12817_, _12816_, _12815_);
  and _21184_ (_12818_, _12817_, _08208_);
  or _21185_ (_12819_, _12818_, _12814_);
  or _21186_ (_12820_, _12819_, _12810_);
  or _21187_ (_12821_, _12820_, _12806_);
  and _21188_ (_12822_, _12821_, _12801_);
  and _21189_ (_12823_, _12822_, _08253_);
  or _21190_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _12823_, _12781_);
  and _21191_ (_12824_, _08254_, word_in[6]);
  nand _21192_ (_12825_, _08174_, _09313_);
  or _21193_ (_12826_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _21194_ (_12827_, _12826_, _12825_);
  and _21195_ (_12828_, _12827_, _08196_);
  or _21196_ (_12829_, _12828_, _08184_);
  nand _21197_ (_12830_, _08174_, _09800_);
  or _21198_ (_12831_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _21199_ (_12832_, _12831_, _12830_);
  and _21200_ (_12833_, _12832_, _08221_);
  nand _21201_ (_12834_, _08174_, _10019_);
  or _21202_ (_12835_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _21203_ (_12836_, _12835_, _12834_);
  and _21204_ (_12837_, _12836_, _08200_);
  nand _21205_ (_12838_, _08174_, _09550_);
  or _21206_ (_12839_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _21207_ (_12840_, _12839_, _12838_);
  and _21208_ (_12841_, _12840_, _08208_);
  or _21209_ (_12842_, _12841_, _12837_);
  or _21210_ (_12843_, _12842_, _12833_);
  or _21211_ (_12844_, _12843_, _12829_);
  nand _21212_ (_12845_, _08174_, _10244_);
  or _21213_ (_12846_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _21214_ (_12847_, _12846_, _12845_);
  and _21215_ (_12848_, _12847_, _08196_);
  or _21216_ (_12849_, _12848_, _08281_);
  nand _21217_ (_12850_, _08174_, _10667_);
  or _21218_ (_12851_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _21219_ (_12852_, _12851_, _12850_);
  and _21220_ (_12853_, _12852_, _08221_);
  nand _21221_ (_12854_, _08174_, _10874_);
  or _21222_ (_12855_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _21223_ (_12856_, _12855_, _12854_);
  and _21224_ (_12857_, _12856_, _08200_);
  nand _21225_ (_12858_, _08174_, _10454_);
  or _21226_ (_12859_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _21227_ (_12860_, _12859_, _12858_);
  and _21228_ (_12861_, _12860_, _08208_);
  or _21229_ (_12862_, _12861_, _12857_);
  or _21230_ (_12863_, _12862_, _12853_);
  or _21231_ (_12864_, _12863_, _12849_);
  and _21232_ (_12865_, _12864_, _12844_);
  and _21233_ (_12866_, _12865_, _08253_);
  or _21234_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _12866_, _12824_);
  and _21235_ (_12867_, _08357_, word_in[8]);
  nand _21236_ (_12868_, _08174_, _09369_);
  or _21237_ (_12869_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _21238_ (_12870_, _12869_, _12868_);
  and _21239_ (_12871_, _12870_, _08359_);
  nand _21240_ (_12872_, _08174_, _09047_);
  or _21241_ (_12873_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _21242_ (_12874_, _12873_, _12872_);
  and _21243_ (_12875_, _12874_, _08358_);
  or _21244_ (_12876_, _12875_, _12871_);
  and _21245_ (_12877_, _12876_, _08321_);
  nand _21246_ (_12878_, _08174_, _10269_);
  or _21247_ (_12879_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _21248_ (_12880_, _12879_, _12878_);
  and _21249_ (_12881_, _12880_, _08359_);
  nand _21250_ (_12882_, _08174_, _10050_);
  or _21251_ (_12883_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _21252_ (_12884_, _12883_, _12882_);
  and _21253_ (_12885_, _12884_, _08358_);
  or _21254_ (_12886_, _12885_, _12881_);
  and _21255_ (_12887_, _12886_, _08323_);
  nand _21256_ (_12888_, _08174_, _09825_);
  or _21257_ (_12889_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _21258_ (_12890_, _12889_, _12888_);
  and _21259_ (_12891_, _12890_, _08359_);
  nand _21260_ (_12892_, _08174_, _09593_);
  or _21261_ (_12893_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _21262_ (_12894_, _12893_, _12892_);
  and _21263_ (_12895_, _12894_, _08358_);
  or _21264_ (_12896_, _12895_, _12891_);
  and _21265_ (_12897_, _12896_, _08346_);
  nand _21266_ (_12898_, _08174_, _10700_);
  or _21267_ (_12899_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _21268_ (_12900_, _12899_, _12898_);
  and _21269_ (_12901_, _12900_, _08359_);
  nand _21270_ (_12902_, _08174_, _10484_);
  or _21271_ (_12903_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _21272_ (_12904_, _12903_, _12902_);
  and _21273_ (_12905_, _12904_, _08358_);
  or _21274_ (_12906_, _12905_, _12901_);
  and _21275_ (_12908_, _12906_, _08350_);
  or _21276_ (_12909_, _12908_, _12897_);
  or _21277_ (_12910_, _12909_, _12887_);
  nor _21278_ (_12911_, _12910_, _12877_);
  nor _21279_ (_12912_, _12911_, _08357_);
  or _21280_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _12912_, _12867_);
  and _21281_ (_12913_, _08357_, word_in[9]);
  nand _21282_ (_12914_, _08174_, _09386_);
  or _21283_ (_12915_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _21284_ (_12916_, _12915_, _12914_);
  and _21285_ (_12918_, _12916_, _08359_);
  nand _21286_ (_12919_, _08174_, _09078_);
  or _21287_ (_12920_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _21288_ (_12921_, _12920_, _12919_);
  and _21289_ (_12922_, _12921_, _08358_);
  or _21290_ (_12923_, _12922_, _12918_);
  and _21291_ (_12924_, _12923_, _08321_);
  nand _21292_ (_12925_, _08174_, _10285_);
  or _21293_ (_12926_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _21294_ (_12927_, _12926_, _12925_);
  and _21295_ (_12928_, _12927_, _08359_);
  nand _21296_ (_12929_, _08174_, _10066_);
  or _21297_ (_12930_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _21298_ (_12931_, _12930_, _12929_);
  and _21299_ (_12932_, _12931_, _08358_);
  or _21300_ (_12933_, _12932_, _12928_);
  and _21301_ (_12934_, _12933_, _08323_);
  nand _21302_ (_12935_, _08174_, _09841_);
  or _21303_ (_12936_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _21304_ (_12937_, _12936_, _12935_);
  and _21305_ (_12938_, _12937_, _08359_);
  nand _21306_ (_12939_, _08174_, _09611_);
  or _21307_ (_12940_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _21308_ (_12941_, _12940_, _12939_);
  and _21309_ (_12942_, _12941_, _08358_);
  or _21310_ (_12943_, _12942_, _12938_);
  and _21311_ (_12944_, _12943_, _08346_);
  nand _21312_ (_12945_, _08174_, _10712_);
  or _21313_ (_12946_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _21314_ (_12947_, _12946_, _12945_);
  and _21315_ (_12948_, _12947_, _08359_);
  nand _21316_ (_12949_, _08174_, _10501_);
  or _21317_ (_12950_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _21318_ (_12951_, _12950_, _12949_);
  and _21319_ (_12952_, _12951_, _08358_);
  or _21320_ (_12953_, _12952_, _12948_);
  and _21321_ (_12954_, _12953_, _08350_);
  or _21322_ (_12955_, _12954_, _12944_);
  or _21323_ (_12956_, _12955_, _12934_);
  nor _21324_ (_12957_, _12956_, _12924_);
  nor _21325_ (_12958_, _12957_, _08357_);
  or _21326_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _12958_, _12913_);
  and _21327_ (_12959_, _08357_, word_in[10]);
  nand _21328_ (_12960_, _08174_, _09400_);
  or _21329_ (_12961_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _21330_ (_12962_, _12961_, _12960_);
  and _21331_ (_12963_, _12962_, _08359_);
  nand _21332_ (_12964_, _08174_, _09093_);
  or _21333_ (_12965_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _21334_ (_12966_, _12965_, _12964_);
  and _21335_ (_12967_, _12966_, _08358_);
  or _21336_ (_12968_, _12967_, _12963_);
  and _21337_ (_12969_, _12968_, _08321_);
  nand _21338_ (_12970_, _08174_, _10298_);
  or _21339_ (_12971_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _21340_ (_12972_, _12971_, _12970_);
  and _21341_ (_12973_, _12972_, _08359_);
  nand _21342_ (_12974_, _08174_, _10079_);
  or _21343_ (_12975_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _21344_ (_12976_, _12975_, _12974_);
  and _21345_ (_12977_, _12976_, _08358_);
  or _21346_ (_12978_, _12977_, _12973_);
  and _21347_ (_12979_, _12978_, _08323_);
  nand _21348_ (_12980_, _08174_, _09853_);
  or _21349_ (_12981_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _21350_ (_12982_, _12981_, _12980_);
  and _21351_ (_12983_, _12982_, _08359_);
  nand _21352_ (_12984_, _08174_, _09623_);
  or _21353_ (_12985_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _21354_ (_12986_, _12985_, _12984_);
  and _21355_ (_12987_, _12986_, _08358_);
  or _21356_ (_12988_, _12987_, _12983_);
  and _21357_ (_12989_, _12988_, _08346_);
  nand _21358_ (_12990_, _08174_, _10724_);
  or _21359_ (_12991_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _21360_ (_12992_, _12991_, _12990_);
  and _21361_ (_12993_, _12992_, _08359_);
  nand _21362_ (_12994_, _08174_, _10513_);
  or _21363_ (_12995_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _21364_ (_12996_, _12995_, _12994_);
  and _21365_ (_12998_, _12996_, _08358_);
  or _21366_ (_12999_, _12998_, _12993_);
  and _21367_ (_13000_, _12999_, _08350_);
  or _21368_ (_13001_, _13000_, _12989_);
  or _21369_ (_13002_, _13001_, _12979_);
  nor _21370_ (_13003_, _13002_, _12969_);
  nor _21371_ (_13004_, _13003_, _08357_);
  or _21372_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13004_, _12959_);
  and _21373_ (_13005_, _08357_, word_in[11]);
  nand _21374_ (_13006_, _08174_, _09413_);
  or _21375_ (_13007_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _21376_ (_13008_, _13007_, _13006_);
  and _21377_ (_13009_, _13008_, _08359_);
  nand _21378_ (_13010_, _08174_, _09105_);
  or _21379_ (_13011_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _21380_ (_13012_, _13011_, _13010_);
  and _21381_ (_13013_, _13012_, _08358_);
  or _21382_ (_13014_, _13013_, _13009_);
  and _21383_ (_13015_, _13014_, _08321_);
  nand _21384_ (_13016_, _08174_, _10310_);
  or _21385_ (_13017_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _21386_ (_13018_, _13017_, _13016_);
  and _21387_ (_13019_, _13018_, _08359_);
  nand _21388_ (_13020_, _08174_, _10095_);
  or _21389_ (_13021_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _21390_ (_13022_, _13021_, _13020_);
  and _21391_ (_13023_, _13022_, _08358_);
  or _21392_ (_13024_, _13023_, _13019_);
  and _21393_ (_13025_, _13024_, _08323_);
  nand _21394_ (_13026_, _08174_, _09865_);
  or _21395_ (_13027_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _21396_ (_13028_, _13027_, _13026_);
  and _21397_ (_13029_, _13028_, _08359_);
  nand _21398_ (_13030_, _08174_, _09636_);
  or _21399_ (_13031_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _21400_ (_13032_, _13031_, _13030_);
  and _21401_ (_13033_, _13032_, _08358_);
  or _21402_ (_13035_, _13033_, _13029_);
  and _21403_ (_13036_, _13035_, _08346_);
  nand _21404_ (_13037_, _08174_, _10736_);
  or _21405_ (_13038_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _21406_ (_13039_, _13038_, _13037_);
  and _21407_ (_13040_, _13039_, _08359_);
  nand _21408_ (_13041_, _08174_, _10525_);
  or _21409_ (_13042_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _21410_ (_13043_, _13042_, _13041_);
  and _21411_ (_13044_, _13043_, _08358_);
  or _21412_ (_13045_, _13044_, _13040_);
  and _21413_ (_13046_, _13045_, _08350_);
  or _21414_ (_13047_, _13046_, _13036_);
  or _21415_ (_13048_, _13047_, _13025_);
  nor _21416_ (_13049_, _13048_, _13015_);
  nor _21417_ (_13050_, _13049_, _08357_);
  or _21418_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13050_, _13005_);
  and _21419_ (_13051_, _08357_, word_in[12]);
  nand _21420_ (_13052_, _08174_, _09424_);
  or _21421_ (_13053_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _21422_ (_13054_, _13053_, _13052_);
  and _21423_ (_13055_, _13054_, _08359_);
  nand _21424_ (_13057_, _08174_, _09120_);
  or _21425_ (_13058_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _21426_ (_13059_, _13058_, _13057_);
  and _21427_ (_13060_, _13059_, _08358_);
  or _21428_ (_13061_, _13060_, _13055_);
  and _21429_ (_13062_, _13061_, _08321_);
  nand _21430_ (_13063_, _08174_, _10323_);
  or _21431_ (_13064_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _21432_ (_13065_, _13064_, _13063_);
  and _21433_ (_13066_, _13065_, _08359_);
  nand _21434_ (_13067_, _08174_, _10110_);
  or _21435_ (_13068_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _21436_ (_13069_, _13068_, _13067_);
  and _21437_ (_13070_, _13069_, _08358_);
  or _21438_ (_13071_, _13070_, _13066_);
  and _21439_ (_13072_, _13071_, _08323_);
  nand _21440_ (_13073_, _08174_, _09878_);
  or _21441_ (_13074_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _21442_ (_13075_, _13074_, _13073_);
  and _21443_ (_13076_, _13075_, _08359_);
  nand _21444_ (_13077_, _08174_, _09648_);
  or _21445_ (_13078_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _21446_ (_13079_, _13078_, _13077_);
  and _21447_ (_13080_, _13079_, _08358_);
  or _21448_ (_13081_, _13080_, _13076_);
  and _21449_ (_13082_, _13081_, _08346_);
  nand _21450_ (_13083_, _08174_, _10747_);
  or _21451_ (_13084_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _21452_ (_13086_, _13084_, _13083_);
  and _21453_ (_13087_, _13086_, _08359_);
  nand _21454_ (_13088_, _08174_, _10537_);
  or _21455_ (_13089_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _21456_ (_13090_, _13089_, _13088_);
  and _21457_ (_13091_, _13090_, _08358_);
  or _21458_ (_13092_, _13091_, _13087_);
  and _21459_ (_13093_, _13092_, _08350_);
  or _21460_ (_13094_, _13093_, _13082_);
  or _21461_ (_13095_, _13094_, _13072_);
  nor _21462_ (_13096_, _13095_, _13062_);
  nor _21463_ (_13097_, _13096_, _08357_);
  or _21464_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13097_, _13051_);
  and _21465_ (_13099_, _08357_, word_in[13]);
  nand _21466_ (_13100_, _08174_, _09435_);
  or _21467_ (_13101_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _21468_ (_13102_, _13101_, _13100_);
  and _21469_ (_13103_, _13102_, _08359_);
  nand _21470_ (_13104_, _08174_, _09131_);
  or _21471_ (_13105_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _21472_ (_13106_, _13105_, _13104_);
  and _21473_ (_13107_, _13106_, _08358_);
  or _21474_ (_13108_, _13107_, _13103_);
  and _21475_ (_13109_, _13108_, _08321_);
  nand _21476_ (_13111_, _08174_, _10334_);
  or _21477_ (_13112_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _21478_ (_13113_, _13112_, _13111_);
  and _21479_ (_13114_, _13113_, _08359_);
  nand _21480_ (_13115_, _08174_, _10121_);
  or _21481_ (_13116_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _21482_ (_13117_, _13116_, _13115_);
  and _21483_ (_13118_, _13117_, _08358_);
  or _21484_ (_13119_, _13118_, _13114_);
  and _21485_ (_13120_, _13119_, _08323_);
  nand _21486_ (_13121_, _08174_, _09891_);
  or _21487_ (_13122_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _21488_ (_13123_, _13122_, _13121_);
  and _21489_ (_13124_, _13123_, _08359_);
  nand _21490_ (_13125_, _08174_, _09661_);
  or _21491_ (_13126_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _21492_ (_13127_, _13126_, _13125_);
  and _21493_ (_13128_, _13127_, _08358_);
  or _21494_ (_13129_, _13128_, _13124_);
  and _21495_ (_13130_, _13129_, _08346_);
  nand _21496_ (_13131_, _08174_, _10761_);
  or _21497_ (_13132_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _21498_ (_13133_, _13132_, _13131_);
  and _21499_ (_13134_, _13133_, _08359_);
  nand _21500_ (_13135_, _08174_, _10549_);
  or _21501_ (_13136_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _21502_ (_13137_, _13136_, _13135_);
  and _21503_ (_13138_, _13137_, _08358_);
  or _21504_ (_13139_, _13138_, _13134_);
  and _21505_ (_13140_, _13139_, _08350_);
  or _21506_ (_13141_, _13140_, _13130_);
  or _21507_ (_13142_, _13141_, _13120_);
  nor _21508_ (_13143_, _13142_, _13109_);
  nor _21509_ (_13144_, _13143_, _08357_);
  or _21510_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13144_, _13099_);
  and _21511_ (_13145_, _08357_, word_in[14]);
  nand _21512_ (_13146_, _08174_, _09448_);
  or _21513_ (_13147_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _21514_ (_13148_, _13147_, _13146_);
  and _21515_ (_13149_, _13148_, _08359_);
  nand _21516_ (_13150_, _08174_, _09144_);
  or _21517_ (_13151_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _21518_ (_13152_, _13151_, _13150_);
  and _21519_ (_13153_, _13152_, _08358_);
  or _21520_ (_13154_, _13153_, _13149_);
  and _21521_ (_13155_, _13154_, _08321_);
  nand _21522_ (_13156_, _08174_, _10346_);
  or _21523_ (_13157_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _21524_ (_13158_, _13157_, _13156_);
  and _21525_ (_13159_, _13158_, _08359_);
  nand _21526_ (_13160_, _08174_, _10134_);
  or _21527_ (_13161_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _21528_ (_13162_, _13161_, _13160_);
  and _21529_ (_13163_, _13162_, _08358_);
  or _21530_ (_13164_, _13163_, _13159_);
  and _21531_ (_13165_, _13164_, _08323_);
  nand _21532_ (_13166_, _08174_, _09910_);
  or _21533_ (_13167_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _21534_ (_13168_, _13167_, _13166_);
  and _21535_ (_13169_, _13168_, _08359_);
  nand _21536_ (_13170_, _08174_, _09673_);
  or _21537_ (_13171_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _21538_ (_13172_, _13171_, _13170_);
  and _21539_ (_13173_, _13172_, _08358_);
  or _21540_ (_13174_, _13173_, _13169_);
  and _21541_ (_13175_, _13174_, _08346_);
  nand _21542_ (_13176_, _08174_, _10773_);
  or _21543_ (_13177_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _21544_ (_13178_, _13177_, _13176_);
  and _21545_ (_13179_, _13178_, _08359_);
  nand _21546_ (_13180_, _08174_, _10561_);
  or _21547_ (_13181_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _21548_ (_13182_, _13181_, _13180_);
  and _21549_ (_13183_, _13182_, _08358_);
  or _21550_ (_13184_, _13183_, _13179_);
  and _21551_ (_13185_, _13184_, _08350_);
  or _21552_ (_13186_, _13185_, _13175_);
  or _21553_ (_13187_, _13186_, _13165_);
  nor _21554_ (_13188_, _13187_, _13155_);
  nor _21555_ (_13189_, _13188_, _08357_);
  or _21556_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13189_, _13145_);
  and _21557_ (_13190_, _08450_, word_in[16]);
  and _21558_ (_13191_, _12579_, _08196_);
  and _21559_ (_13192_, _12566_, _08200_);
  or _21560_ (_13193_, _13192_, _13191_);
  and _21561_ (_13194_, _12575_, _08221_);
  and _21562_ (_13195_, _12571_, _08208_);
  or _21563_ (_13196_, _13195_, _13194_);
  or _21564_ (_13197_, _13196_, _13193_);
  or _21565_ (_13198_, _13197_, _08419_);
  and _21566_ (_13199_, _12595_, _08221_);
  and _21567_ (_13200_, _12599_, _08196_);
  or _21568_ (_13201_, _13200_, _13199_);
  and _21569_ (_13202_, _12591_, _08208_);
  and _21570_ (_13203_, _12586_, _08200_);
  or _21571_ (_13204_, _13203_, _13202_);
  or _21572_ (_13205_, _13204_, _13201_);
  or _21573_ (_13207_, _13205_, _08460_);
  nand _21574_ (_13208_, _13207_, _13198_);
  nor _21575_ (_13209_, _13208_, _08450_);
  or _21576_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13209_, _13190_);
  and _21577_ (_13210_, _08450_, word_in[17]);
  and _21578_ (_13211_, _12623_, _08200_);
  and _21579_ (_13212_, _12610_, _08196_);
  or _21580_ (_13213_, _13212_, _13211_);
  and _21581_ (_13214_, _12615_, _08208_);
  and _21582_ (_13215_, _12619_, _08221_);
  or _21583_ (_13216_, _13215_, _13214_);
  or _21584_ (_13217_, _13216_, _13213_);
  or _21585_ (_13218_, _13217_, _08419_);
  and _21586_ (_13219_, _12636_, _08221_);
  and _21587_ (_13220_, _12631_, _08196_);
  or _21588_ (_13221_, _13220_, _13219_);
  and _21589_ (_13222_, _12640_, _08208_);
  and _21590_ (_13223_, _12645_, _08200_);
  or _21591_ (_13224_, _13223_, _13222_);
  or _21592_ (_13225_, _13224_, _13221_);
  or _21593_ (_13226_, _13225_, _08460_);
  nand _21594_ (_13227_, _13226_, _13218_);
  nor _21595_ (_13228_, _13227_, _08450_);
  or _21596_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13228_, _13210_);
  and _21597_ (_13229_, _08450_, word_in[18]);
  and _21598_ (_13230_, _12663_, _08221_);
  and _21599_ (_13231_, _12654_, _08196_);
  or _21600_ (_13232_, _13231_, _13230_);
  and _21601_ (_13233_, _12659_, _08208_);
  and _21602_ (_13234_, _12667_, _08200_);
  or _21603_ (_13235_, _13234_, _13233_);
  or _21604_ (_13236_, _13235_, _13232_);
  or _21605_ (_13237_, _13236_, _08419_);
  and _21606_ (_13238_, _12674_, _08196_);
  and _21607_ (_13239_, _12688_, _08200_);
  or _21608_ (_13240_, _13239_, _13238_);
  and _21609_ (_13241_, _12679_, _08221_);
  and _21610_ (_13242_, _12683_, _08208_);
  or _21611_ (_13243_, _13242_, _13241_);
  or _21612_ (_13244_, _13243_, _13240_);
  or _21613_ (_13245_, _13244_, _08460_);
  nand _21614_ (_13247_, _13245_, _13237_);
  nor _21615_ (_13248_, _13247_, _08450_);
  or _21616_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13248_, _13229_);
  and _21617_ (_13249_, _08450_, word_in[19]);
  and _21618_ (_13250_, _12707_, _08221_);
  and _21619_ (_13251_, _12698_, _08196_);
  or _21620_ (_13252_, _13251_, _13250_);
  and _21621_ (_13253_, _12703_, _08208_);
  and _21622_ (_13254_, _12711_, _08200_);
  or _21623_ (_13255_, _13254_, _13253_);
  or _21624_ (_13256_, _13255_, _13252_);
  or _21625_ (_13257_, _13256_, _08419_);
  and _21626_ (_13258_, _12723_, _08221_);
  and _21627_ (_13259_, _12718_, _08196_);
  or _21628_ (_13260_, _13259_, _13258_);
  and _21629_ (_13261_, _12727_, _08208_);
  and _21630_ (_13262_, _12732_, _08200_);
  or _21631_ (_13263_, _13262_, _13261_);
  or _21632_ (_13264_, _13263_, _13260_);
  or _21633_ (_13265_, _13264_, _08460_);
  nand _21634_ (_13266_, _13265_, _13257_);
  nor _21635_ (_13267_, _13266_, _08450_);
  or _21636_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13267_, _13249_);
  and _21637_ (_13268_, _08450_, word_in[20]);
  and _21638_ (_13269_, _12750_, _08221_);
  and _21639_ (_13270_, _12754_, _08196_);
  or _21640_ (_13271_, _13270_, _13269_);
  and _21641_ (_13272_, _12746_, _08208_);
  and _21642_ (_13273_, _12741_, _08200_);
  or _21643_ (_13274_, _13273_, _13272_);
  or _21644_ (_13275_, _13274_, _13271_);
  or _21645_ (_13276_, _13275_, _08419_);
  and _21646_ (_13277_, _12770_, _08221_);
  and _21647_ (_13278_, _12774_, _08196_);
  or _21648_ (_13279_, _13278_, _13277_);
  and _21649_ (_13280_, _12766_, _08208_);
  and _21650_ (_13282_, _12761_, _08200_);
  or _21651_ (_13283_, _13282_, _13280_);
  or _21652_ (_13284_, _13283_, _13279_);
  or _21653_ (_13285_, _13284_, _08460_);
  nand _21654_ (_13286_, _13285_, _13276_);
  nor _21655_ (_13287_, _13286_, _08450_);
  or _21656_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13287_, _13268_);
  and _21657_ (_13288_, _08450_, word_in[21]);
  and _21658_ (_13290_, _12793_, _08221_);
  and _21659_ (_13291_, _12797_, _08196_);
  or _21660_ (_13292_, _13291_, _13290_);
  and _21661_ (_13293_, _12789_, _08208_);
  and _21662_ (_13294_, _12784_, _08200_);
  or _21663_ (_13295_, _13294_, _13293_);
  or _21664_ (_13296_, _13295_, _13292_);
  or _21665_ (_13297_, _13296_, _08419_);
  and _21666_ (_13298_, _12817_, _08196_);
  and _21667_ (_13299_, _12804_, _08200_);
  or _21668_ (_13300_, _13299_, _13298_);
  and _21669_ (_13301_, _12813_, _08221_);
  and _21670_ (_13302_, _12809_, _08208_);
  or _21671_ (_13303_, _13302_, _13301_);
  or _21672_ (_13304_, _13303_, _13300_);
  or _21673_ (_13305_, _13304_, _08460_);
  nand _21674_ (_13306_, _13305_, _13297_);
  nor _21675_ (_13307_, _13306_, _08450_);
  or _21676_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13307_, _13288_);
  and _21677_ (_13308_, _08450_, word_in[22]);
  and _21678_ (_13309_, _12836_, _08221_);
  and _21679_ (_13310_, _12840_, _08196_);
  or _21680_ (_13311_, _13310_, _13309_);
  and _21681_ (_13312_, _12832_, _08208_);
  and _21682_ (_13313_, _12827_, _08200_);
  or _21683_ (_13314_, _13313_, _13312_);
  or _21684_ (_13315_, _13314_, _13311_);
  or _21685_ (_13316_, _13315_, _08419_);
  and _21686_ (_13317_, _12860_, _08196_);
  and _21687_ (_13318_, _12847_, _08200_);
  or _21688_ (_13319_, _13318_, _13317_);
  and _21689_ (_13320_, _12856_, _08221_);
  and _21690_ (_13321_, _12852_, _08208_);
  or _21691_ (_13322_, _13321_, _13320_);
  or _21692_ (_13323_, _13322_, _13319_);
  or _21693_ (_13325_, _13323_, _08460_);
  nand _21694_ (_13326_, _13325_, _13316_);
  nor _21695_ (_13327_, _13326_, _08450_);
  or _21696_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13327_, _13308_);
  or _21697_ (_13329_, _11830_, _08748_);
  and _21698_ (_13330_, _13329_, _11889_);
  and _21699_ (_13331_, _11830_, _11395_);
  and _21700_ (_13332_, _11852_, _11415_);
  or _21701_ (_13333_, _13332_, _13331_);
  or _21702_ (_13334_, _13333_, _13330_);
  and _21703_ (_13335_, _11810_, _08750_);
  and _21704_ (_13337_, _11867_, _11415_);
  or _21705_ (_13338_, _13337_, _13335_);
  and _21706_ (_13339_, _11737_, _11810_);
  and _21707_ (_13340_, _11805_, _11415_);
  or _21708_ (_13341_, _13340_, _13339_);
  or _21709_ (_13342_, _13341_, _13338_);
  or _21710_ (_13343_, _13342_, _13334_);
  and _21711_ (_13344_, _11404_, _08757_);
  and _21712_ (_13345_, _11400_, _08757_);
  or _21713_ (_13346_, _13345_, _13344_);
  or _21714_ (_13347_, _13346_, _12536_);
  or _21715_ (_13348_, _13347_, _13343_);
  nor _21716_ (_13349_, _11878_, _08715_);
  and _21717_ (_13350_, _11404_, _11395_);
  and _21718_ (_13351_, _11391_, _08758_);
  and _21719_ (_13352_, _13351_, _08736_);
  or _21720_ (_13353_, _13352_, _13350_);
  or _21721_ (_13354_, _11410_, _11400_);
  and _21722_ (_13355_, _13354_, _11810_);
  or _21723_ (_13356_, _13355_, _13353_);
  or _21724_ (_13357_, _13356_, _13349_);
  or _21725_ (_13358_, _11921_, _11887_);
  and _21726_ (_13360_, _11415_, _11404_);
  or _21727_ (_13361_, _13360_, _12549_);
  or _21728_ (_13362_, _13361_, _13358_);
  or _21729_ (_13364_, _11918_, _11909_);
  or _21730_ (_13365_, _13364_, _11803_);
  or _21731_ (_13367_, _13365_, _13362_);
  or _21732_ (_13368_, _13367_, _13357_);
  or _21733_ (_13370_, _13368_, _13348_);
  and _21734_ (_13372_, _13370_, _06527_);
  and _21735_ (_13373_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _21736_ (_13375_, _08732_, _11390_);
  and _21737_ (_13376_, _13375_, _08749_);
  and _21738_ (_13377_, _13376_, _08754_);
  and _21739_ (_13378_, _08741_, _08736_);
  and _21740_ (_13379_, _13378_, _08746_);
  and _21741_ (_13380_, _13379_, _08757_);
  or _21742_ (_13381_, _13380_, _08767_);
  or _21743_ (_13382_, _13381_, _13377_);
  not _21744_ (_13383_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _21745_ (_13384_, _11795_, _13383_);
  and _21746_ (_13385_, _13384_, _13382_);
  or _21747_ (_13386_, _13385_, _13373_);
  or _21748_ (_13387_, _13386_, _13372_);
  and _21749_ (_11599_, _13387_, _06071_);
  and _21750_ (_13389_, _08508_, word_in[24]);
  and _21751_ (_13390_, _12884_, _08359_);
  and _21752_ (_13391_, _12880_, _08358_);
  or _21753_ (_13393_, _13391_, _13390_);
  and _21754_ (_13394_, _13393_, _08482_);
  and _21755_ (_13395_, _12874_, _08359_);
  and _21756_ (_13396_, _12870_, _08358_);
  or _21757_ (_13397_, _13396_, _13395_);
  and _21758_ (_13398_, _13397_, _08480_);
  and _21759_ (_13399_, _12894_, _08359_);
  and _21760_ (_13400_, _12890_, _08358_);
  or _21761_ (_13401_, _13400_, _13399_);
  and _21762_ (_13402_, _13401_, _08517_);
  and _21763_ (_13403_, _12904_, _08359_);
  and _21764_ (_13404_, _12900_, _08358_);
  or _21765_ (_13405_, _13404_, _13403_);
  and _21766_ (_13406_, _13405_, _08522_);
  or _21767_ (_13407_, _13406_, _13402_);
  or _21768_ (_13408_, _13407_, _13398_);
  nor _21769_ (_13409_, _13408_, _13394_);
  nor _21770_ (_13410_, _13409_, _08508_);
  or _21771_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13410_, _13389_);
  and _21772_ (_13411_, _08508_, word_in[25]);
  and _21773_ (_13412_, _12931_, _08359_);
  and _21774_ (_13414_, _12927_, _08358_);
  or _21775_ (_13415_, _13414_, _13412_);
  and _21776_ (_13417_, _13415_, _08482_);
  and _21777_ (_13418_, _12921_, _08359_);
  and _21778_ (_13419_, _12916_, _08358_);
  or _21779_ (_13420_, _13419_, _13418_);
  and _21780_ (_13421_, _13420_, _08480_);
  and _21781_ (_13422_, _12941_, _08359_);
  and _21782_ (_13423_, _12937_, _08358_);
  or _21783_ (_13425_, _13423_, _13422_);
  and _21784_ (_13426_, _13425_, _08517_);
  and _21785_ (_13428_, _12951_, _08359_);
  and _21786_ (_13429_, _12947_, _08358_);
  or _21787_ (_13431_, _13429_, _13428_);
  and _21788_ (_13432_, _13431_, _08522_);
  or _21789_ (_13434_, _13432_, _13426_);
  or _21790_ (_13435_, _13434_, _13421_);
  nor _21791_ (_13437_, _13435_, _13417_);
  nor _21792_ (_13438_, _13437_, _08508_);
  or _21793_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13438_, _13411_);
  and _21794_ (_13440_, _08508_, word_in[26]);
  and _21795_ (_13442_, _12966_, _08359_);
  and _21796_ (_13443_, _12962_, _08358_);
  or _21797_ (_13444_, _13443_, _13442_);
  and _21798_ (_13445_, _13444_, _08480_);
  and _21799_ (_13446_, _12976_, _08359_);
  and _21800_ (_13447_, _12972_, _08358_);
  or _21801_ (_13448_, _13447_, _13446_);
  and _21802_ (_13449_, _13448_, _08482_);
  and _21803_ (_13450_, _12986_, _08359_);
  and _21804_ (_13451_, _12982_, _08358_);
  or _21805_ (_13452_, _13451_, _13450_);
  and _21806_ (_13453_, _13452_, _08517_);
  and _21807_ (_13454_, _12996_, _08359_);
  and _21808_ (_13455_, _12992_, _08358_);
  or _21809_ (_13456_, _13455_, _13454_);
  and _21810_ (_13458_, _13456_, _08522_);
  or _21811_ (_13459_, _13458_, _13453_);
  or _21812_ (_13460_, _13459_, _13449_);
  nor _21813_ (_13462_, _13460_, _13445_);
  nor _21814_ (_13463_, _13462_, _08508_);
  or _21815_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13463_, _13440_);
  and _21816_ (_13465_, _08508_, word_in[27]);
  and _21817_ (_13466_, _13012_, _08359_);
  and _21818_ (_13467_, _13008_, _08358_);
  or _21819_ (_13468_, _13467_, _13466_);
  and _21820_ (_13469_, _13468_, _08480_);
  and _21821_ (_13470_, _13022_, _08359_);
  and _21822_ (_13471_, _13018_, _08358_);
  or _21823_ (_13472_, _13471_, _13470_);
  and _21824_ (_13473_, _13472_, _08482_);
  and _21825_ (_13474_, _13032_, _08359_);
  and _21826_ (_13476_, _13028_, _08358_);
  or _21827_ (_13477_, _13476_, _13474_);
  and _21828_ (_13479_, _13477_, _08517_);
  and _21829_ (_13480_, _13043_, _08359_);
  and _21830_ (_13481_, _13039_, _08358_);
  or _21831_ (_13482_, _13481_, _13480_);
  and _21832_ (_13483_, _13482_, _08522_);
  or _21833_ (_13484_, _13483_, _13479_);
  or _21834_ (_13485_, _13484_, _13473_);
  nor _21835_ (_13486_, _13485_, _13469_);
  nor _21836_ (_13488_, _13486_, _08508_);
  or _21837_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13488_, _13465_);
  and _21838_ (_13489_, _08508_, word_in[28]);
  and _21839_ (_13490_, _13069_, _08359_);
  and _21840_ (_13491_, _13065_, _08358_);
  or _21841_ (_13492_, _13491_, _13490_);
  and _21842_ (_13493_, _13492_, _08482_);
  and _21843_ (_13494_, _13059_, _08359_);
  and _21844_ (_13495_, _13054_, _08358_);
  or _21845_ (_13496_, _13495_, _13494_);
  and _21846_ (_13498_, _13496_, _08480_);
  and _21847_ (_13499_, _13079_, _08359_);
  and _21848_ (_13500_, _13075_, _08358_);
  or _21849_ (_13501_, _13500_, _13499_);
  and _21850_ (_13503_, _13501_, _08517_);
  and _21851_ (_13504_, _13090_, _08359_);
  and _21852_ (_13506_, _13086_, _08358_);
  or _21853_ (_13507_, _13506_, _13504_);
  and _21854_ (_13509_, _13507_, _08522_);
  or _21855_ (_13510_, _13509_, _13503_);
  or _21856_ (_13511_, _13510_, _13498_);
  nor _21857_ (_13512_, _13511_, _13493_);
  nor _21858_ (_13513_, _13512_, _08508_);
  or _21859_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13513_, _13489_);
  and _21860_ (_13514_, _08508_, word_in[29]);
  and _21861_ (_13515_, _13117_, _08359_);
  and _21862_ (_13516_, _13113_, _08358_);
  or _21863_ (_13518_, _13516_, _13515_);
  and _21864_ (_13519_, _13518_, _08482_);
  and _21865_ (_13521_, _13106_, _08359_);
  and _21866_ (_13522_, _13102_, _08358_);
  or _21867_ (_13523_, _13522_, _13521_);
  and _21868_ (_13524_, _13523_, _08480_);
  and _21869_ (_13525_, _13127_, _08359_);
  and _21870_ (_13526_, _13123_, _08358_);
  or _21871_ (_13527_, _13526_, _13525_);
  and _21872_ (_13528_, _13527_, _08517_);
  and _21873_ (_13529_, _13137_, _08359_);
  and _21874_ (_13530_, _13133_, _08358_);
  or _21875_ (_13531_, _13530_, _13529_);
  and _21876_ (_13532_, _13531_, _08522_);
  or _21877_ (_13533_, _13532_, _13528_);
  or _21878_ (_13534_, _13533_, _13524_);
  nor _21879_ (_13535_, _13534_, _13519_);
  nor _21880_ (_13537_, _13535_, _08508_);
  or _21881_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13537_, _13514_);
  and _21882_ (_13538_, _08508_, word_in[30]);
  and _21883_ (_13539_, _13162_, _08359_);
  and _21884_ (_13540_, _13158_, _08358_);
  or _21885_ (_13541_, _13540_, _13539_);
  and _21886_ (_13543_, _13541_, _08482_);
  and _21887_ (_13544_, _13152_, _08359_);
  and _21888_ (_13546_, _13148_, _08358_);
  or _21889_ (_13547_, _13546_, _13544_);
  and _21890_ (_13549_, _13547_, _08480_);
  and _21891_ (_13550_, _13172_, _08359_);
  and _21892_ (_13551_, _13168_, _08358_);
  or _21893_ (_13552_, _13551_, _13550_);
  and _21894_ (_13553_, _13552_, _08517_);
  and _21895_ (_13554_, _13182_, _08359_);
  and _21896_ (_13555_, _13178_, _08358_);
  or _21897_ (_13556_, _13555_, _13554_);
  and _21898_ (_13557_, _13556_, _08522_);
  or _21899_ (_13558_, _13557_, _13553_);
  or _21900_ (_13559_, _13558_, _13549_);
  nor _21901_ (_13560_, _13559_, _13543_);
  nor _21902_ (_13562_, _13560_, _08508_);
  or _21903_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13562_, _13538_);
  and _21904_ (_13564_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08003_);
  and _21905_ (_13566_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21906_ (_13567_, _13566_, _13564_);
  and _21907_ (_11677_, _13567_, _06071_);
  nor _21908_ (_11692_, _11627_, rst);
  nor _21909_ (_11712_, _11688_, rst);
  or _21910_ (_13569_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _21911_ (_13570_, _06530_, _05760_);
  and _21912_ (_13572_, _13570_, _06071_);
  and _21913_ (_11720_, _13572_, _13569_);
  nand _21914_ (_13574_, _06376_, _06386_);
  or _21915_ (_13576_, _09347_, _13574_);
  and _21916_ (_13577_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _21917_ (_13578_, _07978_, _06966_);
  or _21918_ (_13579_, _06391_, _06381_);
  and _21919_ (_13580_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _21920_ (_13582_, _13580_, _13579_);
  or _21921_ (_13583_, _13582_, _13578_);
  or _21922_ (_13584_, _13583_, _13577_);
  and _21923_ (_11767_, _13584_, _06071_);
  or _21924_ (_13585_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand _21925_ (_13586_, _06530_, _05862_);
  and _21926_ (_13587_, _13586_, _06071_);
  and _21927_ (_11809_, _13587_, _13585_);
  and _21928_ (_13588_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _21929_ (_13589_, _12197_, _06369_);
  or _21930_ (_13590_, _13589_, _13588_);
  and _21931_ (_11820_, _13590_, _06071_);
  nor _21932_ (_13592_, _11242_, _11240_);
  nor _21933_ (_13593_, _13592_, _11243_);
  or _21934_ (_13594_, _13593_, _09711_);
  or _21935_ (_13595_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _21936_ (_13597_, _13595_, _11270_);
  and _21937_ (_13598_, _13597_, _13594_);
  and _21938_ (_13599_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _21939_ (_11832_, _13599_, _13598_);
  nor _21940_ (_11871_, _11607_, rst);
  nand _21941_ (_13602_, _10978_, _08053_);
  or _21942_ (_13603_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _21943_ (_13604_, _13603_, _06071_);
  and _21944_ (_11886_, _13604_, _13602_);
  and _21945_ (_13606_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _21946_ (_13608_, _12120_, _07979_);
  or _21947_ (_13609_, _13608_, _13606_);
  and _21948_ (_11892_, _13609_, _06071_);
  or _21949_ (_13611_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand _21950_ (_13613_, _06530_, _05782_);
  and _21951_ (_13614_, _13613_, _06071_);
  and _21952_ (_11898_, _13614_, _13611_);
  and _21953_ (_13616_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _21954_ (_13617_, _11239_, _11237_);
  nor _21955_ (_13618_, _13617_, _11240_);
  or _21956_ (_13619_, _13618_, _09711_);
  or _21957_ (_13620_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _21958_ (_13621_, _13620_, _11270_);
  and _21959_ (_13623_, _13621_, _13619_);
  or _21960_ (_11941_, _13623_, _13616_);
  and _21961_ (_13625_, _11422_, _11401_);
  and _21962_ (_13627_, _11745_, _08732_);
  or _21963_ (_13628_, _13627_, _13625_);
  and _21964_ (_13629_, _11396_, _08748_);
  or _21965_ (_13630_, _13629_, _11875_);
  and _21966_ (_13631_, _11860_, _08764_);
  or _21967_ (_13632_, _11408_, _11400_);
  and _21968_ (_13633_, _13632_, _11395_);
  or _21969_ (_13634_, _13633_, _13631_);
  or _21970_ (_13635_, _13634_, _13630_);
  or _21971_ (_13636_, _13635_, _13628_);
  and _21972_ (_13637_, _13636_, _11421_);
  and _21973_ (_13638_, _13628_, _11385_);
  and _21974_ (_13639_, _13379_, _08764_);
  and _21975_ (_13640_, _13639_, _11810_);
  or _21976_ (_13641_, _13640_, _11811_);
  and _21977_ (_13642_, _13641_, _13384_);
  or _21978_ (_13643_, _13642_, _13638_);
  or _21979_ (_13644_, _13643_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _21980_ (_13645_, _13644_, _13637_);
  or _21981_ (_13646_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05686_);
  and _21982_ (_13647_, _13646_, _06071_);
  and _21983_ (_11988_, _13647_, _13645_);
  and _21984_ (_13648_, _12161_, _06369_);
  not _21985_ (_13649_, _06376_);
  or _21986_ (_13650_, _06394_, _13649_);
  nor _21987_ (_13651_, _06387_, _06390_);
  or _21988_ (_13652_, _13651_, _13650_);
  and _21989_ (_13653_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or _21990_ (_13654_, _13653_, _13648_);
  and _21991_ (_12012_, _13654_, _06071_);
  and _21992_ (_13655_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _21993_ (_13656_, _11023_, _06369_);
  or _21994_ (_13657_, _13656_, _13655_);
  and _21995_ (_12018_, _13657_, _06071_);
  and _21996_ (_13658_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _21997_ (_13659_, _06611_, _06434_);
  or _21998_ (_13660_, _13659_, _13658_);
  and _21999_ (_12048_, _13660_, _06071_);
  or _22000_ (_13661_, _11254_, _11249_);
  nor _22001_ (_13662_, _11255_, _09711_);
  and _22002_ (_13663_, _13662_, _13661_);
  nor _22003_ (_13664_, _09710_, _06153_);
  nor _22004_ (_13665_, _13664_, _13663_);
  or _22005_ (_13666_, _13665_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand _22006_ (_13667_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _22007_ (_13668_, _13667_, _13666_);
  nor _22008_ (_12089_, _13668_, rst);
  and _22009_ (_13669_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _22010_ (_13670_, _11023_, _06966_);
  and _22011_ (_13671_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _22012_ (_13672_, _13671_, _13579_);
  or _22013_ (_13673_, _13672_, _13670_);
  or _22014_ (_13674_, _13673_, _13669_);
  and _22015_ (_12099_, _13674_, _06071_);
  and _22016_ (_13675_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _22017_ (_13676_, _07945_, _06967_);
  and _22018_ (_13677_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _22019_ (_13678_, _13677_, _13579_);
  or _22020_ (_13679_, _13678_, _13676_);
  or _22021_ (_13680_, _13679_, _13675_);
  and _22022_ (_12101_, _13680_, _06071_);
  and _22023_ (_13681_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _22024_ (_13682_, _11260_, _11258_);
  nor _22025_ (_13683_, _13682_, _11261_);
  or _22026_ (_13684_, _13683_, _09711_);
  or _22027_ (_13685_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _22028_ (_13687_, _13685_, _11270_);
  and _22029_ (_13688_, _13687_, _13684_);
  or _22030_ (_12111_, _13688_, _13681_);
  nor _22031_ (_13689_, _11257_, _11084_);
  nor _22032_ (_13690_, _13689_, _11258_);
  or _22033_ (_13691_, _13690_, _09711_);
  or _22034_ (_13692_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _22035_ (_13693_, _13692_, _11270_);
  and _22036_ (_13694_, _13693_, _13691_);
  and _22037_ (_13695_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _22038_ (_12141_, _13695_, _13694_);
  and _22039_ (_12170_, _08753_, _06071_);
  and _22040_ (_13696_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _22041_ (_13697_, _11256_, _11087_);
  nor _22042_ (_13698_, _13697_, _11257_);
  or _22043_ (_13699_, _13698_, _09711_);
  or _22044_ (_13700_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _22045_ (_13701_, _13700_, _11270_);
  and _22046_ (_13702_, _13701_, _13699_);
  or _22047_ (_12175_, _13702_, _13696_);
  nor _22048_ (_12179_, _11493_, rst);
  not _22049_ (_13703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _22050_ (_13704_, _13703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _22051_ (_13705_, _13704_, _07885_);
  nor _22052_ (_13706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _22053_ (_13707_, _13706_, _13705_);
  or _22054_ (_13708_, _13707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _22055_ (_13709_, _06026_, _05923_);
  and _22056_ (_13710_, _13709_, _10946_);
  and _22057_ (_13711_, _13710_, _06806_);
  or _22058_ (_13712_, _13711_, _13708_);
  and _22059_ (_13713_, _08799_, _06383_);
  or _22060_ (_13714_, _06383_, _07907_);
  nand _22061_ (_13715_, _13714_, _13711_);
  or _22062_ (_13716_, _13715_, _13713_);
  and _22063_ (_13717_, _13716_, _13712_);
  and _22064_ (_13718_, _09248_, _06821_);
  or _22065_ (_13719_, _13718_, _13717_);
  nand _22066_ (_13720_, _13718_, _07977_);
  and _22067_ (_13721_, _13720_, _06071_);
  and _22068_ (_12181_, _13721_, _13719_);
  and _22069_ (_13722_, _07104_, _06805_);
  and _22070_ (_13723_, _13722_, _06840_);
  nand _22071_ (_13724_, _13723_, _09341_);
  or _22072_ (_13725_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _22073_ (_13726_, _13725_, _06071_);
  and _22074_ (_12190_, _13726_, _13724_);
  nand _22075_ (_13727_, _13723_, _09037_);
  or _22076_ (_13728_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _22077_ (_13729_, _13728_, _06071_);
  and _22078_ (_12193_, _13729_, _13727_);
  and _22079_ (_13730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _22080_ (_13731_, _13730_, _07885_);
  and _22081_ (_13732_, _07902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _22082_ (_13733_, _13732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22083_ (_13734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _22084_ (_13735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _22085_ (_13736_, _13735_, _13734_);
  and _22086_ (_13737_, _13736_, _13733_);
  nor _22087_ (_13738_, _13737_, _13731_);
  and _22088_ (_13739_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  not _22089_ (_13740_, _13738_);
  and _22090_ (_13741_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or _22091_ (_13742_, _13741_, _13739_);
  and _22092_ (_13743_, _06380_, _06012_);
  and _22093_ (_13744_, _13743_, _06821_);
  or _22094_ (_13745_, _13744_, _13742_);
  not _22095_ (_13746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand _22096_ (_13747_, _13746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _22097_ (_13748_, _13747_, _07902_);
  nand _22098_ (_13749_, _13748_, _13744_);
  and _22099_ (_13750_, _13749_, _13745_);
  and _22100_ (_12200_, _13750_, _06071_);
  and _22101_ (_13751_, _06362_, _06027_);
  and _22102_ (_13752_, _13751_, _06821_);
  and _22103_ (_13753_, _13752_, _07885_);
  and _22104_ (_13754_, _13753_, _12019_);
  and _22105_ (_13755_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _22106_ (_13756_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _22107_ (_13757_, _13756_, _13755_);
  nor _22108_ (_13758_, _13757_, _13744_);
  and _22109_ (_13759_, _13752_, _07902_);
  not _22110_ (_13760_, _13759_);
  nor _22111_ (_13761_, _13760_, _06434_);
  or _22112_ (_13762_, _13761_, _13758_);
  or _22113_ (_13763_, _13762_, _13754_);
  and _22114_ (_12203_, _13763_, _06071_);
  or _22115_ (_13764_, _13737_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not _22116_ (_13765_, _13731_);
  not _22117_ (_13766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand _22118_ (_13767_, _13737_, _13766_);
  and _22119_ (_13769_, _13767_, _13765_);
  and _22120_ (_13770_, _13769_, _13764_);
  nor _22121_ (_13771_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _22122_ (_13772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _22123_ (_13774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _22124_ (_13776_, _13774_, _13772_);
  and _22125_ (_13777_, _13776_, _13771_);
  not _22126_ (_13778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor _22127_ (_13779_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _22128_ (_13780_, _13779_, _13778_);
  and _22129_ (_13781_, _13780_, _13766_);
  and _22130_ (_13782_, _13781_, _13777_);
  nor _22131_ (_13783_, _13782_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _22132_ (_13784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _22133_ (_13785_, _13784_, _13783_);
  and _22134_ (_13786_, _13785_, _13731_);
  nor _22135_ (_13788_, _13786_, _13770_);
  nor _22136_ (_13789_, _13788_, _13752_);
  and _22137_ (_13790_, _13753_, _07978_);
  or _22138_ (_13791_, _13790_, _13789_);
  and _22139_ (_12206_, _13791_, _06071_);
  and _22140_ (_13792_, _13733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _22141_ (_13793_, _13792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _22142_ (_13794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _22143_ (_13796_, _13794_, _13733_);
  nor _22144_ (_13797_, _13796_, _13793_);
  nor _22145_ (_13798_, _13752_, rst);
  and _22146_ (_12211_, _13798_, _13797_);
  or _22147_ (_13799_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _22148_ (_13800_, _06530_, _05716_);
  and _22149_ (_13802_, _13800_, _06071_);
  and _22150_ (_12214_, _13802_, _13799_);
  and _22151_ (_13803_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _22152_ (_13804_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _22153_ (_13805_, _13804_, _13803_);
  and _22154_ (_12217_, _13805_, _06071_);
  nor _22155_ (_13806_, _11255_, _11091_);
  nor _22156_ (_13807_, _13806_, _11256_);
  or _22157_ (_13808_, _13807_, _09711_);
  or _22158_ (_13809_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _22159_ (_13810_, _13809_, _11270_);
  and _22160_ (_13811_, _13810_, _13808_);
  and _22161_ (_13812_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _22162_ (_12220_, _13812_, _13811_);
  not _22163_ (_13813_, _12167_);
  nor _22164_ (_13814_, _12126_, _13813_);
  not _22165_ (_13815_, _12084_);
  and _22166_ (_13816_, _13815_, _12221_);
  and _22167_ (_13817_, _13816_, _13814_);
  and _22168_ (_13818_, _12386_, _12341_);
  not _22169_ (_13819_, _12030_);
  and _22170_ (_13820_, _12426_, _13819_);
  and _22171_ (_13821_, _13820_, _13818_);
  and _22172_ (_13822_, _13821_, _13817_);
  nor _22173_ (_13823_, _12426_, _12030_);
  and _22174_ (_13824_, _13823_, _13818_);
  and _22175_ (_13825_, _13824_, _13817_);
  nor _22176_ (_13826_, _13825_, _13822_);
  not _22177_ (_13827_, _12341_);
  and _22178_ (_13828_, _12386_, _13827_);
  and _22179_ (_13829_, _13828_, _13823_);
  and _22180_ (_13830_, _13829_, _13817_);
  nor _22181_ (_13831_, _12386_, _13827_);
  and _22182_ (_13832_, _13820_, _13831_);
  and _22183_ (_13833_, _13832_, _13817_);
  nor _22184_ (_13835_, _13833_, _13830_);
  and _22185_ (_13836_, _13835_, _13826_);
  and _22186_ (_13837_, _12126_, _13815_);
  and _22187_ (_13838_, _12221_, _12167_);
  and _22188_ (_13839_, _13838_, _13837_);
  and _22189_ (_13840_, _13821_, _13839_);
  nor _22190_ (_13842_, _12386_, _12341_);
  and _22191_ (_13843_, _13842_, _13820_);
  and _22192_ (_13844_, _13843_, _13817_);
  nor _22193_ (_13845_, _13844_, _13840_);
  not _22194_ (_13846_, _12221_);
  and _22195_ (_13847_, _13837_, _13813_);
  and _22196_ (_13848_, _13847_, _13846_);
  not _22197_ (_13849_, _12426_);
  and _22198_ (_13850_, _13842_, _13849_);
  and _22199_ (_13851_, _13850_, _12030_);
  and _22200_ (_13852_, _13851_, _13848_);
  and _22201_ (_13853_, _13847_, _12221_);
  and _22202_ (_13854_, _13853_, _13821_);
  nor _22203_ (_13856_, _13854_, _13852_);
  and _22204_ (_13857_, _13856_, _13845_);
  and _22205_ (_13858_, _13857_, _13836_);
  and _22206_ (_13860_, _13843_, _13839_);
  and _22207_ (_13861_, _13828_, _13820_);
  and _22208_ (_13863_, _13861_, _13839_);
  nor _22209_ (_13864_, _13863_, _13860_);
  and _22210_ (_13865_, _13832_, _13839_);
  and _22211_ (_13866_, _13829_, _13839_);
  nor _22212_ (_13867_, _13866_, _13865_);
  and _22213_ (_13869_, _13867_, _13864_);
  and _22214_ (_13870_, _13824_, _13839_);
  and _22215_ (_13871_, _13851_, _13839_);
  nor _22216_ (_13872_, _13871_, _13870_);
  nor _22217_ (_13873_, _12221_, _13813_);
  and _22218_ (_13874_, _13873_, _13837_);
  and _22219_ (_13875_, _13874_, _13821_);
  and _22220_ (_13876_, _13861_, _13874_);
  nor _22221_ (_13877_, _13876_, _13875_);
  and _22222_ (_13878_, _13877_, _13872_);
  and _22223_ (_13879_, _13878_, _13869_);
  and _22224_ (_13880_, _13879_, _13858_);
  and _22225_ (_13881_, _12426_, _12030_);
  and _22226_ (_13882_, _13818_, _13881_);
  nor _22227_ (_13883_, _12084_, _12221_);
  and _22228_ (_13884_, _13883_, _13814_);
  and _22229_ (_13885_, _13884_, _13882_);
  and _22230_ (_13886_, _13882_, _12221_);
  nor _22231_ (_13887_, _12126_, _12167_);
  and _22232_ (_13888_, _13887_, _13815_);
  and _22233_ (_13889_, _13888_, _13886_);
  nor _22234_ (_13890_, _13889_, _13885_);
  nand _22235_ (_13891_, _13882_, _13837_);
  and _22236_ (_13892_, _13881_, _13839_);
  and _22237_ (_13893_, _13892_, _13831_);
  and _22238_ (_13894_, _13842_, _13881_);
  and _22239_ (_13895_, _13894_, _13839_);
  nor _22240_ (_13896_, _13895_, _13893_);
  and _22241_ (_13897_, _13828_, _13892_);
  and _22242_ (_13898_, _13882_, _13846_);
  and _22243_ (_13899_, _13888_, _13898_);
  nor _22244_ (_13900_, _13899_, _13897_);
  and _22245_ (_13901_, _13900_, _13896_);
  and _22246_ (_13902_, _13901_, _13891_);
  and _22247_ (_13903_, _13902_, _13890_);
  and _22248_ (_13904_, _13903_, _13880_);
  and _22249_ (_13905_, _13889_, _07823_);
  not _22250_ (_13906_, _12295_);
  and _22251_ (_13907_, _13885_, _13906_);
  nor _22252_ (_13908_, _13907_, _13905_);
  nand _22253_ (_13909_, _13895_, _07429_);
  and _22254_ (_13910_, _13909_, _13908_);
  nor _22255_ (_13911_, _13910_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _22256_ (_13912_, _13911_);
  and _22257_ (_13913_, _13889_, _07766_);
  not _22258_ (_13914_, _10946_);
  nor _22259_ (_13915_, _13850_, _13914_);
  and _22260_ (_13916_, _13915_, _12228_);
  nor _22261_ (_13917_, _13916_, _13913_);
  and _22262_ (_13918_, _13917_, _12435_);
  and _22263_ (_13919_, _13918_, _13912_);
  not _22264_ (_13920_, _13919_);
  nor _22265_ (_13921_, _13920_, _13904_);
  not _22266_ (_13922_, _13921_);
  and _22267_ (_13923_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _22268_ (_13924_, _13893_, _07429_);
  not _22269_ (_13925_, _13924_);
  nand _22270_ (_13926_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand _22271_ (_13927_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _22272_ (_13928_, _13927_, _13926_);
  nand _22273_ (_13929_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _22274_ (_13930_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _22275_ (_13931_, _13930_, _13929_);
  and _22276_ (_13932_, _13931_, _13928_);
  nand _22277_ (_13933_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand _22278_ (_13934_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _22279_ (_13935_, _13934_, _13933_);
  nand _22280_ (_13936_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand _22281_ (_13937_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _22282_ (_13938_, _13937_, _13936_);
  and _22283_ (_13939_, _13938_, _13935_);
  and _22284_ (_13940_, _13939_, _13932_);
  nand _22285_ (_13942_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand _22286_ (_13943_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22287_ (_13944_, _13943_, _13942_);
  nand _22288_ (_13945_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand _22289_ (_13946_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _22290_ (_13947_, _13946_, _13945_);
  and _22291_ (_13948_, _13947_, _13944_);
  nand _22292_ (_13949_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand _22293_ (_13950_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _22294_ (_13951_, _13950_, _13949_);
  nand _22295_ (_13952_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _22296_ (_13953_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22297_ (_13954_, _13953_, _13952_);
  and _22298_ (_13955_, _13954_, _13951_);
  and _22299_ (_13956_, _13955_, _13948_);
  and _22300_ (_13957_, _13956_, _13940_);
  nand _22301_ (_13958_, _13897_, _11961_);
  nand _22302_ (_13959_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22303_ (_13960_, _13959_, _13958_);
  nand _22304_ (_13961_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand _22305_ (_13962_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _22306_ (_13963_, _13962_, _13961_);
  and _22307_ (_13964_, _13963_, _13960_);
  and _22308_ (_13966_, _13898_, _13847_);
  and _22309_ (_13967_, _11399_, _11390_);
  and _22310_ (_13968_, _13967_, _08746_);
  nor _22311_ (_13969_, _13968_, _11918_);
  nor _22312_ (_13970_, _11885_, _11739_);
  nor _22313_ (_13971_, _13331_, _12541_);
  and _22314_ (_13972_, _13971_, _13970_);
  and _22315_ (_13973_, _13972_, _13969_);
  and _22316_ (_13974_, _13973_, _11866_);
  not _22317_ (_13975_, _11855_);
  and _22318_ (_13976_, _11400_, _11395_);
  nor _22319_ (_13977_, _13976_, _13975_);
  not _22320_ (_13978_, _11870_);
  nor _22321_ (_13979_, _13337_, _13978_);
  and _22322_ (_13980_, _13979_, _13977_);
  and _22323_ (_13981_, _13980_, _13974_);
  and _22324_ (_13982_, _13981_, _11851_);
  nor _22325_ (_13983_, _13982_, _11744_);
  nor _22326_ (_13985_, _13983_, p3_in[3]);
  not _22327_ (_13986_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _22328_ (_13987_, _13983_, _13986_);
  nor _22329_ (_13988_, _13987_, _13985_);
  nand _22330_ (_13990_, _13988_, _13966_);
  and _22331_ (_13991_, _13853_, _13882_);
  nor _22332_ (_13993_, _13983_, p2_in[3]);
  not _22333_ (_13994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _22334_ (_13996_, _13983_, _13994_);
  nor _22335_ (_13997_, _13996_, _13993_);
  nand _22336_ (_13998_, _13997_, _13991_);
  and _22337_ (_13999_, _13998_, _13990_);
  and _22338_ (_14000_, _13882_, _13839_);
  nor _22339_ (_14002_, _13983_, p0_in[3]);
  not _22340_ (_14003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _22341_ (_14004_, _13983_, _14003_);
  nor _22342_ (_14005_, _14004_, _14002_);
  nand _22343_ (_14006_, _14005_, _14000_);
  and _22344_ (_14007_, _13874_, _13882_);
  nor _22345_ (_00002_, _13983_, p1_in[3]);
  not _22346_ (_00003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _22347_ (_00004_, _13983_, _00003_);
  nor _22348_ (_00005_, _00004_, _00002_);
  nand _22349_ (_00006_, _00005_, _14007_);
  and _22350_ (_00007_, _00006_, _14006_);
  and _22351_ (_00008_, _00007_, _13999_);
  and _22352_ (_00009_, _00008_, _13964_);
  nand _22353_ (_00010_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _22354_ (_00011_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _22355_ (_00012_, _00011_, _00010_);
  and _22356_ (_00013_, _00012_, _00009_);
  nand _22357_ (_00015_, _00013_, _13957_);
  nand _22358_ (_00016_, _00015_, _13919_);
  nand _22359_ (_00017_, _00016_, _13925_);
  or _22360_ (_00018_, _00017_, _13923_);
  nand _22361_ (_00019_, _13924_, _11791_);
  and _22362_ (_00020_, _00019_, _06071_);
  and _22363_ (_12226_, _00020_, _00018_);
  and _22364_ (_00021_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _22365_ (_00022_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _22366_ (_00023_, _00022_, _00021_);
  and _22367_ (_12229_, _00023_, _06071_);
  and _22368_ (_00024_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _22369_ (_00025_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _22370_ (_00026_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _22371_ (_00027_, _00026_, _00025_);
  and _22372_ (_00028_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _22373_ (_00029_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _22374_ (_00030_, _00029_, _00028_);
  or _22375_ (_00031_, _00030_, _00027_);
  and _22376_ (_00032_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _22377_ (_00033_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _22378_ (_00034_, _00033_, _00032_);
  and _22379_ (_00035_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _22380_ (_00036_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _22381_ (_00037_, _00036_, _00035_);
  or _22382_ (_00038_, _00037_, _00034_);
  or _22383_ (_00039_, _00038_, _00031_);
  and _22384_ (_00040_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _22385_ (_00041_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or _22386_ (_00042_, _00041_, _00040_);
  and _22387_ (_00043_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22388_ (_00044_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _22389_ (_00045_, _00044_, _00043_);
  or _22390_ (_00046_, _00045_, _00042_);
  and _22391_ (_00047_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _22392_ (_00048_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _22393_ (_00049_, _00048_, _00047_);
  and _22394_ (_00050_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22395_ (_00051_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _22396_ (_00052_, _00051_, _00050_);
  or _22397_ (_00053_, _00052_, _00049_);
  or _22398_ (_00054_, _00053_, _00046_);
  or _22399_ (_00055_, _00054_, _00039_);
  and _22400_ (_00056_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _22401_ (_00057_, _13897_, _12398_);
  or _22402_ (_00058_, _00057_, _00056_);
  and _22403_ (_00059_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _22404_ (_00060_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _22405_ (_00061_, _00060_, _00059_);
  or _22406_ (_00062_, _00061_, _00058_);
  or _22407_ (_00063_, _13983_, p0_in[2]);
  not _22408_ (_00064_, _13983_);
  or _22409_ (_00065_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _22410_ (_00066_, _00065_, _00063_);
  and _22411_ (_00067_, _00066_, _14000_);
  or _22412_ (_00068_, _13983_, p1_in[2]);
  or _22413_ (_00069_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _22414_ (_00070_, _00069_, _00068_);
  and _22415_ (_00071_, _00070_, _14007_);
  or _22416_ (_00072_, _00071_, _00067_);
  or _22417_ (_00073_, _13983_, p3_in[2]);
  or _22418_ (_00074_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _22419_ (_00075_, _00074_, _00073_);
  and _22420_ (_00076_, _00075_, _13966_);
  or _22421_ (_00077_, _13983_, p2_in[2]);
  or _22422_ (_00078_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _22423_ (_00079_, _00078_, _00077_);
  and _22424_ (_00080_, _00079_, _13991_);
  or _22425_ (_00081_, _00080_, _00076_);
  or _22426_ (_00082_, _00081_, _00072_);
  or _22427_ (_00083_, _00082_, _00062_);
  and _22428_ (_00084_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _22429_ (_00085_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _22430_ (_00086_, _00085_, _00084_);
  or _22431_ (_00087_, _00086_, _00083_);
  or _22432_ (_00088_, _00087_, _00055_);
  and _22433_ (_00089_, _00088_, _13919_);
  or _22434_ (_00090_, _00089_, _13924_);
  or _22435_ (_00091_, _00090_, _00024_);
  or _22436_ (_00092_, _13925_, _07564_);
  and _22437_ (_00093_, _00092_, _06071_);
  and _22438_ (_12232_, _00093_, _00091_);
  and _22439_ (_00094_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _22440_ (_00095_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _22441_ (_00096_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _22442_ (_00097_, _00096_, _00095_);
  and _22443_ (_00098_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _22444_ (_00099_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _22445_ (_00100_, _00099_, _00098_);
  or _22446_ (_00101_, _00100_, _00097_);
  and _22447_ (_00102_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _22448_ (_00103_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _22449_ (_00104_, _00103_, _00102_);
  and _22450_ (_00105_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _22451_ (_00106_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _22452_ (_00107_, _00106_, _00105_);
  or _22453_ (_00108_, _00107_, _00104_);
  or _22454_ (_00109_, _00108_, _00101_);
  and _22455_ (_00110_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22456_ (_00111_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _22457_ (_00112_, _00111_, _00110_);
  and _22458_ (_00113_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22459_ (_00114_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _22460_ (_00115_, _00114_, _00113_);
  or _22461_ (_00116_, _00115_, _00112_);
  and _22462_ (_00117_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _22463_ (_00118_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _22464_ (_00119_, _00118_, _00117_);
  and _22465_ (_00120_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22466_ (_00121_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _22467_ (_00122_, _00121_, _00120_);
  or _22468_ (_00123_, _00122_, _00119_);
  or _22469_ (_00124_, _00123_, _00116_);
  or _22470_ (_00125_, _00124_, _00109_);
  and _22471_ (_00126_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _22472_ (_00127_, _13897_, _12379_);
  or _22473_ (_00128_, _00127_, _00126_);
  and _22474_ (_00129_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _22475_ (_00130_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _22476_ (_00131_, _00130_, _00129_);
  or _22477_ (_00132_, _00131_, _00128_);
  or _22478_ (_00133_, _13983_, p0_in[1]);
  or _22479_ (_00134_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _22480_ (_00135_, _00134_, _00133_);
  and _22481_ (_00136_, _00135_, _14000_);
  or _22482_ (_00137_, _13983_, p1_in[1]);
  or _22483_ (_00138_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _22484_ (_00139_, _00138_, _00137_);
  and _22485_ (_00140_, _00139_, _14007_);
  or _22486_ (_00141_, _00140_, _00136_);
  or _22487_ (_00142_, _13983_, p2_in[1]);
  or _22488_ (_00143_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _22489_ (_00144_, _00143_, _00142_);
  and _22490_ (_00145_, _00144_, _13991_);
  or _22491_ (_00146_, _13983_, p3_in[1]);
  or _22492_ (_00147_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _22493_ (_00148_, _00147_, _00146_);
  and _22494_ (_00149_, _00148_, _13966_);
  or _22495_ (_00150_, _00149_, _00145_);
  or _22496_ (_00151_, _00150_, _00141_);
  or _22497_ (_00152_, _00151_, _00132_);
  and _22498_ (_00153_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _22499_ (_00154_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _22500_ (_00155_, _00154_, _00153_);
  or _22501_ (_00156_, _00155_, _00152_);
  or _22502_ (_00157_, _00156_, _00125_);
  and _22503_ (_00158_, _00157_, _13919_);
  or _22504_ (_00159_, _00158_, _13924_);
  or _22505_ (_00160_, _00159_, _00094_);
  nand _22506_ (_00161_, _13924_, _08110_);
  and _22507_ (_00162_, _00161_, _06071_);
  and _22508_ (_12235_, _00162_, _00160_);
  or _22509_ (_00163_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _22510_ (_00164_, _06530_, _05749_);
  and _22511_ (_00165_, _00164_, _06071_);
  and _22512_ (_12254_, _00165_, _00163_);
  or _22513_ (_00166_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  nand _22514_ (_00167_, _06530_, _11276_);
  and _22515_ (_00168_, _00167_, _06071_);
  and _22516_ (_12261_, _00168_, _00166_);
  nand _22517_ (_00169_, _13924_, _08053_);
  and _22518_ (_00170_, _00169_, _06071_);
  nand _22519_ (_00171_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _22520_ (_00172_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _22521_ (_00173_, _00172_, _00171_);
  nand _22522_ (_00174_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _22523_ (_00175_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _22524_ (_00176_, _00175_, _00174_);
  and _22525_ (_00177_, _00176_, _00173_);
  nand _22526_ (_00178_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _22527_ (_00179_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _22528_ (_00180_, _00179_, _00178_);
  nand _22529_ (_00181_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _22530_ (_00182_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _22531_ (_00183_, _00182_, _00181_);
  and _22532_ (_00184_, _00183_, _00180_);
  and _22533_ (_00185_, _00184_, _00177_);
  nand _22534_ (_00187_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _22535_ (_00188_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _22536_ (_00189_, _00188_, _00187_);
  nand _22537_ (_00190_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _22538_ (_00191_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _22539_ (_00192_, _00191_, _00190_);
  and _22540_ (_00193_, _00192_, _00189_);
  nand _22541_ (_00194_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand _22542_ (_00195_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _22543_ (_00196_, _00195_, _00194_);
  nand _22544_ (_00197_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22545_ (_00198_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _22546_ (_00199_, _00198_, _00197_);
  and _22547_ (_00200_, _00199_, _00196_);
  and _22548_ (_00201_, _00200_, _00193_);
  and _22549_ (_00202_, _00201_, _00185_);
  nand _22550_ (_00203_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _22551_ (_00204_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _22552_ (_00205_, _00204_, _00203_);
  nand _22553_ (_00206_, _13897_, _12337_);
  nand _22554_ (_00207_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _22555_ (_00208_, _00207_, _00206_);
  and _22556_ (_00209_, _00208_, _00205_);
  nor _22557_ (_00210_, _13983_, p2_in[0]);
  not _22558_ (_00211_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _22559_ (_00212_, _13983_, _00211_);
  nor _22560_ (_00213_, _00212_, _00210_);
  nand _22561_ (_00214_, _00213_, _13991_);
  nor _22562_ (_00215_, _13983_, p3_in[0]);
  not _22563_ (_00216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _22564_ (_00217_, _13983_, _00216_);
  nor _22565_ (_00218_, _00217_, _00215_);
  nand _22566_ (_00219_, _00218_, _13966_);
  and _22567_ (_00220_, _00219_, _00214_);
  nor _22568_ (_00221_, _13983_, p0_in[0]);
  not _22569_ (_00222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _22570_ (_00223_, _13983_, _00222_);
  nor _22571_ (_00224_, _00223_, _00221_);
  nand _22572_ (_00225_, _00224_, _14000_);
  nor _22573_ (_00226_, _13983_, p1_in[0]);
  not _22574_ (_00227_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _22575_ (_00228_, _13983_, _00227_);
  nor _22576_ (_00229_, _00228_, _00226_);
  nand _22577_ (_00230_, _00229_, _14007_);
  and _22578_ (_00231_, _00230_, _00225_);
  and _22579_ (_00232_, _00231_, _00220_);
  and _22580_ (_00233_, _00232_, _00209_);
  nand _22581_ (_00234_, _08811_, _07872_);
  or _22582_ (_00235_, _08811_, _07872_);
  nand _22583_ (_00236_, _00235_, _00234_);
  or _22584_ (_00237_, _07772_, _07715_);
  and _22585_ (_00238_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _22586_ (_00239_, _06006_, _06161_);
  nor _22587_ (_00240_, _00239_, _10928_);
  nor _22588_ (_00241_, _00240_, _08806_);
  nor _22589_ (_00242_, _00241_, _00238_);
  and _22590_ (_00243_, _00242_, _07830_);
  nand _22591_ (_00244_, _00243_, _00237_);
  and _22592_ (_00245_, _07823_, _07746_);
  not _22593_ (_00246_, _00245_);
  and _22594_ (_00247_, _00246_, _00244_);
  or _22595_ (_00248_, _00247_, _08952_);
  nand _22596_ (_00249_, _00247_, _08952_);
  and _22597_ (_00250_, _00249_, _00248_);
  nand _22598_ (_00251_, _00250_, _00236_);
  or _22599_ (_00252_, _00250_, _00236_);
  nand _22600_ (_00253_, _00252_, _00251_);
  or _22601_ (_00254_, _08110_, _07772_);
  and _22602_ (_00255_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not _22603_ (_00256_, _06362_);
  nor _22604_ (_00257_, _06803_, _00256_);
  nor _22605_ (_00259_, _06362_, _06226_);
  nor _22606_ (_00260_, _00259_, _00257_);
  nor _22607_ (_00261_, _00260_, _08806_);
  nor _22608_ (_00262_, _00261_, _00255_);
  and _22609_ (_00263_, _00262_, _07830_);
  nand _22610_ (_00265_, _00263_, _00254_);
  and _22611_ (_00266_, _08169_, _07823_);
  not _22612_ (_00267_, _00266_);
  and _22613_ (_00268_, _00267_, _00265_);
  or _22614_ (_00269_, _00268_, _08964_);
  nand _22615_ (_00270_, _00268_, _08964_);
  nand _22616_ (_00271_, _00270_, _00269_);
  and _22617_ (_00272_, _07773_, _07564_);
  and _22618_ (_00273_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _22619_ (_00274_, _07754_);
  nor _22620_ (_00275_, _00274_, _06803_);
  nor _22621_ (_00276_, _07754_, _06237_);
  or _22622_ (_00277_, _00276_, _00275_);
  and _22623_ (_00278_, _00277_, _08805_);
  or _22624_ (_00279_, _00278_, _00273_);
  or _22625_ (_00280_, _00279_, _07823_);
  or _22626_ (_00281_, _00280_, _00272_);
  or _22627_ (_00282_, _07830_, _07594_);
  and _22628_ (_00283_, _00282_, _00281_);
  or _22629_ (_00284_, _11791_, _07772_);
  and _22630_ (_00285_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _22631_ (_00286_, _07105_, _08799_);
  nor _22632_ (_00287_, _07105_, _06183_);
  nor _22633_ (_00288_, _00287_, _00286_);
  nor _22634_ (_00289_, _00288_, _08806_);
  nor _22635_ (_00290_, _00289_, _00285_);
  and _22636_ (_00291_, _00290_, _07830_);
  and _22637_ (_00292_, _00291_, _00284_);
  and _22638_ (_00293_, _12466_, _07823_);
  or _22639_ (_00294_, _00293_, _00292_);
  nand _22640_ (_00295_, _00294_, _00283_);
  or _22641_ (_00296_, _00294_, _00283_);
  and _22642_ (_00297_, _00296_, _00295_);
  nand _22643_ (_00298_, _00297_, _00271_);
  or _22644_ (_00299_, _00297_, _00271_);
  nand _22645_ (_00300_, _00299_, _00298_);
  nand _22646_ (_00301_, _00300_, _00253_);
  or _22647_ (_00302_, _00300_, _00253_);
  nand _22648_ (_00303_, _00302_, _00301_);
  nand _22649_ (_00304_, _00303_, _13885_);
  nand _22650_ (_00305_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _22651_ (_00306_, _00305_, _00304_);
  and _22652_ (_00307_, _00306_, _00233_);
  and _22653_ (_00308_, _00307_, _00202_);
  nor _22654_ (_00309_, _00308_, _13920_);
  nand _22655_ (_00310_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _22656_ (_00311_, _00310_, _13925_);
  or _22657_ (_00312_, _00311_, _00309_);
  and _22658_ (_12265_, _00312_, _00170_);
  nor _22659_ (_12281_, _12323_, rst);
  nor _22660_ (_12287_, _12122_, rst);
  nor _22661_ (_12290_, _11511_, rst);
  nor _22662_ (_00313_, _11248_, _11095_);
  nor _22663_ (_00314_, _00313_, _11249_);
  or _22664_ (_00315_, _00314_, _09711_);
  or _22665_ (_00317_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _22666_ (_00318_, _00317_, _11270_);
  and _22667_ (_00319_, _00318_, _00315_);
  and _22668_ (_00320_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _22669_ (_12293_, _00320_, _00319_);
  nor _22670_ (_12300_, _11570_, rst);
  or _22671_ (_00322_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _22672_ (_00323_, _00322_, _13711_);
  nand _22673_ (_00324_, _00256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _22674_ (_00325_, _00324_, _13711_);
  or _22675_ (_00326_, _00325_, _00257_);
  and _22676_ (_00327_, _00326_, _00323_);
  or _22677_ (_00328_, _00327_, _13718_);
  nand _22678_ (_00329_, _13718_, _09037_);
  and _22679_ (_00330_, _00329_, _06071_);
  and _22680_ (_12303_, _00330_, _00328_);
  nand _22681_ (_00331_, _13723_, _06434_);
  or _22682_ (_00332_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _22683_ (_00333_, _00332_, _06071_);
  and _22684_ (_12315_, _00333_, _00331_);
  nor _22685_ (_00334_, _11723_, _11471_);
  nor _22686_ (_00335_, _11718_, _11472_);
  or _22687_ (_00336_, _00335_, _00334_);
  nand _22688_ (_00337_, _00336_, _06243_);
  or _22689_ (_00338_, _00336_, _06243_);
  and _22690_ (_00339_, _00338_, _00337_);
  and _22691_ (_00340_, _00339_, _11751_);
  and _22692_ (_00341_, _11827_, _07564_);
  and _22693_ (_00342_, _11748_, _07594_);
  and _22694_ (_00343_, _11628_, _11424_);
  and _22695_ (_00344_, _12469_, _05768_);
  and _22696_ (_00345_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _22697_ (_00346_, _00345_, _00344_);
  or _22698_ (_00347_, _00346_, _00343_);
  nor _22699_ (_00348_, _00347_, _00342_);
  nand _22700_ (_00349_, _00348_, _12437_);
  or _22701_ (_00350_, _00349_, _00341_);
  or _22702_ (_00351_, _00350_, _00340_);
  and _22703_ (_00352_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _22704_ (_00353_, _00352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _22705_ (_00354_, _00353_, _12503_);
  or _22706_ (_00355_, _00354_, _12437_);
  and _22707_ (_00356_, _00355_, _06071_);
  and _22708_ (_12327_, _00356_, _00351_);
  and _22709_ (_00357_, _13753_, _12197_);
  and _22710_ (_00358_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _22711_ (_00360_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _22712_ (_00361_, _00360_, _00358_);
  nor _22713_ (_00362_, _00361_, _13744_);
  nor _22714_ (_00363_, _13760_, _07945_);
  or _22715_ (_00364_, _00363_, _00362_);
  or _22716_ (_00365_, _00364_, _00357_);
  and _22717_ (_12331_, _00365_, _06071_);
  not _22718_ (_00366_, _07643_);
  or _22719_ (_00367_, _12485_, _11748_);
  and _22720_ (_00368_, _00367_, _00366_);
  nor _22721_ (_00369_, _11428_, _11053_);
  and _22722_ (_00370_, _12469_, _12131_);
  nor _22723_ (_00371_, _11533_, _11425_);
  or _22724_ (_00372_, _00371_, _00370_);
  or _22725_ (_00373_, _00372_, _00369_);
  not _22726_ (_00374_, _11709_);
  or _22727_ (_00375_, _11552_, _11553_);
  or _22728_ (_00376_, _00375_, _00374_);
  nand _22729_ (_00377_, _00375_, _00374_);
  and _22730_ (_00378_, _00377_, _11751_);
  and _22731_ (_00379_, _00378_, _00376_);
  or _22732_ (_00380_, _00379_, _00373_);
  nor _22733_ (_00381_, _00380_, _00368_);
  nand _22734_ (_00382_, _00381_, _12437_);
  and _22735_ (_00383_, _11250_, _08178_);
  and _22736_ (_00384_, _00383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _22737_ (_00385_, _00383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _22738_ (_00386_, _00385_, _00384_);
  or _22739_ (_00387_, _00386_, _12437_);
  and _22740_ (_00389_, _00387_, _06071_);
  and _22741_ (_12334_, _00389_, _00382_);
  nor _22742_ (_00390_, _11261_, _11079_);
  nor _22743_ (_00391_, _00390_, _11262_);
  or _22744_ (_00392_, _00391_, _09711_);
  or _22745_ (_00394_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _22746_ (_00395_, _00394_, _11270_);
  and _22747_ (_00396_, _00395_, _00392_);
  and _22748_ (_00397_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _22749_ (_12342_, _00397_, _00396_);
  nor _22750_ (_00398_, _11247_, _11245_);
  nor _22751_ (_00399_, _00398_, _11248_);
  or _22752_ (_00400_, _00399_, _09711_);
  or _22753_ (_00401_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _22754_ (_00402_, _00401_, _11270_);
  and _22755_ (_00403_, _00402_, _00400_);
  and _22756_ (_00404_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _22757_ (_12345_, _00404_, _00403_);
  nor _22758_ (_00405_, _11236_, _06528_);
  nand _22759_ (_00406_, _00405_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _22760_ (_00407_, _00405_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _22761_ (_00408_, _00407_, _11270_);
  and _22762_ (_12358_, _00408_, _00406_);
  and _22763_ (_00409_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _22764_ (_00410_, _00409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _22765_ (_12361_, _00410_, _06071_);
  nor _22766_ (_12367_, _11648_, rst);
  nor _22767_ (_00411_, _13796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _22768_ (_00412_, _13796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _22769_ (_00413_, _00412_, _00411_);
  and _22770_ (_12373_, _00413_, _13798_);
  and _22771_ (_00414_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _08003_);
  and _22772_ (_00415_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22773_ (_00416_, _00415_, _00414_);
  and _22774_ (_12392_, _00416_, _06071_);
  or _22775_ (_00417_, _08992_, rxd_i);
  nand _22776_ (_00418_, _00417_, _07903_);
  or _22777_ (_00419_, _07904_, _07889_);
  and _22778_ (_00420_, _00419_, _00418_);
  not _22779_ (_00421_, _07886_);
  nand _22780_ (_00422_, _07910_, _00421_);
  or _22781_ (_00423_, _00422_, _00420_);
  and _22782_ (_12396_, _00423_, _06560_);
  not _22783_ (_00424_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _22784_ (_00425_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _22785_ (_00426_, _00425_, _00424_);
  and _22786_ (_00427_, _00426_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _22787_ (_00428_, _00425_, _00424_);
  or _22788_ (_00429_, _00428_, _00426_);
  nand _22789_ (_00431_, _00429_, _06071_);
  nor _22790_ (_12415_, _00431_, _00427_);
  or _22791_ (_00432_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _22792_ (_00434_, _00425_, rst);
  and _22793_ (_12440_, _00434_, _00432_);
  nor _22794_ (_12448_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  not _22795_ (_00435_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _22796_ (_00436_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _22797_ (_00437_, _07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _22798_ (_00438_, _00437_, _00436_);
  nor _22799_ (_00439_, _00438_, _00435_);
  and _22800_ (_00440_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _22801_ (_00441_, _00440_, _00439_);
  or _22802_ (_00442_, _00441_, _13711_);
  or _22803_ (_00443_, _07754_, _00435_);
  nand _22804_ (_00444_, _00443_, _13711_);
  or _22805_ (_00445_, _00444_, _00275_);
  and _22806_ (_00446_, _00445_, _00442_);
  or _22807_ (_00447_, _00446_, _13718_);
  nand _22808_ (_00448_, _13718_, _06434_);
  and _22809_ (_00449_, _00448_, _06071_);
  and _22810_ (_12461_, _00449_, _00447_);
  nand _22811_ (_00450_, _13723_, _07945_);
  or _22812_ (_00451_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22813_ (_00452_, _00451_, _06071_);
  and _22814_ (_12468_, _00452_, _00450_);
  and _22815_ (_00453_, _13753_, _12161_);
  and _22816_ (_00454_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _22817_ (_00455_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _22818_ (_00456_, _00455_, _00454_);
  nor _22819_ (_00457_, _00456_, _13744_);
  nor _22820_ (_00458_, _13760_, _06993_);
  or _22821_ (_00459_, _00458_, _00457_);
  or _22822_ (_00460_, _00459_, _00453_);
  and _22823_ (_12471_, _00460_, _06071_);
  or _22824_ (_00461_, _11719_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _22825_ (_00462_, _00461_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _22826_ (_00463_, _00462_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _22827_ (_00464_, _00463_, _11471_);
  and _22828_ (_00465_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _22829_ (_00466_, _00465_, _11722_);
  and _22830_ (_00467_, _00466_, _11716_);
  and _22831_ (_00468_, _00467_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _22832_ (_00469_, _00468_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _22833_ (_00471_, _00469_, _11472_);
  and _22834_ (_00472_, _00471_, _00464_);
  nor _22835_ (_00473_, _00472_, _06261_);
  and _22836_ (_00474_, _00472_, _06261_);
  or _22837_ (_00476_, _00474_, _00473_);
  and _22838_ (_00477_, _00476_, _11751_);
  and _22839_ (_00478_, _11827_, _07425_);
  and _22840_ (_00479_, _11748_, _07520_);
  and _22841_ (_00480_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _22842_ (_00481_, _00480_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _22843_ (_00482_, _00481_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _22844_ (_00483_, _00481_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _22845_ (_00484_, _00483_, _00482_);
  and _22846_ (_00485_, _00484_, _12469_);
  and _22847_ (_00486_, _12090_, _11424_);
  and _22848_ (_00487_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _22849_ (_00488_, _00487_, _00486_);
  or _22850_ (_00489_, _00488_, _00485_);
  or _22851_ (_00490_, _00489_, _00479_);
  nor _22852_ (_00491_, _00490_, _00478_);
  nand _22853_ (_00492_, _00491_, _12437_);
  or _22854_ (_00493_, _00492_, _00477_);
  and _22855_ (_00494_, _00352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _22856_ (_00495_, _00494_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _22857_ (_00496_, _00495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _22858_ (_00497_, _00496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22859_ (_00498_, _00497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _22860_ (_00499_, _00497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _22861_ (_00500_, _00499_, _00498_);
  or _22862_ (_00501_, _00500_, _12437_);
  and _22863_ (_00502_, _00501_, _06071_);
  and _22864_ (_12490_, _00502_, _00493_);
  and _22865_ (_00504_, _00462_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _22866_ (_00505_, _00504_, _00464_);
  or _22867_ (_00506_, _00468_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _22868_ (_00507_, _00506_, _00469_);
  or _22869_ (_00508_, _00507_, _11471_);
  and _22870_ (_00509_, _00508_, _11751_);
  and _22871_ (_00510_, _00509_, _00505_);
  nor _22872_ (_00511_, _11428_, _07643_);
  nor _22873_ (_00512_, _12438_, _07673_);
  nor _22874_ (_00513_, _00480_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _22875_ (_00514_, _00513_, _00481_);
  and _22876_ (_00515_, _00514_, _12469_);
  and _22877_ (_00516_, _12131_, _11424_);
  or _22878_ (_00517_, _00516_, _00515_);
  and _22879_ (_00518_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22880_ (_00519_, _00518_, _00517_);
  nor _22881_ (_00520_, _00519_, _00512_);
  nand _22882_ (_00521_, _00520_, _12437_);
  or _22883_ (_00522_, _00521_, _00511_);
  or _22884_ (_00523_, _00522_, _00510_);
  nor _22885_ (_00524_, _00496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _22886_ (_00525_, _00524_, _00497_);
  or _22887_ (_00526_, _00525_, _12437_);
  and _22888_ (_00527_, _00526_, _06071_);
  and _22889_ (_12496_, _00527_, _00523_);
  and _22890_ (_00528_, _00467_, _11472_);
  nor _22891_ (_00529_, _11721_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _22892_ (_00530_, _00529_, _00528_);
  nand _22893_ (_00532_, _00530_, _06151_);
  or _22894_ (_00533_, _00530_, _06151_);
  and _22895_ (_00534_, _00533_, _00532_);
  and _22896_ (_00535_, _00534_, _11751_);
  nor _22897_ (_00536_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _22898_ (_00537_, _00536_, _00480_);
  and _22899_ (_00538_, _00537_, _12469_);
  nor _22900_ (_00539_, _11428_, _07715_);
  nor _22901_ (_00540_, _12438_, _07746_);
  and _22902_ (_00541_, _11424_, _12172_);
  and _22903_ (_00542_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _22904_ (_00543_, _00542_, _00541_);
  or _22905_ (_00544_, _00543_, _00540_);
  or _22906_ (_00545_, _00544_, _00539_);
  nor _22907_ (_00546_, _00545_, _00538_);
  nand _22908_ (_00547_, _00546_, _12437_);
  or _22909_ (_00548_, _00547_, _00535_);
  nor _22910_ (_00549_, _12505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _22911_ (_00550_, _00549_, _00496_);
  or _22912_ (_00551_, _00550_, _12437_);
  and _22913_ (_00552_, _00551_, _06071_);
  and _22914_ (_12526_, _00552_, _00548_);
  nor _22915_ (_00553_, _07881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _22916_ (_00554_, _00553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _22917_ (_00555_, _00553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _22918_ (_00556_, _00555_, _06071_);
  and _22919_ (_12554_, _00556_, _00554_);
  not _22920_ (_00557_, _13718_);
  and _22921_ (_00558_, _13711_, _07105_);
  and _22922_ (_00559_, _00558_, _06803_);
  nor _22923_ (_00560_, _00558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _22924_ (_00561_, _00560_, _00559_);
  nand _22925_ (_00562_, _00561_, _00557_);
  nand _22926_ (_00564_, _13718_, _07945_);
  and _22927_ (_00565_, _00564_, _06071_);
  and _22928_ (_12557_, _00565_, _00562_);
  and _22929_ (_00566_, _13753_, _12120_);
  and _22930_ (_00567_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _22931_ (_00568_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _22932_ (_00569_, _00568_, _00567_);
  nor _22933_ (_00570_, _00569_, _13744_);
  nor _22934_ (_00571_, _13760_, _06609_);
  or _22935_ (_00573_, _00571_, _00570_);
  or _22936_ (_00575_, _00573_, _00566_);
  and _22937_ (_12560_, _00575_, _06071_);
  not _22938_ (_00576_, _13711_);
  or _22939_ (_00577_, _00576_, _10936_);
  and _22940_ (_00578_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22941_ (_00579_, _00578_, _13718_);
  nor _22942_ (_00580_, _10930_, _08993_);
  or _22943_ (_00581_, _00580_, _10928_);
  and _22944_ (_00582_, _00581_, _13711_);
  or _22945_ (_00583_, _00582_, _00579_);
  nand _22946_ (_00584_, _13718_, _06993_);
  and _22947_ (_00585_, _00584_, _06071_);
  and _22948_ (_12600_, _00585_, _00583_);
  nor _22949_ (_00586_, _09341_, _06611_);
  and _22950_ (_00587_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _22951_ (_00588_, _00587_, _00586_);
  and _22952_ (_12624_, _00588_, _06071_);
  nand _22953_ (_00589_, _11791_, _10978_);
  or _22954_ (_00590_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _22955_ (_00591_, _00590_, _06071_);
  and _22956_ (_12694_, _00591_, _00589_);
  nor _22957_ (_12907_, _11931_, rst);
  not _22958_ (_00593_, _07715_);
  and _22959_ (_00594_, _00367_, _00593_);
  or _22960_ (_00595_, _11707_, _11705_);
  and _22961_ (_00596_, _11751_, _11708_);
  and _22962_ (_00597_, _00596_, _00595_);
  and _22963_ (_00598_, _12469_, _12172_);
  nor _22964_ (_00599_, _11570_, _11425_);
  and _22965_ (_00600_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _22966_ (_00601_, _00600_, _00599_);
  or _22967_ (_00602_, _00601_, _00598_);
  or _22968_ (_00603_, _00602_, _00597_);
  nor _22969_ (_00604_, _00603_, _00594_);
  nand _22970_ (_00605_, _00604_, _12437_);
  nor _22971_ (_00606_, _08180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _22972_ (_00607_, _00606_, _00383_);
  or _22973_ (_00608_, _00607_, _12437_);
  and _22974_ (_00609_, _00608_, _06071_);
  and _22975_ (_13034_, _00609_, _00605_);
  or _22976_ (_00610_, _12437_, _08181_);
  and _22977_ (_00611_, _00610_, _06071_);
  not _22978_ (_00612_, _11791_);
  and _22979_ (_00613_, _00367_, _00612_);
  or _22980_ (_00614_, _11610_, _11611_);
  not _22981_ (_00615_, _00614_);
  nand _22982_ (_00616_, _00615_, _11703_);
  or _22983_ (_00617_, _00615_, _11703_);
  and _22984_ (_00619_, _00617_, _11751_);
  and _22985_ (_00620_, _00619_, _00616_);
  nor _22986_ (_00622_, _11591_, _11425_);
  and _22987_ (_00623_, _12469_, _12024_);
  or _22988_ (_00624_, _00623_, _00622_);
  or _22989_ (_00625_, _00624_, _00620_);
  or _22990_ (_00626_, _00625_, _00613_);
  nand _22991_ (_00627_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand _22992_ (_00628_, _00627_, _12437_);
  or _22993_ (_00629_, _00628_, _00626_);
  and _22994_ (_13056_, _00629_, _00611_);
  or _22995_ (_00630_, _12437_, _08192_);
  and _22996_ (_00631_, _00630_, _06071_);
  and _22997_ (_00632_, _00367_, _07564_);
  or _22998_ (_00633_, _11700_, _11698_);
  and _22999_ (_00634_, _11751_, _11702_);
  and _23000_ (_00635_, _00634_, _00633_);
  nor _23001_ (_00636_, _11428_, _08177_);
  and _23002_ (_00637_, _11424_, _11612_);
  and _23003_ (_00638_, _12469_, _11628_);
  or _23004_ (_00639_, _00638_, _00637_);
  or _23005_ (_00640_, _00639_, _00636_);
  or _23006_ (_00642_, _00640_, _00635_);
  nor _23007_ (_00643_, _00642_, _00632_);
  nand _23008_ (_00644_, _00643_, _12437_);
  and _23009_ (_13085_, _00644_, _00631_);
  not _23010_ (_00645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _23011_ (_00646_, _12437_, _11428_);
  nor _23012_ (_00647_, _00646_, _00645_);
  and _23013_ (_00648_, _11649_, _11424_);
  and _23014_ (_00649_, _12469_, _11651_);
  or _23015_ (_00650_, _00649_, _00648_);
  or _23016_ (_00651_, _11695_, _11693_);
  and _23017_ (_00652_, _11751_, _11697_);
  and _23018_ (_00653_, _00652_, _00651_);
  or _23019_ (_00654_, _00653_, _00650_);
  not _23020_ (_00655_, _08110_);
  and _23021_ (_00656_, _00367_, _00655_);
  or _23022_ (_00657_, _00656_, _00654_);
  and _23023_ (_00658_, _00657_, _12437_);
  or _23024_ (_00659_, _00658_, _00647_);
  and _23025_ (_13098_, _00659_, _06071_);
  not _23026_ (_00660_, _08053_);
  and _23027_ (_00661_, _00367_, _00660_);
  or _23028_ (_00662_, _11691_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _23029_ (_00663_, _11693_);
  and _23030_ (_00664_, _11751_, _00663_);
  and _23031_ (_00665_, _00664_, _00662_);
  and _23032_ (_00666_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _23033_ (_00667_, _11672_, _11424_);
  and _23034_ (_00668_, _12469_, _11689_);
  or _23035_ (_00669_, _00668_, _00667_);
  or _23036_ (_00670_, _00669_, _00666_);
  or _23037_ (_00671_, _00670_, _00665_);
  nor _23038_ (_00672_, _00671_, _00661_);
  nand _23039_ (_00673_, _00672_, _12437_);
  or _23040_ (_00674_, _12437_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _23041_ (_00675_, _00674_, _06071_);
  and _23042_ (_13110_, _00675_, _00673_);
  or _23043_ (_00676_, _07819_, _07757_);
  or _23044_ (_00677_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _23045_ (_00678_, _00677_, _06071_);
  and _23046_ (_13206_, _00678_, _00676_);
  and _23047_ (_00679_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _23048_ (_00680_, _07819_, _07530_);
  or _23049_ (_00681_, _00680_, _00679_);
  or _23050_ (_00682_, _00681_, _07429_);
  or _23051_ (_00683_, _07870_, _07433_);
  and _23052_ (_00684_, _00683_, _06071_);
  and _23053_ (_13246_, _00684_, _00682_);
  and _23054_ (_00685_, _00367_, _07425_);
  or _23055_ (_00686_, _11711_, _11516_);
  and _23056_ (_00687_, _11751_, _11713_);
  and _23057_ (_00688_, _00687_, _00686_);
  nor _23058_ (_00689_, _11428_, _11052_);
  and _23059_ (_00690_, _12469_, _12090_);
  nor _23060_ (_00691_, _11493_, _11425_);
  or _23061_ (_00692_, _00691_, _00690_);
  or _23062_ (_00693_, _00692_, _00689_);
  or _23063_ (_00694_, _00693_, _00688_);
  nor _23064_ (_00695_, _00694_, _00685_);
  nand _23065_ (_00696_, _00695_, _12437_);
  and _23066_ (_00697_, _00384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _23067_ (_00698_, _00384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _23068_ (_00699_, _00698_, _00697_);
  or _23069_ (_00700_, _00699_, _12437_);
  and _23070_ (_00701_, _00700_, _06071_);
  and _23071_ (_13281_, _00701_, _00696_);
  and _23072_ (_00702_, _11716_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _23073_ (_00703_, _00702_, _11471_);
  and _23074_ (_00704_, _11717_, _11471_);
  nor _23075_ (_00705_, _00704_, _00703_);
  and _23076_ (_00706_, _00705_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _23077_ (_00707_, _00705_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _23078_ (_00708_, _00707_, _11751_);
  nor _23079_ (_00709_, _00708_, _00706_);
  nor _23080_ (_00710_, _11428_, _08110_);
  nor _23081_ (_00711_, _12438_, _08169_);
  and _23082_ (_00712_, _11424_, _11651_);
  and _23083_ (_00713_, _12469_, _05747_);
  or _23084_ (_00714_, _00713_, _00712_);
  and _23085_ (_00715_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _23086_ (_00716_, _00715_, _00714_);
  or _23087_ (_00717_, _00716_, _00711_);
  nor _23088_ (_00718_, _00717_, _00710_);
  nand _23089_ (_00719_, _00718_, _12437_);
  or _23090_ (_00720_, _00719_, _00709_);
  nor _23091_ (_00721_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _23092_ (_00722_, _00721_, _00352_);
  or _23093_ (_00723_, _00722_, _12437_);
  and _23094_ (_00724_, _00723_, _06071_);
  and _23095_ (_13289_, _00724_, _00720_);
  and _23096_ (_00726_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor _23097_ (_00727_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23098_ (_00729_, _00727_, _06510_);
  or _23099_ (_00730_, _06486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _23100_ (_00731_, _06499_, _06445_);
  and _23101_ (_00732_, _00731_, _00730_);
  or _23102_ (_00733_, _00732_, _06474_);
  and _23103_ (_00734_, _00733_, _00729_);
  or _23104_ (_00735_, _00734_, _00726_);
  and _23105_ (_00736_, _06505_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23106_ (_00737_, _00736_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _23107_ (_00738_, _00737_, _06071_);
  and _23108_ (_13324_, _00738_, _00735_);
  nor _23109_ (_00739_, _11428_, _08053_);
  nand _23110_ (_00740_, _11716_, _06193_);
  or _23111_ (_00741_, _11716_, _06193_);
  and _23112_ (_00742_, _00741_, _00740_);
  and _23113_ (_00743_, _00742_, _11471_);
  and _23114_ (_00744_, _00703_, _11717_);
  or _23115_ (_00745_, _00744_, _00743_);
  and _23116_ (_00746_, _00745_, _11751_);
  and _23117_ (_00747_, _11748_, _08139_);
  and _23118_ (_00748_, _12469_, _05726_);
  and _23119_ (_00749_, _11689_, _11424_);
  and _23120_ (_00750_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _23121_ (_00751_, _00750_, _00749_);
  nor _23122_ (_00752_, _00751_, _00748_);
  nand _23123_ (_00753_, _00752_, _12437_);
  or _23124_ (_00754_, _00753_, _00747_);
  or _23125_ (_00755_, _00754_, _00746_);
  or _23126_ (_00756_, _00755_, _00739_);
  nor _23127_ (_00757_, _12500_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _23128_ (_00758_, _00757_, _12501_);
  or _23129_ (_00759_, _00758_, _12437_);
  and _23130_ (_00760_, _00759_, _06071_);
  and _23131_ (_13328_, _00760_, _00756_);
  and _23132_ (_00761_, _07105_, _06027_);
  and _23133_ (_00762_, _00761_, _06840_);
  nand _23134_ (_00763_, _00762_, _09341_);
  not _23135_ (_00764_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _23136_ (_00765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00764_);
  not _23137_ (_00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23138_ (_00767_, _00766_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _23139_ (_00768_, t1_i);
  and _23140_ (_00769_, _00768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23141_ (_00770_, _00769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _23142_ (_00771_, _00770_, _00767_);
  and _23143_ (_00772_, _00771_, _00765_);
  and _23144_ (_00773_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23145_ (_00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23146_ (_00775_, _00774_, _00773_);
  and _23147_ (_00776_, _00775_, _00772_);
  and _23148_ (_00777_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23149_ (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _23150_ (_00779_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23151_ (_00780_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23152_ (_00782_, _00780_, _00779_);
  not _23153_ (_00783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _23154_ (_00784_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _23155_ (_00785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23156_ (_00786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00785_);
  nor _23157_ (_00787_, _00786_, _00784_);
  and _23158_ (_00788_, _09244_, _06012_);
  and _23159_ (_00789_, _06840_, _00788_);
  nor _23160_ (_00790_, _00789_, _00787_);
  and _23161_ (_00791_, _00790_, _00782_);
  not _23162_ (_00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23163_ (_00793_, _00790_, _00792_);
  and _23164_ (_00794_, _06840_, _06032_);
  and _23165_ (_00795_, _00794_, _06027_);
  and _23166_ (_00796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23167_ (_00797_, _00796_, _00778_);
  and _23168_ (_00798_, _00797_, _00784_);
  nand _23169_ (_00799_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23170_ (_00800_, _00799_, _00795_);
  or _23171_ (_00801_, _00800_, _00793_);
  or _23172_ (_00802_, _00801_, _00791_);
  or _23173_ (_00803_, _00762_, _00802_);
  and _23174_ (_00804_, _00803_, _06071_);
  and _23175_ (_13336_, _00804_, _00763_);
  and _23176_ (_00805_, _00367_, _07819_);
  nor _23177_ (_00806_, _11453_, _11425_);
  and _23178_ (_00807_, _12469_, _12080_);
  or _23179_ (_00808_, _00807_, _00806_);
  or _23180_ (_00809_, _11473_, _11474_);
  not _23181_ (_00810_, _00809_);
  nand _23182_ (_00811_, _00810_, _11714_);
  or _23183_ (_00812_, _00810_, _11714_);
  and _23184_ (_00813_, _00812_, _11751_);
  and _23185_ (_00814_, _00813_, _00811_);
  or _23186_ (_00815_, _00814_, _00808_);
  or _23187_ (_00816_, _00815_, _00805_);
  or _23188_ (_00817_, _11428_, _11051_);
  nand _23189_ (_00818_, _00817_, _12437_);
  or _23190_ (_00819_, _00818_, _00816_);
  nor _23191_ (_00820_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _23192_ (_00821_, _00820_, _12500_);
  or _23193_ (_00822_, _00821_, _12437_);
  and _23194_ (_00823_, _00822_, _06071_);
  and _23195_ (_13359_, _00823_, _00819_);
  nand _23196_ (_00824_, _00762_, _06993_);
  and _23197_ (_00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _23198_ (_00827_, _00825_, _00789_);
  not _23199_ (_00828_, _00827_);
  and _23200_ (_00829_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23201_ (_00830_, _00780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _23202_ (_00831_, _00830_, _00784_);
  and _23203_ (_00832_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _23204_ (_00833_, _00825_);
  nor _23205_ (_00834_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _23206_ (_00835_, _00834_, _00777_);
  and _23207_ (_00836_, _00835_, _00833_);
  nor _23208_ (_00837_, _00836_, _00832_);
  nor _23209_ (_00838_, _00837_, _00789_);
  or _23210_ (_00839_, _00838_, _00829_);
  or _23211_ (_00840_, _00839_, _00762_);
  and _23212_ (_00841_, _00840_, _06071_);
  and _23213_ (_13363_, _00841_, _00824_);
  and _23214_ (_00842_, _00774_, _00772_);
  and _23215_ (_00843_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _23216_ (_00844_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _23217_ (_00845_, _00844_, _00776_);
  and _23218_ (_00846_, _00845_, _00827_);
  and _23219_ (_00847_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _23220_ (_00848_, _00847_, _00846_);
  nand _23221_ (_00849_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23222_ (_00850_, _00849_, _00789_);
  or _23223_ (_00851_, _00850_, _00762_);
  or _23224_ (_00852_, _00851_, _00848_);
  nand _23225_ (_00853_, _00762_, _07945_);
  and _23226_ (_00854_, _00853_, _06071_);
  and _23227_ (_13366_, _00854_, _00852_);
  nor _23228_ (_00855_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _23229_ (_00856_, _00855_, _00843_);
  nand _23230_ (_00857_, _00856_, _00827_);
  or _23231_ (_00858_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23232_ (_00859_, _00858_, _00857_);
  and _23233_ (_00860_, _07106_, _06027_);
  nand _23234_ (_00861_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23235_ (_00862_, _00861_, _00795_);
  or _23236_ (_00863_, _00862_, _00860_);
  or _23237_ (_00865_, _00863_, _00859_);
  nand _23238_ (_00866_, _00860_, _06434_);
  and _23239_ (_00867_, _00866_, _06071_);
  and _23240_ (_13369_, _00867_, _00865_);
  and _23241_ (_00868_, _06435_, _06369_);
  or _23242_ (_00869_, _06438_, _06394_);
  and _23243_ (_00870_, _00869_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or _23244_ (_00871_, _00870_, _00868_);
  and _23245_ (_13371_, _00871_, _06071_);
  nand _23246_ (_00873_, _00762_, _06609_);
  nor _23247_ (_00874_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _23248_ (_00875_, _00874_, _00778_);
  and _23249_ (_00876_, _00875_, _00790_);
  not _23250_ (_00877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _23251_ (_00878_, _00790_, _00877_);
  nand _23252_ (_00879_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _23253_ (_00880_, _00879_, _00795_);
  or _23254_ (_00881_, _00880_, _00878_);
  or _23255_ (_00882_, _00881_, _00876_);
  or _23256_ (_00883_, _00882_, _00762_);
  and _23257_ (_00884_, _00883_, _06071_);
  and _23258_ (_13374_, _00884_, _00873_);
  and _23259_ (_00885_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23260_ (_00887_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23261_ (_00888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23262_ (_00889_, _00888_, _00796_);
  and _23263_ (_00890_, _00889_, _00887_);
  and _23264_ (_00891_, _00890_, _00784_);
  and _23265_ (_00892_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _23266_ (_00893_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _23267_ (_00894_, _00893_, _00892_);
  and _23268_ (_00895_, _00894_, _00833_);
  nor _23269_ (_00896_, _00895_, _00891_);
  nor _23270_ (_00898_, _00896_, _00789_);
  or _23271_ (_00899_, _00898_, _00860_);
  or _23272_ (_00900_, _00899_, _00885_);
  nand _23273_ (_00901_, _00762_, _07977_);
  and _23274_ (_00902_, _00901_, _06071_);
  and _23275_ (_13388_, _00902_, _00900_);
  nor _23276_ (_00903_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _23277_ (_00904_, _00903_, _00842_);
  nand _23278_ (_00905_, _00904_, _00827_);
  or _23279_ (_00906_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23280_ (_00907_, _00906_, _00905_);
  nand _23281_ (_00908_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _23282_ (_00909_, _00908_, _00795_);
  or _23283_ (_00910_, _00909_, _00860_);
  or _23284_ (_00911_, _00910_, _00907_);
  nand _23285_ (_00912_, _00762_, _09037_);
  and _23286_ (_00913_, _00912_, _06071_);
  and _23287_ (_13392_, _00913_, _00911_);
  not _23288_ (_00914_, _00762_);
  not _23289_ (_00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _23290_ (_00916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23291_ (_00917_, _00916_, _00777_);
  and _23292_ (_00918_, _00797_, _00786_);
  nor _23293_ (_00919_, _00918_, _00917_);
  and _23294_ (_00920_, _00919_, _00915_);
  nor _23295_ (_00921_, _00919_, _00915_);
  nor _23296_ (_00922_, _00921_, _00920_);
  nor _23297_ (_00923_, _00922_, _00789_);
  and _23298_ (_00924_, _00789_, _07977_);
  or _23299_ (_00925_, _00924_, _00923_);
  nand _23300_ (_00926_, _00925_, _00914_);
  nand _23301_ (_00927_, _00762_, _00915_);
  and _23302_ (_00928_, _00927_, _06071_);
  and _23303_ (_13413_, _00928_, _00926_);
  nand _23304_ (_00929_, _00789_, _09037_);
  or _23305_ (_00930_, _00921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _23306_ (_00931_, _00921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23307_ (_00932_, _00931_, _00930_);
  or _23308_ (_00933_, _00932_, _00789_);
  and _23309_ (_00934_, _00933_, _00914_);
  and _23310_ (_00935_, _00934_, _00929_);
  and _23311_ (_00936_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _23312_ (_00937_, _00936_, _00935_);
  and _23313_ (_13416_, _00937_, _06071_);
  nand _23314_ (_00938_, _00789_, _07945_);
  and _23315_ (_00939_, _00887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23316_ (_00940_, _00939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23317_ (_00941_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23318_ (_00942_, _00941_, _00940_);
  and _23319_ (_00943_, _00942_, _00916_);
  and _23320_ (_00944_, _00889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23321_ (_00945_, _00944_, _00939_);
  and _23322_ (_00946_, _00945_, _00772_);
  and _23323_ (_00947_, _00946_, _00786_);
  nor _23324_ (_00948_, _00947_, _00943_);
  and _23325_ (_00949_, _00948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23326_ (_00950_, _00948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23327_ (_00951_, _00950_, _00949_);
  or _23328_ (_00952_, _00951_, _00789_);
  and _23329_ (_00953_, _00952_, _00914_);
  and _23330_ (_00954_, _00953_, _00938_);
  and _23331_ (_00955_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23332_ (_00956_, _00955_, _00954_);
  and _23333_ (_13424_, _00956_, _06071_);
  nand _23334_ (_00957_, _00789_, _06609_);
  and _23335_ (_00958_, _00946_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23336_ (_00959_, _00958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23337_ (_00960_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _23338_ (_00961_, _00786_);
  and _23339_ (_00962_, _00890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23340_ (_00963_, _00962_, _00941_);
  and _23341_ (_00964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23342_ (_00965_, _00964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23343_ (_00966_, _00965_, _00963_);
  nor _23344_ (_00967_, _00966_, _00961_);
  and _23345_ (_00968_, _00967_, _00960_);
  and _23346_ (_00969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23347_ (_00970_, _00942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23348_ (_00971_, _00970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23349_ (_00972_, _00971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _23350_ (_00973_, _00916_);
  and _23351_ (_00974_, _00965_, _00942_);
  nor _23352_ (_00975_, _00974_, _00973_);
  and _23353_ (_00976_, _00975_, _00972_);
  or _23354_ (_00977_, _00976_, _00969_);
  or _23355_ (_00978_, _00977_, _00968_);
  or _23356_ (_00979_, _00978_, _00789_);
  and _23357_ (_00980_, _00979_, _00914_);
  and _23358_ (_00981_, _00980_, _00957_);
  and _23359_ (_00982_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _23360_ (_00983_, _00982_, _00981_);
  and _23361_ (_13427_, _00983_, _06071_);
  nand _23362_ (_00984_, _00789_, _06993_);
  or _23363_ (_00985_, _00958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _23364_ (_00986_, _00959_, _00961_);
  and _23365_ (_00987_, _00986_, _00985_);
  and _23366_ (_00988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _23367_ (_00989_, _00970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _23368_ (_00990_, _00971_, _00973_);
  and _23369_ (_00991_, _00990_, _00989_);
  or _23370_ (_00992_, _00991_, _00988_);
  or _23371_ (_00993_, _00992_, _00987_);
  or _23372_ (_00994_, _00993_, _00789_);
  and _23373_ (_00995_, _00994_, _00914_);
  and _23374_ (_00996_, _00995_, _00984_);
  and _23375_ (_00997_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23376_ (_00998_, _00997_, _00996_);
  and _23377_ (_13430_, _00998_, _06071_);
  not _23378_ (_01000_, _00795_);
  and _23379_ (_01001_, _00931_, _01000_);
  or _23380_ (_01003_, _01001_, _00860_);
  and _23381_ (_01004_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23382_ (_01005_, _01000_, _06434_);
  or _23383_ (_01007_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23384_ (_01008_, _01007_, _00795_);
  nor _23385_ (_01010_, _01008_, _01005_);
  nor _23386_ (_01011_, _01010_, _00860_);
  or _23387_ (_01012_, _01011_, _01004_);
  and _23388_ (_13433_, _01012_, _06071_);
  and _23389_ (_01014_, _09576_, _06381_);
  and _23390_ (_01016_, _13574_, _06011_);
  nand _23391_ (_01017_, _06392_, _06011_);
  or _23392_ (_01018_, _01017_, _01016_);
  and _23393_ (_01020_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _23394_ (_01021_, _01020_, _01014_);
  and _23395_ (_13436_, _01021_, _06071_);
  not _23396_ (_01022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _23397_ (_01023_, t0_i);
  and _23398_ (_01025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01023_);
  nor _23399_ (_01027_, _01025_, _01022_);
  not _23400_ (_01029_, _01027_);
  not _23401_ (_01030_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _23402_ (_01031_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _23403_ (_01032_, _01031_, _01030_);
  and _23404_ (_01033_, _01032_, _01029_);
  not _23405_ (_01034_, _01033_);
  and _23406_ (_01035_, _06840_, _06028_);
  nor _23407_ (_01037_, _01035_, _01034_);
  or _23408_ (_01038_, _01037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _23409_ (_01040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23410_ (_01041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _23411_ (_01043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _23412_ (_01044_, _01043_, _01041_);
  and _23413_ (_01046_, _01044_, _01040_);
  and _23414_ (_01047_, _01046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23415_ (_01050_, _01047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _23416_ (_01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23417_ (_01053_, _01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23418_ (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23419_ (_01055_, _01054_, _01050_);
  and _23420_ (_01057_, _01033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _23421_ (_01058_, _01057_, _01055_);
  or _23422_ (_01060_, _01058_, _01035_);
  and _23423_ (_01061_, _01060_, _01038_);
  and _23424_ (_01062_, _07754_, _06027_);
  and _23425_ (_01063_, _01062_, _06840_);
  or _23426_ (_01064_, _01063_, _01061_);
  nand _23427_ (_01065_, _01063_, _07977_);
  and _23428_ (_01066_, _01065_, _06071_);
  and _23429_ (_13439_, _01066_, _01064_);
  nor _23430_ (_01068_, _10945_, _06026_);
  and _23431_ (_01069_, _01068_, _05923_);
  and _23432_ (_01070_, _01069_, _06807_);
  and _23433_ (_01072_, _01070_, _06806_);
  and _23434_ (_01074_, _01072_, _06383_);
  or _23435_ (_01076_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23436_ (_01077_, _01076_, _09250_);
  nand _23437_ (_01079_, _01074_, _06803_);
  and _23438_ (_01080_, _01079_, _01077_);
  and _23439_ (_01081_, _09249_, _07978_);
  or _23440_ (_01082_, _01081_, _01080_);
  and _23441_ (_13441_, _01082_, _06071_);
  nor _23442_ (_01084_, _01057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _23443_ (_01085_, _01057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _23444_ (_01087_, _01085_, _01084_);
  and _23445_ (_01088_, _01050_, _01033_);
  and _23446_ (_01089_, _01088_, _01053_);
  and _23447_ (_01090_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _23448_ (_01091_, _01090_, _01087_);
  nor _23449_ (_01092_, _01091_, _01035_);
  and _23450_ (_01093_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _23451_ (_01094_, _01093_, _01092_);
  or _23452_ (_01095_, _01094_, _01063_);
  nand _23453_ (_01096_, _01063_, _09037_);
  and _23454_ (_01097_, _01096_, _06071_);
  and _23455_ (_13457_, _01097_, _01095_);
  not _23456_ (_01098_, _01063_);
  and _23457_ (_01099_, _01044_, _01033_);
  and _23458_ (_01100_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _23459_ (_01101_, _01100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _23460_ (_01102_, _01101_, _01099_);
  and _23461_ (_01103_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _23462_ (_01104_, _01103_, _01102_);
  nor _23463_ (_01105_, _01104_, _01035_);
  and _23464_ (_01106_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _23465_ (_01107_, _01106_, _01105_);
  and _23466_ (_01108_, _01107_, _01098_);
  nor _23467_ (_01109_, _01098_, _07945_);
  or _23468_ (_01110_, _01109_, _01108_);
  and _23469_ (_13461_, _01110_, _06071_);
  nor _23470_ (_01111_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _23471_ (_01112_, _01111_, _01100_);
  and _23472_ (_01113_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _23473_ (_01114_, _01113_, _01112_);
  nor _23474_ (_01115_, _01114_, _01035_);
  and _23475_ (_01116_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _23476_ (_01117_, _01116_, _01115_);
  and _23477_ (_01118_, _01117_, _01098_);
  nor _23478_ (_01119_, _01098_, _06434_);
  or _23479_ (_01120_, _01119_, _01118_);
  and _23480_ (_13464_, _01120_, _06071_);
  or _23481_ (_01121_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23482_ (_01122_, _01121_, _06071_);
  or _23483_ (_01123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _23484_ (_01124_, _01123_, _06453_);
  or _23485_ (_01125_, _01124_, _06459_);
  and _23486_ (_01126_, _06463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23487_ (_01127_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23488_ (_01128_, _06467_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23489_ (_01129_, _01128_, _06470_);
  and _23490_ (_01130_, _01129_, _01127_);
  nand _23491_ (_01131_, _09237_, _06470_);
  nand _23492_ (_01132_, _01131_, _06458_);
  or _23493_ (_01133_, _01132_, _01130_);
  and _23494_ (_01134_, _01133_, _01125_);
  and _23495_ (_01136_, _09237_, _06452_);
  or _23496_ (_01137_, _01136_, _01134_);
  and _23497_ (_01139_, _01137_, _06474_);
  and _23498_ (_01140_, _01123_, _06491_);
  or _23499_ (_01141_, _01140_, _06498_);
  and _23500_ (_01142_, _09237_, _06483_);
  not _23501_ (_01143_, _06497_);
  and _23502_ (_01144_, _06480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23503_ (_01146_, _01144_, _06483_);
  and _23504_ (_01147_, _06478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23505_ (_01148_, _01147_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23506_ (_01150_, _01148_, _01146_);
  or _23507_ (_01151_, _01150_, _01143_);
  or _23508_ (_01153_, _01151_, _01142_);
  and _23509_ (_01155_, _01153_, _01141_);
  nand _23510_ (_01156_, _09237_, _06490_);
  nand _23511_ (_01158_, _01156_, _06519_);
  or _23512_ (_01159_, _01158_, _01155_);
  or _23513_ (_01160_, _06519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23514_ (_01161_, _01160_, _01159_);
  and _23515_ (_01163_, _01161_, _06564_);
  or _23516_ (_01164_, _01163_, _01139_);
  or _23517_ (_01165_, _01164_, _06508_);
  and _23518_ (_13475_, _01165_, _01122_);
  nor _23519_ (_01166_, _06562_, _06508_);
  not _23520_ (_01167_, _01166_);
  and _23521_ (_01168_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not _23522_ (_01169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23523_ (_01170_, _01126_, _01169_);
  nand _23524_ (_01171_, _01170_, _01129_);
  or _23525_ (_01172_, _09226_, _06471_);
  and _23526_ (_01173_, _01172_, _01171_);
  or _23527_ (_01174_, _01173_, _06457_);
  not _23528_ (_01176_, _06455_);
  not _23529_ (_01177_, _06457_);
  or _23530_ (_01178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23531_ (_01179_, _01178_, _01177_);
  and _23532_ (_01181_, _01179_, _01176_);
  and _23533_ (_01182_, _01181_, _01174_);
  and _23534_ (_01183_, _09226_, _06455_);
  or _23535_ (_01184_, _01183_, _06452_);
  or _23536_ (_01185_, _01184_, _01182_);
  or _23537_ (_01186_, _01178_, _06453_);
  and _23538_ (_01187_, _01186_, _06474_);
  and _23539_ (_01188_, _01187_, _01185_);
  or _23540_ (_01190_, _01178_, _06491_);
  and _23541_ (_01192_, _06519_, _06564_);
  or _23542_ (_01193_, _01147_, _01169_);
  nand _23543_ (_01194_, _01193_, _01146_);
  or _23544_ (_01195_, _09226_, _06484_);
  and _23545_ (_01197_, _01195_, _01194_);
  or _23546_ (_01198_, _01197_, _06494_);
  not _23547_ (_01200_, _06496_);
  not _23548_ (_01201_, _06494_);
  or _23549_ (_01203_, _01178_, _01201_);
  and _23550_ (_01204_, _01203_, _01200_);
  and _23551_ (_01205_, _01204_, _01198_);
  and _23552_ (_01206_, _09226_, _06496_);
  or _23553_ (_01207_, _01206_, _06490_);
  or _23554_ (_01208_, _01207_, _01205_);
  and _23555_ (_01209_, _01208_, _01192_);
  and _23556_ (_01210_, _01209_, _01190_);
  or _23557_ (_01211_, _01210_, _01188_);
  and _23558_ (_01212_, _01211_, _06509_);
  or _23559_ (_01213_, _01212_, _01168_);
  and _23560_ (_13478_, _01213_, _06071_);
  and _23561_ (_01214_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _23562_ (_01215_, _09576_, _06368_);
  or _23563_ (_01216_, _01215_, _01214_);
  and _23564_ (_13487_, _01216_, _06071_);
  nand _23565_ (_01217_, _00789_, _09341_);
  and _23566_ (_01218_, _00974_, _00916_);
  and _23567_ (_01219_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23568_ (_01220_, _01219_, _00786_);
  nor _23569_ (_01221_, _01220_, _01218_);
  and _23570_ (_01222_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23571_ (_01223_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23572_ (_01225_, _01223_, _01222_);
  or _23573_ (_01226_, _01225_, _00789_);
  and _23574_ (_01227_, _01226_, _00914_);
  and _23575_ (_01228_, _01227_, _01217_);
  and _23576_ (_01229_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23577_ (_01230_, _01229_, _01228_);
  and _23578_ (_13497_, _01230_, _06071_);
  nand _23579_ (_01231_, _01063_, _06609_);
  nor _23580_ (_01232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _23581_ (_01233_, _01232_);
  and _23582_ (_01234_, _01099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23583_ (_01235_, _01234_, _01233_);
  not _23584_ (_01237_, _01235_);
  nor _23585_ (_01238_, _01237_, _01035_);
  and _23586_ (_01239_, _01238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _23587_ (_01240_, _01238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor _23588_ (_01241_, _01240_, _01239_);
  nand _23589_ (_01242_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23590_ (_01243_, _01242_, _01035_);
  or _23591_ (_01244_, _01243_, _01241_);
  or _23592_ (_01245_, _01244_, _01063_);
  and _23593_ (_01246_, _01245_, _06071_);
  and _23594_ (_13502_, _01246_, _01231_);
  nand _23595_ (_01248_, _01063_, _09341_);
  not _23596_ (_01249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _23597_ (_01250_, _01035_, _01249_);
  and _23598_ (_01251_, _01232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23599_ (_01252_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23600_ (_01253_, _01252_, _01251_);
  and _23601_ (_01254_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _23602_ (_01255_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _23603_ (_01256_, _01047_, _01033_);
  and _23604_ (_01257_, _01256_, _01233_);
  or _23605_ (_01258_, _01257_, _01035_);
  and _23606_ (_01259_, _01258_, _01255_);
  or _23607_ (_01260_, _01259_, _01253_);
  and _23608_ (_01261_, _01260_, _01250_);
  or _23609_ (_01262_, _01261_, _01063_);
  and _23610_ (_01263_, _01262_, _06071_);
  and _23611_ (_13505_, _01263_, _01248_);
  nand _23612_ (_01264_, _01063_, _06993_);
  not _23613_ (_01265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand _23614_ (_01266_, _01035_, _01265_);
  and _23615_ (_01267_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23616_ (_01268_, _01099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _23617_ (_01269_, _01268_, _01234_);
  or _23618_ (_01270_, _01269_, _01267_);
  or _23619_ (_01271_, _01270_, _01035_);
  and _23620_ (_01272_, _01271_, _01266_);
  or _23621_ (_01273_, _01272_, _01063_);
  and _23622_ (_01274_, _01273_, _06071_);
  and _23623_ (_13508_, _01274_, _01264_);
  nor _23624_ (_01276_, _06508_, _06474_);
  or _23625_ (_01277_, _01276_, _06445_);
  nand _23626_ (_01279_, _00727_, _06562_);
  and _23627_ (_01280_, _01279_, _06071_);
  and _23628_ (_13517_, _01280_, _01277_);
  and _23629_ (_13520_, _07336_, _06071_);
  not _23630_ (_01281_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nor _23631_ (_01282_, _01166_, _01281_);
  or _23632_ (_01283_, _06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _23633_ (_01284_, _01283_, _06453_);
  and _23634_ (_01285_, _01284_, _06474_);
  and _23635_ (_01286_, _06467_, _06445_);
  nor _23636_ (_01287_, _01286_, _06470_);
  and _23637_ (_01288_, _06463_, _06445_);
  or _23638_ (_01290_, _01288_, _01281_);
  nand _23639_ (_01291_, _01290_, _01287_);
  or _23640_ (_01293_, _09225_, _06471_);
  and _23641_ (_01294_, _01293_, _01291_);
  or _23642_ (_01295_, _01294_, _06457_);
  or _23643_ (_01296_, _01283_, _01177_);
  and _23644_ (_01297_, _01296_, _01176_);
  and _23645_ (_01298_, _01297_, _01295_);
  and _23646_ (_01300_, _09225_, _06455_);
  or _23647_ (_01301_, _01300_, _06452_);
  or _23648_ (_01302_, _01301_, _01298_);
  and _23649_ (_01303_, _01302_, _01285_);
  or _23650_ (_01304_, _06494_, _06484_);
  and _23651_ (_01305_, _01304_, _01200_);
  or _23652_ (_01307_, _01305_, _09225_);
  and _23653_ (_01308_, _06480_, _06445_);
  nor _23654_ (_01309_, _01308_, _06483_);
  and _23655_ (_01310_, _06478_, _06445_);
  nor _23656_ (_01311_, _01310_, _01281_);
  nor _23657_ (_01312_, _01311_, _01143_);
  nand _23658_ (_01313_, _01312_, _01309_);
  and _23659_ (_01314_, _01313_, _01307_);
  or _23660_ (_01315_, _01314_, _06490_);
  or _23661_ (_01316_, _06496_, _01201_);
  and _23662_ (_01318_, _01316_, _06491_);
  or _23663_ (_01319_, _01318_, _01283_);
  and _23664_ (_01320_, _01319_, _01192_);
  and _23665_ (_01321_, _01320_, _01315_);
  or _23666_ (_01322_, _01321_, _01303_);
  and _23667_ (_01323_, _01322_, _06509_);
  or _23668_ (_01324_, _01323_, _01282_);
  and _23669_ (_13536_, _01324_, _06071_);
  and _23670_ (_01325_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _23671_ (_01326_, _06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23672_ (_01327_, _01326_, _06453_);
  or _23673_ (_01329_, _01327_, _06459_);
  or _23674_ (_01330_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23675_ (_01331_, _01330_, _01287_);
  nand _23676_ (_01332_, _09236_, _06470_);
  nand _23677_ (_01333_, _01332_, _06458_);
  or _23678_ (_01334_, _01333_, _01331_);
  and _23679_ (_01335_, _01334_, _01329_);
  and _23680_ (_01336_, _09236_, _06452_);
  or _23681_ (_01337_, _01336_, _01335_);
  and _23682_ (_01338_, _01337_, _06474_);
  and _23683_ (_01339_, _06497_, _06483_);
  or _23684_ (_01340_, _01339_, _06490_);
  and _23685_ (_01341_, _01340_, _09236_);
  or _23686_ (_01342_, _01326_, _06497_);
  and _23687_ (_01343_, _01342_, _06491_);
  or _23688_ (_01344_, _01310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23689_ (_01345_, _01344_, _01309_);
  or _23690_ (_01346_, _01345_, _01143_);
  and _23691_ (_01347_, _01346_, _01343_);
  or _23692_ (_01349_, _01347_, _01341_);
  and _23693_ (_01350_, _01349_, _01192_);
  or _23694_ (_01351_, _01350_, _01338_);
  and _23695_ (_01352_, _01351_, _06509_);
  or _23696_ (_01353_, _01352_, _01325_);
  and _23697_ (_13542_, _01353_, _06071_);
  nand _23698_ (_01354_, _01035_, _09341_);
  and _23699_ (_01355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23700_ (_01356_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23701_ (_01357_, _01356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23702_ (_01358_, _01357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23703_ (_01360_, _01358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23704_ (_01361_, _01360_, _01234_);
  nand _23705_ (_01362_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23706_ (_01363_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23707_ (_01364_, _01363_, _01232_);
  and _23708_ (_01365_, _01364_, _01362_);
  and _23709_ (_01366_, _01360_, _01088_);
  or _23710_ (_01368_, _01366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _23711_ (_01369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23712_ (_01370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _01369_);
  and _23713_ (_01371_, _01358_, _01088_);
  and _23714_ (_01372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23715_ (_01373_, _01372_, _01371_);
  not _23716_ (_01374_, _01373_);
  and _23717_ (_01375_, _01374_, _01370_);
  and _23718_ (_01376_, _01375_, _01368_);
  not _23719_ (_01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23720_ (_01378_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _23721_ (_01379_, _01378_, _01357_);
  and _23722_ (_01380_, _01379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand _23723_ (_01381_, _01380_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23724_ (_01382_, _01381_, _01377_);
  or _23725_ (_01383_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _23726_ (_01384_, _01372_);
  or _23727_ (_01385_, _01381_, _01384_);
  and _23728_ (_01386_, _01385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23729_ (_01387_, _01386_, _01383_);
  or _23730_ (_01388_, _01387_, _01376_);
  or _23731_ (_01389_, _01388_, _01365_);
  or _23732_ (_01390_, _01389_, _01035_);
  and _23733_ (_01391_, _01390_, _01098_);
  and _23734_ (_01392_, _01391_, _01354_);
  and _23735_ (_01393_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23736_ (_01394_, _01393_, _01392_);
  and _23737_ (_13545_, _01394_, _06071_);
  nand _23738_ (_01395_, _01035_, _06609_);
  or _23739_ (_01396_, _01370_, _01053_);
  and _23740_ (_01397_, _01371_, _01369_);
  nor _23741_ (_01398_, _01397_, _01377_);
  and _23742_ (_01399_, _01397_, _01377_);
  or _23743_ (_01400_, _01399_, _01398_);
  and _23744_ (_01401_, _01400_, _01396_);
  and _23745_ (_01402_, _01378_, _01358_);
  or _23746_ (_01403_, _01402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23747_ (_01404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _23748_ (_01405_, _01402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23749_ (_01406_, _01405_, _01404_);
  and _23750_ (_01407_, _01406_, _01403_);
  and _23751_ (_01409_, _01358_, _01234_);
  or _23752_ (_01410_, _01409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23753_ (_01411_, _01361_, _01233_);
  and _23754_ (_01412_, _01411_, _01410_);
  or _23755_ (_01413_, _01412_, _01407_);
  or _23756_ (_01414_, _01413_, _01401_);
  or _23757_ (_01415_, _01414_, _01035_);
  and _23758_ (_01416_, _01415_, _01098_);
  and _23759_ (_01417_, _01416_, _01395_);
  and _23760_ (_01418_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _23761_ (_01419_, _01418_, _01417_);
  and _23762_ (_13548_, _01419_, _06071_);
  nand _23763_ (_01420_, _01035_, _09037_);
  and _23764_ (_01421_, _01088_, _01369_);
  and _23765_ (_01422_, _01421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23766_ (_01423_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _23767_ (_01424_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23768_ (_01425_, _01424_, _01396_);
  and _23769_ (_01426_, _01425_, _01423_);
  not _23770_ (_01427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _23771_ (_01428_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23772_ (_01429_, _01428_, _01427_);
  and _23773_ (_01430_, _01355_, _01234_);
  nor _23774_ (_01431_, _01430_, _01233_);
  and _23775_ (_01432_, _01431_, _01429_);
  and _23776_ (_01433_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23777_ (_01434_, _01433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23778_ (_01435_, _01378_, _01355_);
  not _23779_ (_01436_, _01435_);
  and _23780_ (_01437_, _01436_, _01404_);
  and _23781_ (_01438_, _01437_, _01434_);
  or _23782_ (_01439_, _01438_, _01432_);
  or _23783_ (_01440_, _01439_, _01426_);
  or _23784_ (_01441_, _01440_, _01035_);
  and _23785_ (_01443_, _01441_, _01420_);
  or _23786_ (_01444_, _01443_, _01063_);
  nand _23787_ (_01445_, _01063_, _01427_);
  and _23788_ (_01446_, _01445_, _06071_);
  and _23789_ (_13561_, _01446_, _01444_);
  nand _23790_ (_01447_, _01035_, _06434_);
  or _23791_ (_01448_, _01430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23792_ (_01449_, _01356_, _01234_);
  nor _23793_ (_01450_, _01449_, _01233_);
  and _23794_ (_01451_, _01450_, _01448_);
  and _23795_ (_01452_, _01355_, _01088_);
  or _23796_ (_01453_, _01452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23797_ (_01454_, _01356_, _01088_);
  not _23798_ (_01455_, _01454_);
  and _23799_ (_01456_, _01455_, _01370_);
  and _23800_ (_01457_, _01456_, _01453_);
  and _23801_ (_01458_, _01435_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _23802_ (_01459_, _01458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23803_ (_01460_, _01378_, _01356_);
  nand _23804_ (_01462_, _01460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23805_ (_01463_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23806_ (_01465_, _01463_, _01459_);
  or _23807_ (_01466_, _01465_, _01457_);
  or _23808_ (_01467_, _01466_, _01451_);
  or _23809_ (_01468_, _01467_, _01035_);
  and _23810_ (_01469_, _01468_, _01098_);
  and _23811_ (_01470_, _01469_, _01447_);
  and _23812_ (_01471_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _23813_ (_01472_, _01471_, _01470_);
  and _23814_ (_13563_, _01472_, _06071_);
  and _23815_ (_01473_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23816_ (_01474_, _01473_, _01166_);
  and _23817_ (_13565_, _01474_, _06071_);
  nor _23818_ (_01475_, _06478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23819_ (_01476_, _01475_, _06480_);
  or _23820_ (_01477_, _01476_, _06483_);
  and _23821_ (_01478_, _01477_, _01201_);
  or _23822_ (_01479_, _01478_, _06496_);
  and _23823_ (_01480_, _01479_, _06491_);
  and _23824_ (_01481_, _01480_, _01192_);
  and _23825_ (_01482_, _06474_, _06453_);
  nor _23826_ (_01483_, _06463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23827_ (_01484_, _01483_, _06467_);
  or _23828_ (_01485_, _01484_, _06470_);
  and _23829_ (_01486_, _01485_, _01177_);
  or _23830_ (_01487_, _01486_, _06455_);
  and _23831_ (_01488_, _01487_, _01482_);
  or _23832_ (_01489_, _01488_, _06508_);
  or _23833_ (_01490_, _01489_, _01481_);
  or _23834_ (_01491_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23835_ (_01492_, _01491_, _06071_);
  and _23836_ (_13568_, _01492_, _01490_);
  nand _23837_ (_01493_, _01035_, _07945_);
  and _23838_ (_01494_, _01454_, _01369_);
  or _23839_ (_01495_, _01494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _23840_ (_01496_, _01494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23841_ (_01497_, _01496_, _01495_);
  and _23842_ (_01498_, _01497_, _01396_);
  or _23843_ (_01499_, _01449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23844_ (_01500_, _01357_, _01234_);
  nor _23845_ (_01502_, _01500_, _01233_);
  and _23846_ (_01503_, _01502_, _01499_);
  or _23847_ (_01504_, _01460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23848_ (_01506_, _01379_);
  and _23849_ (_01507_, _01506_, _01404_);
  and _23850_ (_01508_, _01507_, _01504_);
  or _23851_ (_01509_, _01508_, _01503_);
  or _23852_ (_01510_, _01509_, _01498_);
  or _23853_ (_01511_, _01510_, _01035_);
  and _23854_ (_01513_, _01511_, _01098_);
  and _23855_ (_01514_, _01513_, _01493_);
  and _23856_ (_01516_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _23857_ (_01518_, _01516_, _01514_);
  and _23858_ (_13571_, _01518_, _06071_);
  and _23859_ (_13573_, _10924_, _06508_);
  nand _23860_ (_01519_, _01035_, _06993_);
  and _23861_ (_01521_, _01357_, _01088_);
  or _23862_ (_01522_, _01521_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _23863_ (_01523_, _01371_);
  and _23864_ (_01524_, _01523_, _01370_);
  and _23865_ (_01525_, _01524_, _01522_);
  or _23866_ (_01526_, _01500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _23867_ (_01527_, _01409_, _01233_);
  and _23868_ (_01528_, _01527_, _01526_);
  or _23869_ (_01529_, _01380_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23870_ (_01530_, _01381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23871_ (_01531_, _01530_, _01529_);
  or _23872_ (_01532_, _01531_, _01528_);
  or _23873_ (_01533_, _01532_, _01525_);
  or _23874_ (_01534_, _01533_, _01035_);
  and _23875_ (_01535_, _01534_, _01098_);
  and _23876_ (_01536_, _01535_, _01519_);
  and _23877_ (_01537_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23878_ (_01538_, _01537_, _01536_);
  and _23879_ (_13575_, _01538_, _06071_);
  and _23880_ (_01539_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _23881_ (_01540_, _01539_, _01166_);
  and _23882_ (_13581_, _01540_, _06071_);
  nand _23883_ (_01541_, _01035_, _07977_);
  or _23884_ (_01542_, _01421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _23885_ (_01543_, _01422_);
  and _23886_ (_01544_, _01543_, _01396_);
  and _23887_ (_01545_, _01544_, _01542_);
  or _23888_ (_01546_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23889_ (_01547_, _01428_, _01232_);
  and _23890_ (_01548_, _01547_, _01546_);
  or _23891_ (_01549_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _23892_ (_01550_, _01433_);
  and _23893_ (_01551_, _01550_, _01404_);
  and _23894_ (_01552_, _01551_, _01549_);
  or _23895_ (_01553_, _01552_, _01548_);
  or _23896_ (_01554_, _01553_, _01545_);
  or _23897_ (_01555_, _01554_, _01035_);
  and _23898_ (_01556_, _01555_, _01541_);
  or _23899_ (_01557_, _01556_, _01063_);
  or _23900_ (_01558_, _01098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23901_ (_01559_, _01558_, _06071_);
  and _23902_ (_13591_, _01559_, _01557_);
  and _23903_ (_13596_, _11017_, _06508_);
  and _23904_ (_01560_, _13743_, _06840_);
  nand _23905_ (_01561_, _01560_, _07977_);
  or _23906_ (_01562_, _01560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23907_ (_01563_, _01562_, _06071_);
  and _23908_ (_13600_, _01563_, _01561_);
  nor _23909_ (_01564_, _06481_, _06488_);
  nand _23910_ (_01565_, _06517_, _01564_);
  nor _23911_ (_01566_, _01565_, _06474_);
  and _23912_ (_01567_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or _23913_ (_01568_, _06508_, _06470_);
  nor _23914_ (_01569_, _01568_, _06450_);
  not _23915_ (_01570_, _06468_);
  and _23916_ (_01571_, _01570_, _06459_);
  and _23917_ (_01573_, _01571_, _01569_);
  or _23918_ (_01574_, _01573_, _01567_);
  or _23919_ (_01576_, _01574_, _01566_);
  and _23920_ (_13601_, _01576_, _06071_);
  and _23921_ (_01577_, _12019_, _06369_);
  and _23922_ (_01578_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or _23923_ (_01579_, _01578_, _01577_);
  and _23924_ (_13605_, _01579_, _06071_);
  and _23925_ (_01581_, _13751_, _06840_);
  or _23926_ (_01582_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _23927_ (_01583_, _01582_, _06071_);
  nand _23928_ (_01584_, _01581_, _06434_);
  and _23929_ (_13607_, _01584_, _01583_);
  or _23930_ (_01585_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _23931_ (_01586_, _06530_, _05833_);
  and _23932_ (_01587_, _01586_, _06071_);
  and _23933_ (_13610_, _01587_, _01585_);
  or _23934_ (_01588_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _23935_ (_01589_, _01588_, _06071_);
  nand _23936_ (_01590_, _01581_, _07945_);
  and _23937_ (_13612_, _01590_, _01589_);
  nand _23938_ (_01591_, _01560_, _09037_);
  or _23939_ (_01592_, _01560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23940_ (_01593_, _01592_, _06071_);
  and _23941_ (_13615_, _01593_, _01591_);
  or _23942_ (_01594_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23943_ (_01595_, _01594_, _06071_);
  nand _23944_ (_01596_, _01581_, _06609_);
  and _23945_ (_13622_, _01596_, _01595_);
  or _23946_ (_01597_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23947_ (_01598_, _01597_, _06071_);
  nand _23948_ (_01599_, _01581_, _09341_);
  and _23949_ (_13624_, _01599_, _01598_);
  or _23950_ (_01600_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _23951_ (_01601_, _01600_, _06071_);
  nand _23952_ (_01602_, _01581_, _06993_);
  and _23953_ (_13626_, _01602_, _01601_);
  and _23954_ (_01603_, _12120_, _06369_);
  and _23955_ (_01604_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _23956_ (_01605_, _01604_, _01603_);
  and _23957_ (_13686_, _01605_, _06071_);
  nor _23958_ (_01606_, _05937_, _05923_);
  and _23959_ (_01607_, _01606_, _06820_);
  and _23960_ (_01608_, _01607_, _13722_);
  and _23961_ (_01609_, _13710_, _10943_);
  not _23962_ (_01610_, _01609_);
  or _23963_ (_01611_, _01610_, _10936_);
  and _23964_ (_01612_, _01611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _23965_ (_01613_, _01612_, _01608_);
  nor _23966_ (_01614_, _10930_, _06479_);
  or _23967_ (_01615_, _01614_, _10928_);
  and _23968_ (_01617_, _01615_, _01609_);
  or _23969_ (_01619_, _01617_, _01613_);
  nand _23970_ (_01621_, _01608_, _06993_);
  and _23971_ (_01622_, _01621_, _06071_);
  and _23972_ (_13768_, _01622_, _01619_);
  not _23973_ (_01623_, _01608_);
  and _23974_ (_01625_, _01609_, _07105_);
  or _23975_ (_01626_, _01625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _23976_ (_01627_, _01626_, _01623_);
  nand _23977_ (_01628_, _01625_, _06803_);
  and _23978_ (_01629_, _01628_, _01627_);
  nor _23979_ (_01630_, _01623_, _07945_);
  or _23980_ (_01631_, _01630_, _01629_);
  and _23981_ (_13773_, _01631_, _06071_);
  nor _23982_ (_01632_, _07753_, _06361_);
  or _23983_ (_01633_, _01610_, _01632_);
  and _23984_ (_01634_, _01633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23985_ (_01635_, _01634_, _01608_);
  and _23986_ (_01636_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23987_ (_01637_, _01636_, _00275_);
  and _23988_ (_01638_, _01637_, _01609_);
  or _23989_ (_01639_, _01638_, _01635_);
  nand _23990_ (_01640_, _01608_, _06434_);
  and _23991_ (_01641_, _01640_, _06071_);
  and _23992_ (_13775_, _01641_, _01639_);
  and _23993_ (_13787_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  and _23994_ (_01643_, _01609_, _08801_);
  or _23995_ (_01644_, _01643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _23996_ (_01645_, _01644_, _01623_);
  nand _23997_ (_01646_, _01643_, _06803_);
  and _23998_ (_01647_, _01646_, _01645_);
  nor _23999_ (_01649_, _01623_, _09341_);
  or _24000_ (_01650_, _01649_, _01647_);
  and _24001_ (_13795_, _01650_, _06071_);
  and _24002_ (_01652_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _24003_ (_01653_, _11023_, _06610_);
  or _24004_ (_01654_, _01653_, _01652_);
  and _24005_ (_13801_, _01654_, _06071_);
  and _24006_ (_01655_, _10948_, _06362_);
  or _24007_ (_01656_, _01655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _24008_ (_01657_, _01656_, _10953_);
  nand _24009_ (_01659_, _01655_, _06803_);
  and _24010_ (_01660_, _01659_, _01657_);
  nor _24011_ (_01661_, _10953_, _09037_);
  or _24012_ (_01662_, _01661_, _01660_);
  and _24013_ (_13834_, _01662_, _06071_);
  and _24014_ (_01664_, _10948_, _06383_);
  and _24015_ (_01665_, _01664_, _06803_);
  nor _24016_ (_01666_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _24017_ (_01667_, _01666_, _01665_);
  nand _24018_ (_01668_, _01667_, _10953_);
  nand _24019_ (_01669_, _10952_, _07977_);
  and _24020_ (_01670_, _01669_, _06071_);
  and _24021_ (_13841_, _01670_, _01668_);
  and _24022_ (_01671_, _10948_, _08801_);
  and _24023_ (_01672_, _01671_, _06803_);
  nor _24024_ (_01674_, _01671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _24025_ (_01675_, _01674_, _01672_);
  nand _24026_ (_01676_, _01675_, _10953_);
  nand _24027_ (_01677_, _10952_, _09341_);
  and _24028_ (_01678_, _01677_, _06071_);
  and _24029_ (_13855_, _01678_, _01676_);
  or _24030_ (_01680_, _05993_, _05981_);
  nand _24031_ (_01681_, _01680_, _10948_);
  and _24032_ (_01682_, _01681_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _24033_ (_01683_, _01682_, _10952_);
  or _24034_ (_01684_, _06005_, _05981_);
  and _24035_ (_01685_, _01684_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _24036_ (_01686_, _01685_, _08943_);
  and _24037_ (_01687_, _01686_, _10948_);
  or _24038_ (_01688_, _01687_, _01683_);
  nand _24039_ (_01689_, _10952_, _06609_);
  and _24040_ (_01690_, _01689_, _06071_);
  and _24041_ (_13859_, _01690_, _01688_);
  not _24042_ (_01691_, _10948_);
  or _24043_ (_01692_, _01691_, _10936_);
  and _24044_ (_01693_, _01692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _24045_ (_01694_, _01693_, _10952_);
  nor _24046_ (_01695_, _10930_, _06464_);
  or _24047_ (_01696_, _01695_, _10928_);
  and _24048_ (_01697_, _01696_, _10948_);
  or _24049_ (_01698_, _01697_, _01694_);
  nand _24050_ (_01699_, _10952_, _06993_);
  and _24051_ (_01700_, _01699_, _06071_);
  and _24052_ (_13862_, _01700_, _01698_);
  and _24053_ (_01701_, _10948_, _07105_);
  or _24054_ (_01702_, _01701_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _24055_ (_01703_, _01702_, _10953_);
  nand _24056_ (_01704_, _01701_, _06803_);
  and _24057_ (_01706_, _01704_, _01703_);
  nor _24058_ (_01707_, _10953_, _07945_);
  or _24059_ (_01708_, _01707_, _01706_);
  and _24060_ (_13868_, _01708_, _06071_);
  nor _24061_ (_13941_, _12084_, rst);
  nand _24062_ (_13965_, _12397_, _06071_);
  nor _24063_ (_13984_, _12098_, rst);
  nor _24064_ (_13989_, _12142_, rst);
  nor _24065_ (_13992_, _12212_, rst);
  and _24066_ (_13995_, _11961_, _06071_);
  nand _24067_ (_14001_, _12378_, _06071_);
  and _24068_ (_00014_, _07342_, _06071_);
  and _24069_ (_00186_, _08028_, _06071_);
  and _24070_ (_00258_, t2ex_i, _06071_);
  and _24071_ (_01709_, _09348_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand _24072_ (_01710_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _24073_ (_01711_, _01710_, _09346_);
  nor _24074_ (_01712_, _06609_, _06400_);
  or _24075_ (_01713_, _01712_, _01711_);
  or _24076_ (_01714_, _01713_, _01709_);
  and _24077_ (_00264_, _01714_, _06071_);
  and _24078_ (_00321_, _12076_, _06071_);
  and _24079_ (_00359_, _07781_, _06071_);
  nor _24080_ (_01715_, _12274_, _11403_);
  nor _24081_ (_01717_, _01715_, _11795_);
  or _24082_ (_01718_, _11876_, _11869_);
  or _24083_ (_01720_, _01718_, _12268_);
  or _24084_ (_01721_, _11845_, _11828_);
  or _24085_ (_01722_, _11881_, _11865_);
  or _24086_ (_01723_, _01722_, _01721_);
  or _24087_ (_01724_, _01723_, _01720_);
  or _24088_ (_01725_, _01724_, _11843_);
  and _24089_ (_01726_, _01725_, _11421_);
  or _24090_ (_01727_, _01726_, _01717_);
  and _24091_ (_00388_, _01727_, _06071_);
  and _24092_ (_01728_, _09228_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _24093_ (_01729_, _09239_, _09233_);
  nand _24094_ (_01731_, _01729_, _01728_);
  nand _24095_ (_01733_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _24096_ (_01735_, _01733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _24097_ (_01737_, _06840_, _06380_);
  nor _24098_ (_01738_, _01737_, _10945_);
  or _24099_ (_01740_, _01738_, _01735_);
  nand _24100_ (_01741_, _01738_, _08799_);
  and _24101_ (_01742_, _01741_, _01740_);
  nand _24102_ (_01744_, _01742_, _09250_);
  nand _24103_ (_01745_, _09249_, _09037_);
  and _24104_ (_01746_, _01745_, _06071_);
  and _24105_ (_00430_, _01746_, _01744_);
  nand _24106_ (_01747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _24107_ (_01748_, _01728_, _09240_);
  nor _24108_ (_01749_, _01748_, _01747_);
  and _24109_ (_01750_, _07105_, _06378_);
  nand _24110_ (_01751_, _01750_, _06840_);
  or _24111_ (_01752_, _01751_, _10945_);
  nand _24112_ (_01753_, _01752_, _01749_);
  or _24113_ (_01754_, _01752_, _06803_);
  and _24114_ (_01755_, _01754_, _01753_);
  nand _24115_ (_01757_, _01755_, _09250_);
  nand _24116_ (_01758_, _09249_, _07945_);
  and _24117_ (_01759_, _01758_, _06071_);
  and _24118_ (_00433_, _01759_, _01757_);
  and _24119_ (_01760_, _01609_, _06805_);
  or _24120_ (_01761_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _24121_ (_01762_, _01761_, _01623_);
  nand _24122_ (_01764_, _01760_, _06803_);
  and _24123_ (_01765_, _01764_, _01762_);
  nor _24124_ (_01766_, _01623_, _06359_);
  or _24125_ (_01767_, _01766_, _01765_);
  and _24126_ (_00470_, _01767_, _06071_);
  and _24127_ (_01768_, _01068_, _06805_);
  and _24128_ (_01769_, _01768_, _06840_);
  and _24129_ (_01770_, _01769_, _06803_);
  and _24130_ (_01771_, _09238_, _09233_);
  nand _24131_ (_01772_, _01771_, _09229_);
  nand _24132_ (_01773_, _01772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand _24133_ (_01774_, _01773_, _07876_);
  nor _24134_ (_01775_, _01774_, _01769_);
  or _24135_ (_01776_, _01775_, _01770_);
  nand _24136_ (_01777_, _01776_, _09250_);
  nand _24137_ (_01778_, _09249_, _06359_);
  and _24138_ (_01779_, _01778_, _06071_);
  and _24139_ (_00475_, _01779_, _01777_);
  and _24140_ (_00531_, _11392_, _06071_);
  nor _24141_ (_00563_, _11533_, rst);
  and _24142_ (_00574_, _00646_, _06071_);
  and _24143_ (_01780_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08003_);
  and _24144_ (_01781_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _24145_ (_01782_, _01781_, _01780_);
  and _24146_ (_00592_, _01782_, _06071_);
  and _24147_ (_01783_, _07824_, _06809_);
  nand _24148_ (_01784_, _01783_, _06383_);
  or _24149_ (_01785_, _01784_, _00593_);
  not _24150_ (_01786_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _24151_ (_01787_, _01784_, _01786_);
  and _24152_ (_01788_, _01787_, _06012_);
  and _24153_ (_01789_, _01788_, _01785_);
  nor _24154_ (_01790_, _06814_, _01786_);
  not _24155_ (_01791_, _01783_);
  or _24156_ (_01792_, _01791_, _10936_);
  and _24157_ (_01793_, _01792_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor _24158_ (_01794_, _10930_, _01786_);
  or _24159_ (_01795_, _01794_, _10928_);
  and _24160_ (_01796_, _01795_, _01783_);
  or _24161_ (_01797_, _01796_, _01793_);
  and _24162_ (_01798_, _01797_, _06815_);
  or _24163_ (_01799_, _01798_, _01790_);
  or _24164_ (_01800_, _01799_, _01789_);
  and _24165_ (_00618_, _01800_, _06071_);
  or _24166_ (_01801_, _01784_, _00612_);
  not _24167_ (_01802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _24168_ (_01803_, _01784_, _01802_);
  and _24169_ (_01804_, _01803_, _06012_);
  and _24170_ (_01805_, _01804_, _01801_);
  nor _24171_ (_01806_, _06814_, _01802_);
  and _24172_ (_01807_, _01783_, _07105_);
  nand _24173_ (_01808_, _01807_, _06803_);
  or _24174_ (_01809_, _01807_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _24175_ (_01810_, _01809_, _06815_);
  and _24176_ (_01811_, _01810_, _01808_);
  or _24177_ (_01812_, _01811_, _01806_);
  or _24178_ (_01813_, _01812_, _01805_);
  and _24179_ (_00621_, _01813_, _06071_);
  or _24180_ (_01814_, _01784_, _07425_);
  not _24181_ (_01815_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _24182_ (_01817_, _01784_, _01815_);
  and _24183_ (_01818_, _01817_, _06012_);
  and _24184_ (_01819_, _01818_, _01814_);
  nor _24185_ (_01820_, _06814_, _01815_);
  and _24186_ (_01821_, _01783_, _08801_);
  nand _24187_ (_01822_, _01821_, _06803_);
  or _24188_ (_01823_, _01821_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _24189_ (_01824_, _01823_, _06815_);
  and _24190_ (_01825_, _01824_, _01822_);
  or _24191_ (_01826_, _01825_, _01820_);
  or _24192_ (_01827_, _01826_, _01819_);
  and _24193_ (_00641_, _01827_, _06071_);
  and _24194_ (pc_log_change, _08705_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _24195_ (_01828_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _24196_ (_01830_, pc_log_change, _06086_);
  and _24197_ (_01831_, _01830_, _06071_);
  and _24198_ (_00725_, _01831_, _01828_);
  and _24199_ (_01832_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08003_);
  and _24200_ (_01833_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _24201_ (_01834_, _01833_, _01832_);
  and _24202_ (_00728_, _01834_, _06071_);
  and _24203_ (_01836_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _24204_ (_01837_, _07945_, _06611_);
  or _24205_ (_01838_, _01837_, _01836_);
  and _24206_ (_00781_, _01838_, _06071_);
  and _24207_ (_01839_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _24208_ (_01840_, _06611_, _06359_);
  or _24209_ (_01841_, _01840_, _01839_);
  and _24210_ (_00826_, _01841_, _06071_);
  nor _24211_ (_00864_, _11965_, rst);
  nand _24212_ (_01842_, _07977_, _07946_);
  or _24213_ (_01843_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _24214_ (_01844_, _01843_, _01842_);
  and _24215_ (_00872_, _01844_, _06071_);
  or _24216_ (_01845_, _01784_, _00655_);
  not _24217_ (_01846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _24218_ (_01847_, _01784_, _01846_);
  and _24219_ (_01848_, _01847_, _06012_);
  and _24220_ (_01849_, _01848_, _01845_);
  nor _24221_ (_01850_, _06814_, _01846_);
  and _24222_ (_01852_, _01783_, _06362_);
  nand _24223_ (_01853_, _01852_, _06803_);
  or _24224_ (_01854_, _01852_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _24225_ (_01855_, _01854_, _06815_);
  and _24226_ (_01856_, _01855_, _01853_);
  or _24227_ (_01857_, _01856_, _01850_);
  or _24228_ (_01858_, _01857_, _01849_);
  and _24229_ (_00886_, _01858_, _06071_);
  or _24230_ (_01859_, _01784_, _00660_);
  not _24231_ (_01860_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _24232_ (_01861_, _01784_, _01860_);
  and _24233_ (_01862_, _01861_, _06012_);
  and _24234_ (_01863_, _01862_, _01859_);
  nor _24235_ (_01864_, _06814_, _01860_);
  or _24236_ (_01865_, _01784_, _08799_);
  and _24237_ (_01866_, _01861_, _06815_);
  and _24238_ (_01867_, _01866_, _01865_);
  or _24239_ (_01868_, _01867_, _01864_);
  or _24240_ (_01869_, _01868_, _01863_);
  and _24241_ (_00897_, _01869_, _06071_);
  or _24242_ (_01871_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not _24243_ (_01872_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _24244_ (_01873_, pc_log_change, _01872_);
  and _24245_ (_01874_, _01873_, _06071_);
  and _24246_ (_00999_, _01874_, _01871_);
  or _24247_ (_01875_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not _24248_ (_01876_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _24249_ (_01877_, pc_log_change, _01876_);
  and _24250_ (_01878_, _01877_, _06071_);
  and _24251_ (_01002_, _01878_, _01875_);
  or _24252_ (_01879_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not _24253_ (_01880_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _24254_ (_01881_, pc_log_change, _01880_);
  and _24255_ (_01882_, _01881_, _06071_);
  and _24256_ (_01006_, _01882_, _01879_);
  and _24257_ (_01883_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _24258_ (_01884_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _24259_ (_01885_, pc_log_change, _01884_);
  or _24260_ (_01886_, _01885_, _01883_);
  and _24261_ (_01009_, _01886_, _06071_);
  not _24262_ (_01887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _24263_ (_01888_, _06062_, _01887_);
  or _24264_ (_01889_, _01888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _24265_ (_01891_, _10947_, _09026_);
  or _24266_ (_01892_, _01891_, _01889_);
  not _24267_ (_01893_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _24268_ (_01894_, _08801_, _01893_);
  nand _24269_ (_01895_, _01894_, _01891_);
  or _24270_ (_01896_, _01895_, _08802_);
  and _24271_ (_01897_, _01896_, _01892_);
  and _24272_ (_01898_, _09248_, _05969_);
  or _24273_ (_01899_, _01898_, _01897_);
  nand _24274_ (_01900_, _01898_, _09341_);
  and _24275_ (_01901_, _01900_, _06071_);
  and _24276_ (_01013_, _01901_, _01899_);
  not _24277_ (_01903_, _01898_);
  and _24278_ (_01904_, _01891_, _06032_);
  or _24279_ (_01905_, _01904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _24280_ (_01906_, _01905_, _01903_);
  nand _24281_ (_01907_, _01904_, _06803_);
  and _24282_ (_01908_, _01907_, _01906_);
  nor _24283_ (_01909_, _01903_, _06609_);
  or _24284_ (_01910_, _01909_, _01908_);
  and _24285_ (_01015_, _01910_, _06071_);
  not _24286_ (_01911_, _01891_);
  or _24287_ (_01912_, _01911_, _10936_);
  and _24288_ (_01913_, _01912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _24289_ (_01915_, _01913_, _01898_);
  not _24290_ (_01916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor _24291_ (_01917_, _10930_, _01916_);
  or _24292_ (_01918_, _01917_, _10928_);
  and _24293_ (_01919_, _01918_, _01891_);
  or _24294_ (_01920_, _01919_, _01915_);
  nand _24295_ (_01921_, _01898_, _06993_);
  and _24296_ (_01922_, _01921_, _06071_);
  and _24297_ (_01019_, _01922_, _01920_);
  nor _24298_ (_01923_, _01035_, rst);
  and _24299_ (_01924_, _01034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _24300_ (_01925_, _01372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24301_ (_01926_, _01925_, _01358_);
  nand _24302_ (_01927_, _01926_, _01234_);
  and _24303_ (_01928_, _01927_, _01232_);
  or _24304_ (_01929_, _01926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _24305_ (_01930_, _01929_, _01088_);
  nor _24306_ (_01931_, _01930_, _01232_);
  nor _24307_ (_01932_, _01931_, _01928_);
  nor _24308_ (_01933_, _01932_, _01924_);
  nor _24309_ (_01934_, _01933_, _01063_);
  and _24310_ (_01024_, _01934_, _01923_);
  and _24311_ (_01935_, _01373_, _01369_);
  or _24312_ (_01936_, _01935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24313_ (_01937_, _01925_, _01397_);
  and _24314_ (_01938_, _01937_, _01396_);
  and _24315_ (_01939_, _01938_, _01936_);
  not _24316_ (_01940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24317_ (_01941_, _01362_, _01940_);
  and _24318_ (_01942_, _01941_, _01928_);
  and _24319_ (_01943_, _01402_, _01372_);
  or _24320_ (_01944_, _01943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24321_ (_01945_, _01925_, _01402_);
  not _24322_ (_01946_, _01945_);
  and _24323_ (_01947_, _01946_, _01404_);
  and _24324_ (_01948_, _01947_, _01944_);
  or _24325_ (_01949_, _01948_, _01942_);
  nor _24326_ (_01950_, _01949_, _01939_);
  nor _24327_ (_01951_, _01950_, _01035_);
  and _24328_ (_01952_, _01035_, _06360_);
  or _24329_ (_01953_, _01952_, _01951_);
  and _24330_ (_01954_, _01953_, _01098_);
  and _24331_ (_01955_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24332_ (_01956_, _01955_, _01954_);
  and _24333_ (_01026_, _01956_, _06071_);
  nand _24334_ (_01957_, _01063_, _06359_);
  and _24335_ (_01958_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _24336_ (_01959_, _01958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _24337_ (_01960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01369_);
  nand _24338_ (_01961_, _01960_, _01051_);
  nand _24339_ (_01962_, _01961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _24340_ (_01963_, _01962_, _01256_);
  or _24341_ (_01964_, _01963_, _01035_);
  and _24342_ (_01965_, _01964_, _01959_);
  or _24343_ (_01966_, _01965_, _01063_);
  and _24344_ (_01967_, _01966_, _06071_);
  and _24345_ (_01028_, _01967_, _01957_);
  and _24346_ (_01968_, _01891_, _07105_);
  or _24347_ (_01969_, _01968_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _24348_ (_01970_, _01969_, _01903_);
  nand _24349_ (_01971_, _01968_, _06803_);
  and _24350_ (_01972_, _01971_, _01970_);
  nor _24351_ (_01973_, _01903_, _07945_);
  or _24352_ (_01974_, _01973_, _01972_);
  and _24353_ (_01036_, _01974_, _06071_);
  or _24354_ (_01975_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _24355_ (_01976_, _01975_, _06071_);
  nand _24356_ (_01977_, _01581_, _06359_);
  and _24357_ (_01039_, _01977_, _01976_);
  or _24358_ (_01978_, _01911_, _01632_);
  and _24359_ (_01979_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _24360_ (_01980_, _01979_, _01898_);
  and _24361_ (_01981_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _24362_ (_01982_, _01981_, _00275_);
  and _24363_ (_01983_, _01982_, _01891_);
  or _24364_ (_01984_, _01983_, _01980_);
  nand _24365_ (_01985_, _01898_, _06434_);
  and _24366_ (_01986_, _01985_, _06071_);
  and _24367_ (_01042_, _01986_, _01984_);
  or _24368_ (_01987_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _24369_ (_01988_, pc_log_change, _06243_);
  and _24370_ (_01989_, _01988_, _06071_);
  and _24371_ (_01045_, _01989_, _01987_);
  not _24372_ (_01990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _24373_ (_01991_, _01378_, _01990_);
  or _24374_ (_01992_, _01991_, _01945_);
  nand _24375_ (_01993_, _01992_, _01404_);
  nor _24376_ (_01994_, _01993_, _01063_);
  and _24377_ (_01049_, _01994_, _01923_);
  and _24378_ (_01995_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _24379_ (_01996_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _24380_ (_01997_, pc_log_change, _01996_);
  or _24381_ (_01998_, _01997_, _01995_);
  and _24382_ (_01052_, _01998_, _06071_);
  and _24383_ (_01999_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _24384_ (_02000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _24385_ (_02001_, pc_log_change, _02000_);
  or _24386_ (_02002_, _02001_, _01999_);
  and _24387_ (_01056_, _02002_, _06071_);
  and _24388_ (_02003_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _24389_ (_02004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _24390_ (_02005_, pc_log_change, _02004_);
  or _24391_ (_02006_, _02005_, _02003_);
  and _24392_ (_01059_, _02006_, _06071_);
  and _24393_ (_01067_, t0_i, _06071_);
  nand _24394_ (_02007_, _00762_, _06359_);
  not _24395_ (_02008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24396_ (_02009_, _00790_, _02008_);
  or _24397_ (_02010_, _00780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24398_ (_02011_, _00797_, _00787_);
  and _24399_ (_02012_, _02011_, _02010_);
  and _24400_ (_02013_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _24401_ (_02014_, _02013_, _02012_);
  nor _24402_ (_02015_, _02014_, _00789_);
  or _24403_ (_02016_, _02015_, _02009_);
  or _24404_ (_02017_, _02016_, _00762_);
  and _24405_ (_02018_, _02017_, _06071_);
  and _24406_ (_01071_, _02018_, _02007_);
  not _24407_ (_02019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _24408_ (_02020_, _00772_, _02019_);
  and _24409_ (_02021_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24410_ (_02022_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _24411_ (_02023_, _00965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _24412_ (_02024_, _02023_, _02022_);
  and _24413_ (_02026_, _02024_, _02021_);
  or _24414_ (_02027_, _02026_, _02020_);
  and _24415_ (_02028_, _02027_, _00916_);
  and _24416_ (_02029_, _02021_, _02023_);
  and _24417_ (_02030_, _02029_, _00945_);
  or _24418_ (_02031_, _02030_, _02020_);
  and _24419_ (_02032_, _02031_, _00786_);
  nand _24420_ (_02033_, _00772_, _00783_);
  and _24421_ (_02034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _24422_ (_02035_, _02034_, _02033_);
  or _24423_ (_02036_, _02035_, _02032_);
  or _24424_ (_02037_, _02036_, _00798_);
  or _24425_ (_02038_, _02037_, _02028_);
  nand _24426_ (_02039_, _02038_, _06071_);
  nor _24427_ (_02040_, _02039_, _00860_);
  and _24428_ (_01073_, _02040_, _01000_);
  nand _24429_ (_02042_, _00789_, _06359_);
  nand _24430_ (_02043_, _01220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _24431_ (_02044_, _00916_, _00772_);
  and _24432_ (_02045_, _02044_, _02023_);
  nand _24433_ (_02046_, _02045_, _02022_);
  and _24434_ (_02047_, _02046_, _02043_);
  nor _24435_ (_02048_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24436_ (_02049_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24437_ (_02050_, _02049_, _02048_);
  or _24438_ (_02051_, _02050_, _00789_);
  and _24439_ (_02052_, _02051_, _00914_);
  and _24440_ (_02053_, _02052_, _02042_);
  and _24441_ (_02054_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24442_ (_02055_, _02054_, _02053_);
  and _24443_ (_01075_, _02055_, _06071_);
  and _24444_ (_01078_, t1_i, _06071_);
  and _24445_ (_02056_, _01891_, _06362_);
  or _24446_ (_02057_, _02056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _24447_ (_02058_, _02057_, _01903_);
  nand _24448_ (_02059_, _02056_, _06803_);
  and _24449_ (_02060_, _02059_, _02058_);
  nor _24450_ (_02061_, _01903_, _09037_);
  or _24451_ (_02062_, _02061_, _02060_);
  and _24452_ (_01083_, _02062_, _06071_);
  and _24453_ (_02063_, _01891_, _06383_);
  or _24454_ (_02064_, _02063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _24455_ (_02065_, _02064_, _01903_);
  nand _24456_ (_02066_, _02063_, _06803_);
  and _24457_ (_02067_, _02066_, _02065_);
  and _24458_ (_02068_, _01898_, _07978_);
  or _24459_ (_02069_, _02068_, _02067_);
  and _24460_ (_01086_, _02069_, _06071_);
  or _24461_ (_02070_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _24462_ (_02071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _24463_ (_02072_, pc_log_change, _02071_);
  and _24464_ (_02073_, _02072_, _06071_);
  and _24465_ (_01135_, _02073_, _02070_);
  or _24466_ (_02075_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not _24467_ (_02076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _24468_ (_02077_, pc_log_change, _02076_);
  and _24469_ (_02078_, _02077_, _06071_);
  and _24470_ (_01138_, _02078_, _02075_);
  and _24471_ (_02079_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _24472_ (_02081_, pc_log_change, _01872_);
  or _24473_ (_02082_, _02081_, _02079_);
  and _24474_ (_01145_, _02082_, _06071_);
  nand _24475_ (_02083_, _09341_, _06035_);
  or _24476_ (_02084_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _24477_ (_02085_, _06541_, _06065_);
  and _24478_ (_02086_, _02085_, _02084_);
  or _24479_ (_02087_, _06548_, _06065_);
  and _24480_ (_02088_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _24481_ (_02089_, _02088_, _02086_);
  nand _24482_ (_02090_, _02089_, _06036_);
  not _24483_ (_02091_, _06029_);
  or _24484_ (_02092_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _24485_ (_02093_, _02092_, _06071_);
  and _24486_ (_02095_, _02093_, _02090_);
  and _24487_ (_01149_, _02095_, _02083_);
  and _24488_ (_02096_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _24489_ (_02097_, pc_log_change, _01880_);
  or _24490_ (_02098_, _02097_, _02096_);
  and _24491_ (_01152_, _02098_, _06071_);
  and _24492_ (_02100_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not _24493_ (_02101_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand _24494_ (_02102_, _06065_, _02101_);
  not _24495_ (_02103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _24496_ (_02105_, _06538_, _06045_);
  and _24497_ (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _24498_ (_02107_, _02106_, _02103_);
  nor _24499_ (_02108_, _02106_, _02103_);
  and _24500_ (_02109_, _06548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _24501_ (_02110_, _02109_, _06065_);
  or _24502_ (_02111_, _02110_, _02108_);
  or _24503_ (_02112_, _02111_, _02107_);
  and _24504_ (_02113_, _02112_, _02102_);
  and _24505_ (_02114_, _02113_, _06036_);
  or _24506_ (_02115_, _02114_, _02100_);
  nor _24507_ (_02116_, _06609_, _06555_);
  or _24508_ (_02117_, _02116_, _02115_);
  and _24509_ (_01154_, _02117_, _06071_);
  nand _24510_ (_02118_, _06993_, _06035_);
  or _24511_ (_02119_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _24512_ (_02120_, _02106_, _06065_);
  and _24513_ (_02121_, _02120_, _02119_);
  and _24514_ (_02122_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _24515_ (_02123_, _02122_, _02121_);
  nand _24516_ (_02124_, _02123_, _06036_);
  or _24517_ (_02125_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _24518_ (_02126_, _02125_, _06071_);
  and _24519_ (_02127_, _02126_, _02124_);
  and _24520_ (_01157_, _02127_, _02118_);
  and _24521_ (_02128_, _06044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _24522_ (_02129_, _02128_, _06059_);
  and _24523_ (_02130_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _24524_ (_02131_, _02130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor _24525_ (_02132_, _02105_, _06065_);
  and _24526_ (_02133_, _02132_, _02131_);
  and _24527_ (_02134_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _24528_ (_02135_, _02134_, _02133_);
  nand _24529_ (_02136_, _02135_, _06036_);
  nand _24530_ (_02137_, _07945_, _06035_);
  or _24531_ (_02138_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _24532_ (_02139_, _02138_, _06071_);
  and _24533_ (_02140_, _02139_, _02137_);
  and _24534_ (_01162_, _02140_, _02136_);
  and _24535_ (_02141_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _24536_ (_02142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _24537_ (_02143_, pc_log_change, _02142_);
  or _24538_ (_02144_, _02143_, _02141_);
  and _24539_ (_01175_, _02144_, _06071_);
  and _24540_ (_02145_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24541_ (_02146_, pc_log_change, _02071_);
  or _24542_ (_02147_, _02146_, _02145_);
  and _24543_ (_01180_, _02147_, _06071_);
  and _24544_ (_02148_, _11023_, _08864_);
  and _24545_ (_02150_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _24546_ (_02151_, _02150_, _02148_);
  and _24547_ (_01189_, _02151_, _06071_);
  nor _24548_ (_02152_, _06538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _24549_ (_02153_, _02152_, _02130_);
  and _24550_ (_02154_, _02153_, _06066_);
  and _24551_ (_02155_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _24552_ (_02156_, _02155_, _02154_);
  nand _24553_ (_02157_, _02156_, _06036_);
  nand _24554_ (_02158_, _06434_, _06035_);
  or _24555_ (_02159_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _24556_ (_02160_, _02159_, _06071_);
  and _24557_ (_02161_, _02160_, _02158_);
  and _24558_ (_01191_, _02161_, _02157_);
  and _24559_ (_02162_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _24560_ (_02163_, _06537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _24561_ (_02164_, _06538_, _06065_);
  and _24562_ (_02165_, _02164_, _02163_);
  nor _24563_ (_02166_, _02165_, _02162_);
  nand _24564_ (_02167_, _02166_, _06036_);
  nand _24565_ (_02168_, _09037_, _06035_);
  or _24566_ (_02169_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _24567_ (_02170_, _02169_, _06071_);
  and _24568_ (_02171_, _02170_, _02168_);
  and _24569_ (_01196_, _02171_, _02167_);
  or _24570_ (_02172_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _24571_ (_02173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _24572_ (_02174_, pc_log_change, _02173_);
  and _24573_ (_02176_, _02174_, _06071_);
  and _24574_ (_01199_, _02176_, _02172_);
  and _24575_ (_02177_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _24576_ (_02178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _24577_ (_02179_, pc_log_change, _02178_);
  or _24578_ (_02180_, _02179_, _02177_);
  and _24579_ (_01202_, _02180_, _06071_);
  or _24580_ (_02181_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _24581_ (_02182_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _24582_ (_02183_, _02182_, _06547_);
  and _24583_ (_02184_, _06059_, _06043_);
  nor _24584_ (_02185_, _02184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor _24585_ (_02187_, _02185_, _06537_);
  or _24586_ (_02188_, _02187_, _06065_);
  or _24587_ (_02189_, _02188_, _02183_);
  and _24588_ (_02190_, _02189_, _02181_);
  and _24589_ (_02191_, _02190_, _06036_);
  and _24590_ (_02192_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _24591_ (_02193_, _00788_, _05969_);
  and _24592_ (_02194_, _07978_, _02193_);
  or _24593_ (_02195_, _02194_, _02192_);
  or _24594_ (_02196_, _02195_, _02191_);
  and _24595_ (_01224_, _02196_, _06071_);
  nor _24596_ (_02198_, _08865_, _06434_);
  and _24597_ (_02199_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or _24598_ (_02200_, _02199_, _02198_);
  and _24599_ (_01236_, _02200_, _06071_);
  and _24600_ (_02201_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _24601_ (_02202_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  or _24602_ (_02203_, _02202_, _02201_);
  and _24603_ (_01247_, _02203_, _06071_);
  nor _24604_ (_02204_, _06609_, _02091_);
  not _24605_ (_02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _24606_ (_02206_, _06059_, _06040_);
  nor _24607_ (_02207_, _02206_, _02205_);
  and _24608_ (_02208_, _02206_, _02205_);
  or _24609_ (_02209_, _02208_, _02207_);
  and _24610_ (_02210_, _02209_, _06066_);
  and _24611_ (_02211_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _24612_ (_02212_, _02211_, _02210_);
  and _24613_ (_02213_, _02212_, _06036_);
  and _24614_ (_02214_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _24615_ (_02215_, _02214_, _02213_);
  or _24616_ (_02216_, _02215_, _02204_);
  and _24617_ (_01275_, _02216_, _06071_);
  nor _24618_ (_01278_, _11591_, rst);
  nor _24619_ (_02217_, _09341_, _02091_);
  or _24620_ (_02218_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _24621_ (_02219_, _06041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _24622_ (_02220_, _06059_, _06042_);
  and _24623_ (_02221_, _02220_, _02219_);
  and _24624_ (_02222_, _06547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _24625_ (_02223_, _02222_, _02221_);
  and _24626_ (_02224_, _02223_, _02218_);
  or _24627_ (_02225_, _02224_, _06065_);
  not _24628_ (_02226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand _24629_ (_02227_, _06065_, _02226_);
  and _24630_ (_02228_, _02227_, _02225_);
  and _24631_ (_02229_, _02228_, _06036_);
  and _24632_ (_02230_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _24633_ (_02231_, _02230_, _02229_);
  or _24634_ (_02232_, _02231_, _02217_);
  and _24635_ (_01289_, _02232_, _06071_);
  nor _24636_ (_02233_, _06993_, _02091_);
  and _24637_ (_02234_, _06059_, _06039_);
  or _24638_ (_02235_, _02234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _24639_ (_02236_, _02206_, _06065_);
  and _24640_ (_02237_, _02236_, _02235_);
  and _24641_ (_02238_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _24642_ (_02240_, _02238_, _02237_);
  and _24643_ (_02241_, _02240_, _06036_);
  and _24644_ (_02242_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _24645_ (_02243_, _02242_, _02241_);
  or _24646_ (_02244_, _02243_, _02233_);
  and _24647_ (_01292_, _02244_, _06071_);
  and _24648_ (_01299_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06071_);
  and _24649_ (_02245_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _24650_ (_01306_, _02245_, _08574_);
  nor _24651_ (_02246_, _07344_, _06861_);
  and _24652_ (_02247_, _06866_, _07344_);
  or _24653_ (_02248_, _02247_, _02246_);
  and _24654_ (_01317_, _02248_, _06071_);
  and _24655_ (_02249_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _24656_ (_02250_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _24657_ (_02251_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24658_ (_02252_, _06059_, _06037_);
  nor _24659_ (_02253_, _02252_, _06065_);
  and _24660_ (_02254_, _02253_, _02251_);
  or _24661_ (_02256_, _02254_, _02249_);
  and _24662_ (_02257_, _02256_, _06036_);
  nor _24663_ (_02258_, _09037_, _02091_);
  and _24664_ (_02259_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _24665_ (_02260_, _02259_, _02258_);
  or _24666_ (_02262_, _02260_, _02257_);
  and _24667_ (_01328_, _02262_, _06071_);
  nand _24668_ (_02263_, _07945_, _06029_);
  and _24669_ (_02264_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _24670_ (_02265_, _06059_, _06038_);
  or _24671_ (_02266_, _02265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _24672_ (_02267_, _02234_, _06065_);
  and _24673_ (_02268_, _02267_, _02266_);
  or _24674_ (_02269_, _02268_, _02264_);
  or _24675_ (_02270_, _02269_, _06029_);
  and _24676_ (_02271_, _02270_, _02263_);
  or _24677_ (_02272_, _02271_, _02193_);
  not _24678_ (_02273_, _02193_);
  or _24679_ (_02275_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _24680_ (_02276_, _02275_, _06071_);
  and _24681_ (_01348_, _02276_, _02272_);
  nand _24682_ (_02277_, _06434_, _06029_);
  and _24683_ (_02278_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _24684_ (_02279_, _02252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _24685_ (_02280_, _02265_, _06065_);
  and _24686_ (_02281_, _02280_, _02279_);
  or _24687_ (_02282_, _02281_, _02278_);
  or _24688_ (_02283_, _02282_, _06029_);
  and _24689_ (_02284_, _02283_, _02277_);
  or _24690_ (_02285_, _02284_, _02193_);
  or _24691_ (_02286_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _24692_ (_02287_, _02286_, _06071_);
  and _24693_ (_01359_, _02287_, _02285_);
  or _24694_ (_02288_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _24695_ (_02289_, _06547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _24696_ (_02290_, _02289_, _02250_);
  and _24697_ (_02291_, _02290_, _02288_);
  or _24698_ (_02292_, _02291_, _06065_);
  not _24699_ (_02293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _24700_ (_02294_, _06065_, _02293_);
  and _24701_ (_02295_, _02294_, _02292_);
  and _24702_ (_02296_, _02295_, _06036_);
  and _24703_ (_02297_, _07978_, _06029_);
  and _24704_ (_02298_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _24705_ (_02299_, _02298_, _02297_);
  or _24706_ (_02300_, _02299_, _02296_);
  and _24707_ (_01367_, _02300_, _06071_);
  and _24708_ (_02301_, _00437_, _08993_);
  nor _24709_ (_02302_, _02301_, _07890_);
  and _24710_ (_02303_, _07901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _24711_ (_02304_, _02303_, _02302_);
  and _24712_ (_02305_, _02304_, _07913_);
  nand _24713_ (_02306_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _24714_ (_02307_, _02306_, _06560_);
  or _24715_ (_01408_, _02307_, _02305_);
  nand _24716_ (_02308_, _09341_, _07946_);
  or _24717_ (_02309_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _24718_ (_02310_, _02309_, _06071_);
  and _24719_ (_01442_, _02310_, _02308_);
  nor _24720_ (_01461_, _07874_, rst);
  and _24721_ (_02311_, _00761_, _05969_);
  nand _24722_ (_02312_, _02311_, _09341_);
  and _24723_ (_02313_, _06545_, _06062_);
  not _24724_ (_02314_, _02313_);
  and _24725_ (_02315_, _01062_, _05969_);
  nor _24726_ (_02316_, _02315_, _02314_);
  not _24727_ (_02317_, _02316_);
  and _24728_ (_02318_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _24729_ (_02319_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _24730_ (_02320_, _02319_, _02318_);
  or _24731_ (_02321_, _02311_, _02320_);
  and _24732_ (_02322_, _02321_, _06071_);
  and _24733_ (_01464_, _02322_, _02312_);
  and _24734_ (_02323_, _07105_, _06033_);
  or _24735_ (_02324_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _24736_ (_02325_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _24737_ (_02326_, _02325_, _02324_);
  or _24738_ (_02327_, _02326_, _02323_);
  nand _24739_ (_02328_, _02311_, _09037_);
  and _24740_ (_02329_, _02328_, _06071_);
  and _24741_ (_01501_, _02329_, _02327_);
  nand _24742_ (_02330_, _02311_, _06609_);
  nor _24743_ (_02331_, _02316_, _02101_);
  and _24744_ (_02332_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _24745_ (_02333_, _02332_, _02331_);
  or _24746_ (_02334_, _02333_, _02311_);
  and _24747_ (_02335_, _02334_, _06071_);
  and _24748_ (_01505_, _02335_, _02330_);
  nand _24749_ (_02336_, _02311_, _06993_);
  and _24750_ (_02337_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _24751_ (_02338_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _24752_ (_02339_, _02338_, _02337_);
  or _24753_ (_02340_, _02339_, _02311_);
  and _24754_ (_02341_, _02340_, _06071_);
  and _24755_ (_01512_, _02341_, _02336_);
  and _24756_ (_02342_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _24757_ (_02343_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _24758_ (_02344_, _02343_, _02342_);
  or _24759_ (_02345_, _02344_, _02311_);
  nand _24760_ (_02346_, _02311_, _07945_);
  and _24761_ (_02347_, _02346_, _06071_);
  and _24762_ (_01515_, _02347_, _02345_);
  and _24763_ (_02348_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _24764_ (_02349_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _24765_ (_02350_, _02349_, _02348_);
  or _24766_ (_02351_, _02350_, _02311_);
  nand _24767_ (_02352_, _02311_, _06434_);
  and _24768_ (_02353_, _02352_, _06071_);
  and _24769_ (_01517_, _02353_, _02351_);
  or _24770_ (_02354_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _24771_ (_02355_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _24772_ (_02356_, _02355_, _02354_);
  or _24773_ (_02357_, _02356_, _02323_);
  nand _24774_ (_02358_, _02311_, _07977_);
  and _24775_ (_02359_, _02358_, _06071_);
  and _24776_ (_01520_, _02359_, _02357_);
  not _24777_ (_02360_, _02315_);
  nor _24778_ (_02361_, _02360_, _09341_);
  nor _24779_ (_02362_, _02313_, _02226_);
  and _24780_ (_02363_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _24781_ (_02364_, _02363_, _02362_);
  nor _24782_ (_02365_, _02364_, _02315_);
  or _24783_ (_02366_, _02365_, _02323_);
  or _24784_ (_02367_, _02366_, _02361_);
  nand _24785_ (_02368_, _02323_, _02226_);
  and _24786_ (_02369_, _02368_, _06071_);
  and _24787_ (_01572_, _02369_, _02367_);
  nand _24788_ (_02370_, _02315_, _06609_);
  not _24789_ (_02371_, _02311_);
  and _24790_ (_02372_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _24791_ (_02373_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _24792_ (_02374_, _02373_, _02372_);
  or _24793_ (_02375_, _02374_, _02315_);
  and _24794_ (_02376_, _02375_, _02371_);
  and _24795_ (_02377_, _02376_, _02370_);
  and _24796_ (_02378_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _24797_ (_02379_, _02378_, _02377_);
  and _24798_ (_01575_, _02379_, _06071_);
  nand _24799_ (_02380_, _02315_, _06993_);
  and _24800_ (_02381_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _24801_ (_02382_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _24802_ (_02383_, _02382_, _02381_);
  or _24803_ (_02384_, _02383_, _02315_);
  and _24804_ (_02385_, _02384_, _02371_);
  and _24805_ (_02386_, _02385_, _02380_);
  and _24806_ (_02387_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _24807_ (_02388_, _02387_, _02386_);
  and _24808_ (_01580_, _02388_, _06071_);
  nand _24809_ (_02389_, _02315_, _07945_);
  and _24810_ (_02390_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _24811_ (_02391_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _24812_ (_02392_, _02391_, _02390_);
  or _24813_ (_02393_, _02392_, _02315_);
  and _24814_ (_02394_, _02393_, _02371_);
  and _24815_ (_02395_, _02394_, _02389_);
  and _24816_ (_02396_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _24817_ (_02397_, _02396_, _02395_);
  and _24818_ (_01616_, _02397_, _06071_);
  nand _24819_ (_02399_, _02315_, _06434_);
  and _24820_ (_02401_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _24821_ (_02402_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _24822_ (_02403_, _02402_, _02401_);
  or _24823_ (_02404_, _02403_, _02315_);
  and _24824_ (_02405_, _02404_, _02371_);
  and _24825_ (_02406_, _02405_, _02399_);
  and _24826_ (_02407_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _24827_ (_02408_, _02407_, _02406_);
  and _24828_ (_01618_, _02408_, _06071_);
  nand _24829_ (_02409_, _02315_, _09037_);
  or _24830_ (_02410_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _24831_ (_02411_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _24832_ (_02412_, _02411_, _02410_);
  or _24833_ (_02413_, _02412_, _02315_);
  and _24834_ (_02414_, _02413_, _02371_);
  and _24835_ (_02415_, _02414_, _02409_);
  and _24836_ (_02416_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _24837_ (_02417_, _02416_, _02415_);
  and _24838_ (_01620_, _02417_, _06071_);
  nor _24839_ (_02418_, _02313_, _02293_);
  and _24840_ (_02419_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _24841_ (_02420_, _02419_, _02418_);
  or _24842_ (_02421_, _02420_, _02315_);
  nand _24843_ (_02422_, _02315_, _07977_);
  and _24844_ (_02423_, _02422_, _02421_);
  or _24845_ (_02424_, _02423_, _02323_);
  nand _24846_ (_02425_, _02311_, _02293_);
  and _24847_ (_02426_, _02425_, _06071_);
  and _24848_ (_01624_, _02426_, _02424_);
  and _24849_ (_02428_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _24850_ (_02429_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _24851_ (_02430_, pc_log_change, _02429_);
  or _24852_ (_02431_, _02430_, _02428_);
  and _24853_ (_01642_, _02431_, _06071_);
  and _24854_ (_02432_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _24855_ (_02433_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _24856_ (_02434_, pc_log_change, _02433_);
  or _24857_ (_02435_, _02434_, _02432_);
  and _24858_ (_01648_, _02435_, _06071_);
  and _24859_ (_02436_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not _24860_ (_02437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor _24861_ (_02438_, pc_log_change, _02437_);
  or _24862_ (_02439_, _02438_, _02436_);
  and _24863_ (_01651_, _02439_, _06071_);
  and _24864_ (_02440_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _24865_ (_02441_, pc_log_change, _02076_);
  or _24866_ (_02442_, _02441_, _02440_);
  and _24867_ (_01658_, _02442_, _06071_);
  or _24868_ (_02443_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _24869_ (_02444_, pc_log_change, _06210_);
  and _24870_ (_02445_, _02444_, _06071_);
  and _24871_ (_01663_, _02445_, _02443_);
  and _24872_ (_02446_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _24873_ (_02447_, pc_log_change, _01876_);
  or _24874_ (_02448_, _02447_, _02446_);
  and _24875_ (_01673_, _02448_, _06071_);
  and _24876_ (_02449_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _24877_ (_02450_, pc_log_change, _02173_);
  or _24878_ (_02451_, _02450_, _02449_);
  and _24879_ (_01679_, _02451_, _06071_);
  and _24880_ (_01705_, t2_i, _06071_);
  and _24881_ (_02452_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _24882_ (_02453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _24883_ (_02454_, pc_log_change, _02453_);
  or _24884_ (_02455_, _02454_, _02452_);
  and _24885_ (_01716_, _02455_, _06071_);
  and _24886_ (_02456_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _24887_ (_02457_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _24888_ (_02458_, pc_log_change, _02457_);
  or _24889_ (_02459_, _02458_, _02456_);
  and _24890_ (_01719_, _02459_, _06071_);
  and _24891_ (_02460_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _24892_ (_02461_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _24893_ (_02462_, pc_log_change, _02461_);
  or _24894_ (_02463_, _02462_, _02460_);
  and _24895_ (_01730_, _02463_, _06071_);
  or _24896_ (_02464_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand _24897_ (_02465_, pc_log_change, _01996_);
  and _24898_ (_02467_, _02465_, _06071_);
  and _24899_ (_01732_, _02467_, _02464_);
  or _24900_ (_02468_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand _24901_ (_02469_, pc_log_change, _02437_);
  and _24902_ (_02470_, _02469_, _06071_);
  and _24903_ (_01734_, _02470_, _02468_);
  and _24904_ (_02471_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not _24905_ (_02472_, pc_log_change);
  and _24906_ (_02473_, _02472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _24907_ (_02474_, _02473_, _02471_);
  and _24908_ (_01736_, _02474_, _06071_);
  nor _24909_ (_02475_, _06359_, _02091_);
  not _24910_ (_02476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand _24911_ (_02477_, _06065_, _02476_);
  and _24912_ (_02478_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _24913_ (_02479_, _02478_, _06547_);
  not _24914_ (_02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _24915_ (_02481_, _02220_, _02480_);
  nor _24916_ (_02482_, _02481_, _02184_);
  or _24917_ (_02483_, _02482_, _06065_);
  or _24918_ (_02484_, _02483_, _02479_);
  and _24919_ (_02485_, _02484_, _02477_);
  and _24920_ (_02486_, _02485_, _06036_);
  and _24921_ (_02487_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _24922_ (_02488_, _02487_, _02486_);
  or _24923_ (_02489_, _02488_, _02475_);
  and _24924_ (_01739_, _02489_, _06071_);
  and _24925_ (_02491_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _24926_ (_02492_, _02472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _24927_ (_02493_, _02492_, _02491_);
  and _24928_ (_01743_, _02493_, _06071_);
  and _24929_ (_01763_, _07515_, _06071_);
  or _24930_ (_02494_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _24931_ (_02495_, _06530_, _05754_);
  and _24932_ (_02496_, _02495_, _06071_);
  and _24933_ (_01816_, _02496_, _02494_);
  nor _24934_ (_01829_, _11549_, rst);
  and _24935_ (_02497_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _24936_ (_02498_, _09341_, _06400_);
  and _24937_ (_02500_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and _24938_ (_02501_, _02500_, _09345_);
  or _24939_ (_02502_, _02501_, _02498_);
  or _24940_ (_02503_, _02502_, _02497_);
  and _24941_ (_01835_, _02503_, _06071_);
  and _24942_ (_01851_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and _24943_ (_02504_, _09583_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _24944_ (_02505_, _09003_, _09579_);
  and _24945_ (_02507_, _02505_, _09005_);
  or _24946_ (_02508_, _02507_, _02504_);
  and _24947_ (_01870_, _02508_, _06071_);
  and _24948_ (_02509_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _24949_ (_02510_, _11023_, _07979_);
  and _24950_ (_02511_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _24951_ (_02512_, _02511_, _07983_);
  or _24952_ (_02513_, _02512_, _02510_);
  or _24953_ (_02514_, _02513_, _02509_);
  and _24954_ (_01902_, _02514_, _06071_);
  and _24955_ (_02515_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _24956_ (_02516_, _08865_, _06993_);
  or _24957_ (_02517_, _02516_, _02515_);
  and _24958_ (_01914_, _02517_, _06071_);
  nor _24959_ (_02518_, _07011_, rst);
  or _24960_ (_02519_, _06528_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _24961_ (_04199_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06071_);
  and _24962_ (_02520_, _04199_, _02519_);
  or _24963_ (_02025_, _02520_, _02518_);
  and _24964_ (_02521_, _09576_, _06375_);
  nand _24965_ (_02522_, _06375_, _06011_);
  and _24966_ (_02523_, _02522_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _24967_ (_02524_, _02523_, _02521_);
  and _24968_ (_02041_, _02524_, _06071_);
  nor _24969_ (_02525_, _07945_, _06996_);
  and _24970_ (_02526_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _24971_ (_02527_, _02526_, _06390_);
  or _24972_ (_02528_, _02527_, _02525_);
  or _24973_ (_02529_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _24974_ (_02530_, _02529_, _06071_);
  and _24975_ (_02074_, _02530_, _02528_);
  and _24976_ (_02531_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _24977_ (_02532_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _24978_ (_02533_, _02532_, _02531_);
  and _24979_ (_02080_, _02533_, _06071_);
  nand _24980_ (_02534_, _11791_, _07759_);
  or _24981_ (_02535_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _24982_ (_02536_, _02535_, _06071_);
  and _24983_ (_02094_, _02536_, _02534_);
  or _24984_ (_02538_, _07757_, _07425_);
  or _24985_ (_02539_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _24986_ (_02540_, _02539_, _06071_);
  and _24987_ (_02099_, _02540_, _02538_);
  nor _24988_ (_02541_, _11791_, _07107_);
  and _24989_ (_02542_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _24990_ (_02543_, _02542_, _07429_);
  or _24991_ (_02544_, _02543_, _02541_);
  nand _24992_ (_02546_, _12466_, _07429_);
  and _24993_ (_02548_, _02546_, _06071_);
  and _24994_ (_02104_, _02548_, _02544_);
  and _24995_ (_02274_, _10978_, _06071_);
  and _24996_ (_03772_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06071_);
  and _24997_ (_02550_, _03772_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _24998_ (_02149_, _02550_, _02274_);
  and _24999_ (_02552_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _25000_ (_02553_, _08865_, _06359_);
  or _25001_ (_02554_, _02553_, _02552_);
  and _25002_ (_02175_, _02554_, _06071_);
  and _25003_ (_02556_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _25004_ (_02197_, _02556_, _08597_);
  nor _25005_ (_02239_, _11671_, rst);
  nand _25006_ (_02557_, _07946_, _06993_);
  or _25007_ (_02558_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _25008_ (_02560_, _02558_, _06071_);
  and _25009_ (_02255_, _02560_, _02557_);
  not _25010_ (_02562_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _25011_ (_02563_, _02562_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _25012_ (_02261_, _02563_, _06071_);
  and _25013_ (_02564_, _13711_, _06032_);
  or _25014_ (_02565_, _02564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _25015_ (_02566_, _02565_, _00557_);
  nand _25016_ (_02567_, _02564_, _06803_);
  and _25017_ (_02568_, _02567_, _02566_);
  nor _25018_ (_02569_, _00557_, _06609_);
  or _25019_ (_02570_, _02569_, _02568_);
  and _25020_ (_02398_, _02570_, _06071_);
  and _25021_ (_02571_, _13711_, _08801_);
  and _25022_ (_02572_, _02571_, _06803_);
  nor _25023_ (_02573_, _02571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _25024_ (_02574_, _02573_, _02572_);
  nand _25025_ (_02575_, _02574_, _00557_);
  nand _25026_ (_02576_, _13718_, _09341_);
  and _25027_ (_02577_, _02576_, _06071_);
  and _25028_ (_02400_, _02577_, _02575_);
  nand _25029_ (_02578_, _11825_, _06071_);
  nor _25030_ (_02427_, _02578_, _11933_);
  and _25031_ (_02579_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _25032_ (_02466_, _02579_, _08588_);
  and _25033_ (_02490_, _07848_, _06071_);
  and _25034_ (_02580_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _25035_ (_02581_, _09576_, _06385_);
  or _25036_ (_02582_, _02581_, _02580_);
  and _25037_ (_02499_, _02582_, _06071_);
  and _25038_ (_02506_, _07003_, _06508_);
  and _25039_ (_02537_, _00268_, _06071_);
  nor _25040_ (_02583_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _25041_ (_02584_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _25042_ (_02585_, _02584_, _02583_);
  nand _25043_ (_02586_, _02585_, _00472_);
  nand _25044_ (_02587_, _02586_, _06086_);
  or _25045_ (_02588_, _02586_, _06086_);
  and _25046_ (_02589_, _02588_, _02587_);
  and _25047_ (_02590_, _02589_, _11751_);
  and _25048_ (_02591_, _11827_, _07819_);
  and _25049_ (_02592_, _11748_, _07870_);
  nor _25050_ (_02593_, _00482_, _06086_);
  and _25051_ (_02594_, _00482_, _06086_);
  or _25052_ (_02595_, _02594_, _02593_);
  and _25053_ (_02596_, _02595_, _12469_);
  and _25054_ (_02597_, _12080_, _11424_);
  or _25055_ (_02598_, _02597_, _02596_);
  and _25056_ (_02599_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _25057_ (_02600_, _02599_, _02598_);
  nor _25058_ (_02601_, _02600_, _02592_);
  nand _25059_ (_02602_, _02601_, _12437_);
  or _25060_ (_02603_, _02602_, _02591_);
  or _25061_ (_02604_, _02603_, _02590_);
  and _25062_ (_02605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _25063_ (_02606_, _02605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _25064_ (_02607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _25065_ (_02608_, _02607_, _12502_);
  and _25066_ (_02609_, _02608_, _02606_);
  and _25067_ (_02610_, _02609_, _12500_);
  or _25068_ (_02611_, _02610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _25069_ (_02612_, _02610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _25070_ (_02613_, _02612_, _02611_);
  or _25071_ (_02614_, _02613_, _12437_);
  and _25072_ (_02615_, _02614_, _06071_);
  and _25073_ (_02545_, _02615_, _02604_);
  and _25074_ (_02616_, _05764_, _05722_);
  and _25075_ (_02617_, _02616_, _05875_);
  nor _25076_ (_02618_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _25077_ (_02619_, _02618_, _08705_);
  and _25078_ (_02620_, _02619_, _05805_);
  and _25079_ (_02621_, _05786_, _05743_);
  and _25080_ (_02622_, _02621_, _02620_);
  and _25081_ (_02623_, _05843_, _05825_);
  and _25082_ (_02624_, _02623_, _02622_);
  and _25083_ (_02547_, _02624_, _02617_);
  and _25084_ (_02625_, _10959_, _06006_);
  or _25085_ (_02626_, _02625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25086_ (_02627_, _02626_, _09250_);
  nand _25087_ (_02628_, _02625_, _06803_);
  and _25088_ (_02629_, _02628_, _02627_);
  nor _25089_ (_02630_, _09250_, _06993_);
  or _25090_ (_02631_, _02630_, _02629_);
  and _25091_ (_02549_, _02631_, _06071_);
  and _25092_ (_02632_, _01609_, _06362_);
  or _25093_ (_02633_, _02632_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _25094_ (_02634_, _02633_, _01623_);
  nand _25095_ (_02635_, _02632_, _06803_);
  and _25096_ (_02636_, _02635_, _02634_);
  nor _25097_ (_02637_, _01623_, _09037_);
  or _25098_ (_02638_, _02637_, _02636_);
  and _25099_ (_02551_, _02638_, _06071_);
  and _25100_ (_02639_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _25101_ (_02555_, _02639_, _07989_);
  and _25102_ (_02640_, _10972_, rxd_i);
  not _25103_ (_02641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor _25104_ (_02642_, _10972_, _02641_);
  or _25105_ (_02643_, _02642_, _02640_);
  and _25106_ (_02559_, _02643_, _06071_);
  or _25107_ (_02644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _25108_ (_02645_, _02644_, _01891_);
  not _25109_ (_02646_, _06805_);
  nor _25110_ (_02647_, _02646_, _06803_);
  nand _25111_ (_02648_, _02646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _25112_ (_02649_, _02648_, _01891_);
  or _25113_ (_02650_, _02649_, _02647_);
  and _25114_ (_02651_, _02650_, _02645_);
  or _25115_ (_02652_, _02651_, _01898_);
  nand _25116_ (_02653_, _01898_, _06359_);
  and _25117_ (_02654_, _02653_, _06071_);
  and _25118_ (_02561_, _02654_, _02652_);
  nand _25119_ (_02655_, _13723_, _06359_);
  or _25120_ (_02656_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _25121_ (_02657_, _02656_, _06071_);
  and _25122_ (_02665_, _02657_, _02655_);
  and _25123_ (_02658_, _13782_, _13731_);
  and _25124_ (_02659_, _13784_, _13736_);
  and _25125_ (_02660_, _02659_, _13780_);
  and _25126_ (_02661_, _02660_, _13777_);
  nand _25127_ (_02662_, _02661_, _13732_);
  nand _25128_ (_02663_, _02662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _25129_ (_02664_, _02663_, _02658_);
  or _25130_ (_02666_, _02664_, _13744_);
  and _25131_ (_02673_, _02666_, _06071_);
  and _25132_ (_02667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25133_ (_02668_, _07875_, _01916_);
  or _25134_ (_02669_, _02668_, _07879_);
  nor _25135_ (_02670_, _02669_, _02667_);
  or _25136_ (_02671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _25137_ (_02672_, _02671_, _06071_);
  nor _25138_ (_02674_, _02672_, _02670_);
  nor _25139_ (_02688_, _11453_, rst);
  nor _25140_ (_02675_, _13736_, _00436_);
  or _25141_ (_02676_, _02675_, _02661_);
  and _25142_ (_02677_, _02676_, _13733_);
  nand _25143_ (_02678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _25144_ (_02679_, _02678_, _13732_);
  or _25145_ (_02680_, _02679_, _02677_);
  and _25146_ (_02681_, _02680_, _13765_);
  or _25147_ (_02682_, _02681_, _02658_);
  and _25148_ (_02707_, _02682_, _13798_);
  or _25149_ (_02683_, _01691_, _01632_);
  and _25150_ (_02684_, _02683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _25151_ (_02685_, _02684_, _10952_);
  and _25152_ (_02686_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _25153_ (_02687_, _02686_, _00275_);
  and _25154_ (_02689_, _02687_, _10948_);
  or _25155_ (_02690_, _02689_, _02685_);
  nand _25156_ (_02691_, _10952_, _06434_);
  and _25157_ (_02692_, _02691_, _06071_);
  and _25158_ (_02737_, _02692_, _02690_);
  and _25159_ (_02693_, _01609_, _06383_);
  or _25160_ (_02694_, _02693_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _25161_ (_02695_, _02694_, _01623_);
  nand _25162_ (_02696_, _02693_, _06803_);
  and _25163_ (_02697_, _02696_, _02695_);
  and _25164_ (_02698_, _01608_, _07978_);
  or _25165_ (_02699_, _02698_, _02697_);
  and _25166_ (_02741_, _02699_, _06071_);
  and _25167_ (_02700_, _01609_, _06032_);
  or _25168_ (_02701_, _02700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _25169_ (_02702_, _02701_, _01623_);
  nand _25170_ (_02703_, _02700_, _06803_);
  and _25171_ (_02704_, _02703_, _02702_);
  nor _25172_ (_02705_, _01623_, _06609_);
  or _25173_ (_02706_, _02705_, _02704_);
  and _25174_ (_02752_, _02706_, _06071_);
  nor _25175_ (_02708_, _07912_, _07951_);
  or _25176_ (_02709_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _25177_ (_02710_, _02709_, _07896_);
  or _25178_ (_02711_, _02710_, _07887_);
  and _25179_ (_02712_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _25180_ (_02713_, _02712_, rxd_i);
  and _25181_ (_02714_, _02713_, _02711_);
  or _25182_ (_02715_, _02714_, _02708_);
  nand _25183_ (_02716_, _07887_, _09002_);
  and _25184_ (_02717_, _02716_, _06560_);
  and _25185_ (_02718_, _02717_, _02715_);
  and _25186_ (_02719_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _25187_ (_02754_, _02719_, _02718_);
  and _25188_ (_02720_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _25189_ (_02765_, _02720_, _07950_);
  nor _25190_ (_02721_, _02670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _25191_ (_02722_, _02721_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _25192_ (_02723_, _02721_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _25193_ (_02724_, _02723_, _06071_);
  and _25194_ (_02769_, _02724_, _02722_);
  and _25195_ (_02725_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _25196_ (_02726_, _02725_, _13798_);
  and _25197_ (_02727_, _13752_, _06071_);
  and _25198_ (_02728_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _25199_ (_02780_, _02728_, _02726_);
  nand _25200_ (_02729_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or _25201_ (_02730_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _25202_ (_02731_, _02730_, _02729_);
  and _25203_ (_02782_, _02731_, _13798_);
  and _25204_ (_02732_, _13711_, _06805_);
  or _25205_ (_02733_, _02732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _25206_ (_02734_, _02733_, _00557_);
  nand _25207_ (_02735_, _02732_, _06803_);
  and _25208_ (_02736_, _02735_, _02734_);
  nor _25209_ (_02738_, _00557_, _06359_);
  or _25210_ (_02739_, _02738_, _02736_);
  and _25211_ (_02786_, _02739_, _06071_);
  and _25212_ (_02740_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _25213_ (_02742_, _06530_, _05789_);
  or _25214_ (_02743_, _02742_, _02740_);
  and _25215_ (_02792_, _02743_, _06071_);
  nor _25216_ (_02744_, _06496_, _06490_);
  or _25217_ (_02745_, _06494_, _06483_);
  and _25218_ (_02746_, _06481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _25219_ (_02747_, _02746_, _02745_);
  and _25220_ (_02748_, _02747_, _02744_);
  and _25221_ (_02749_, _02748_, _01192_);
  or _25222_ (_02750_, _06470_, _06457_);
  and _25223_ (_02751_, _06468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _25224_ (_02753_, _02751_, _02750_);
  and _25225_ (_02755_, _02753_, _01176_);
  and _25226_ (_02756_, _02755_, _01482_);
  or _25227_ (_02757_, _02756_, _06508_);
  or _25228_ (_02758_, _02757_, _02749_);
  or _25229_ (_02759_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _25230_ (_02760_, _02759_, _06071_);
  and _25231_ (_02794_, _02760_, _02758_);
  nand _25232_ (_02761_, _01192_, _06511_);
  and _25233_ (_02762_, _06511_, _06474_);
  or _25234_ (_02763_, _02762_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _25235_ (_02764_, _02763_, _06071_);
  and _25236_ (_02810_, _02764_, _02761_);
  nand _25237_ (_02766_, _00727_, _01192_);
  and _25238_ (_02767_, _00727_, _06474_);
  or _25239_ (_02768_, _02767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _25240_ (_02770_, _02768_, _06071_);
  and _25241_ (_02813_, _02770_, _02766_);
  and _25242_ (_02771_, _10959_, _07754_);
  or _25243_ (_02772_, _02771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _25244_ (_02773_, _02772_, _09250_);
  nand _25245_ (_02774_, _02771_, _06803_);
  and _25246_ (_02775_, _02774_, _02773_);
  nor _25247_ (_02776_, _09250_, _06434_);
  or _25248_ (_02777_, _02776_, _02775_);
  and _25249_ (_02825_, _02777_, _06071_);
  and _25250_ (_02778_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _25251_ (_02779_, _06530_, _05773_);
  or _25252_ (_02781_, _02779_, _02778_);
  and _25253_ (_02874_, _02781_, _06071_);
  and _25254_ (_02783_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _25255_ (_02784_, _06530_, _05835_);
  or _25256_ (_02785_, _02784_, _02783_);
  and _25257_ (_02895_, _02785_, _06071_);
  and _25258_ (_02787_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _25259_ (_02788_, _06530_, _05817_);
  or _25260_ (_02789_, _02788_, _02787_);
  and _25261_ (_02908_, _02789_, _06071_);
  nor _25262_ (_02980_, _11904_, rst);
  or _25263_ (_02983_, _08776_, _08770_);
  and _25264_ (_03013_, _08032_, _06071_);
  nor _25265_ (_02790_, _13733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _25266_ (_02791_, _02790_, _13792_);
  and _25267_ (_03057_, _02791_, _13798_);
  and _25268_ (_02793_, _10943_, _06833_);
  and _25269_ (_02795_, _02793_, _06032_);
  nand _25270_ (_02796_, _02795_, _06803_);
  or _25271_ (_02797_, _02795_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25272_ (_02798_, _02797_, _06815_);
  and _25273_ (_02799_, _02798_, _02796_);
  and _25274_ (_02800_, _10951_, _06372_);
  not _25275_ (_02801_, _02800_);
  nor _25276_ (_02802_, _02801_, _06609_);
  not _25277_ (_02803_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor _25278_ (_02804_, _02800_, _02803_);
  or _25279_ (_02805_, _02804_, _02802_);
  and _25280_ (_02806_, _02805_, _06012_);
  nor _25281_ (_02807_, _06814_, _02803_);
  or _25282_ (_02808_, _02807_, rst);
  or _25283_ (_02809_, _02808_, _02806_);
  or _25284_ (_03119_, _02809_, _02799_);
  and _25285_ (_02811_, _06810_, _08801_);
  nand _25286_ (_02812_, _02811_, _06803_);
  or _25287_ (_02814_, _02811_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25288_ (_02815_, _02814_, _06815_);
  and _25289_ (_02816_, _02815_, _02812_);
  nand _25290_ (_02817_, _09341_, _06822_);
  or _25291_ (_02818_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25292_ (_02819_, _02818_, _06012_);
  and _25293_ (_02820_, _02819_, _02817_);
  not _25294_ (_02821_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor _25295_ (_02822_, _06814_, _02821_);
  or _25296_ (_02823_, _02822_, rst);
  or _25297_ (_02824_, _02823_, _02820_);
  or _25298_ (_03122_, _02824_, _02816_);
  and _25299_ (_02826_, _06810_, _06362_);
  nand _25300_ (_02827_, _02826_, _06803_);
  or _25301_ (_02828_, _02826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25302_ (_02829_, _02828_, _06815_);
  and _25303_ (_02830_, _02829_, _02827_);
  nand _25304_ (_02831_, _09037_, _06822_);
  or _25305_ (_02832_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25306_ (_02833_, _02832_, _06012_);
  and _25307_ (_02834_, _02833_, _02831_);
  and _25308_ (_02835_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _25309_ (_02836_, _02835_, rst);
  or _25310_ (_02837_, _02836_, _02834_);
  or _25311_ (_03124_, _02837_, _02830_);
  not _25312_ (_02838_, _06834_);
  or _25313_ (_02839_, _02838_, _01632_);
  and _25314_ (_02840_, _02839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25315_ (_02841_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25316_ (_02842_, _02841_, _00275_);
  and _25317_ (_02843_, _02842_, _06834_);
  or _25318_ (_02844_, _02843_, _02840_);
  and _25319_ (_02845_, _02844_, _06815_);
  nand _25320_ (_02846_, _06841_, _06434_);
  or _25321_ (_02847_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25322_ (_02848_, _02847_, _06012_);
  and _25323_ (_02849_, _02848_, _02846_);
  and _25324_ (_02850_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25325_ (_02851_, _02850_, rst);
  or _25326_ (_02852_, _02851_, _02849_);
  or _25327_ (_03127_, _02852_, _02845_);
  nor _25328_ (_03136_, _11469_, rst);
  and _25329_ (_02853_, _10943_, _06809_);
  and _25330_ (_02854_, _02853_, _06006_);
  nand _25331_ (_02855_, _02854_, _06803_);
  or _25332_ (_02856_, _02854_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25333_ (_02857_, _02856_, _06815_);
  and _25334_ (_02858_, _02857_, _02855_);
  and _25335_ (_02859_, _01607_, _06372_);
  not _25336_ (_02860_, _02859_);
  nor _25337_ (_02861_, _02860_, _06993_);
  not _25338_ (_02862_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor _25339_ (_02863_, _02859_, _02862_);
  or _25340_ (_02864_, _02863_, _02861_);
  and _25341_ (_02865_, _02864_, _06012_);
  nor _25342_ (_02866_, _06814_, _02862_);
  or _25343_ (_02867_, _02866_, rst);
  or _25344_ (_02868_, _02867_, _02865_);
  or _25345_ (_03146_, _02868_, _02858_);
  and _25346_ (_02869_, _02793_, _06006_);
  nand _25347_ (_02870_, _02869_, _06803_);
  or _25348_ (_02871_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _25349_ (_02872_, _02871_, _06815_);
  and _25350_ (_02873_, _02872_, _02870_);
  nor _25351_ (_02875_, _02801_, _06993_);
  not _25352_ (_02876_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor _25353_ (_02877_, _02800_, _02876_);
  or _25354_ (_02878_, _02877_, _02875_);
  and _25355_ (_02879_, _02878_, _06012_);
  nor _25356_ (_02880_, _06814_, _02876_);
  or _25357_ (_02881_, _02880_, rst);
  or _25358_ (_02882_, _02881_, _02879_);
  or _25359_ (_03148_, _02882_, _02873_);
  and _25360_ (_02883_, _06810_, _06032_);
  nand _25361_ (_02884_, _02883_, _06803_);
  or _25362_ (_02885_, _02883_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25363_ (_02886_, _02885_, _06815_);
  and _25364_ (_02887_, _02886_, _02884_);
  nand _25365_ (_02888_, _06822_, _06609_);
  or _25366_ (_02889_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25367_ (_02890_, _02889_, _06012_);
  and _25368_ (_02891_, _02890_, _02888_);
  not _25369_ (_02892_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor _25370_ (_02893_, _06814_, _02892_);
  or _25371_ (_02894_, _02893_, rst);
  or _25372_ (_02896_, _02894_, _02891_);
  or _25373_ (_03151_, _02896_, _02887_);
  and _25374_ (_02897_, _06810_, _06383_);
  nand _25375_ (_02898_, _02897_, _06803_);
  or _25376_ (_02899_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _25377_ (_02900_, _02899_, _06815_);
  and _25378_ (_02901_, _02900_, _02898_);
  nand _25379_ (_02902_, _07977_, _06822_);
  and _25380_ (_02903_, _02902_, _06012_);
  and _25381_ (_02904_, _02903_, _02899_);
  nor _25382_ (_02905_, _06814_, _00227_);
  or _25383_ (_02906_, _02905_, rst);
  or _25384_ (_02907_, _02906_, _02904_);
  or _25385_ (_03153_, _02907_, _02901_);
  and _25386_ (_02909_, _06810_, _07105_);
  nand _25387_ (_02910_, _02909_, _06803_);
  or _25388_ (_02911_, _02909_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25389_ (_02912_, _02911_, _06815_);
  and _25390_ (_02913_, _02912_, _02910_);
  nand _25391_ (_02914_, _07945_, _06822_);
  or _25392_ (_02915_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25393_ (_02916_, _02915_, _06012_);
  and _25394_ (_02917_, _02916_, _02914_);
  nor _25395_ (_02918_, _06814_, _00003_);
  or _25396_ (_02919_, _02918_, rst);
  or _25397_ (_02920_, _02919_, _02917_);
  or _25398_ (_03155_, _02920_, _02913_);
  and _25399_ (_02921_, _06834_, _08801_);
  nand _25400_ (_02922_, _02921_, _06803_);
  or _25401_ (_02923_, _02921_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25402_ (_02924_, _02923_, _06815_);
  and _25403_ (_02925_, _02924_, _02922_);
  nand _25404_ (_02926_, _09341_, _06841_);
  or _25405_ (_02927_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25406_ (_02928_, _02927_, _06012_);
  and _25407_ (_02929_, _02928_, _02926_);
  not _25408_ (_02930_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor _25409_ (_02931_, _06814_, _02930_);
  or _25410_ (_02932_, _02931_, rst);
  or _25411_ (_02933_, _02932_, _02929_);
  or _25412_ (_03157_, _02933_, _02925_);
  and _25413_ (_02934_, _06840_, _06363_);
  nand _25414_ (_02935_, _02934_, _06803_);
  or _25415_ (_02936_, _02934_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25416_ (_02937_, _02936_, _06815_);
  and _25417_ (_02938_, _02937_, _02935_);
  nand _25418_ (_02939_, _09037_, _06841_);
  or _25419_ (_02940_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25420_ (_02941_, _02940_, _06012_);
  and _25421_ (_02942_, _02941_, _02939_);
  and _25422_ (_02943_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _25423_ (_02944_, _02943_, rst);
  or _25424_ (_02945_, _02944_, _02942_);
  or _25425_ (_03159_, _02945_, _02938_);
  and _25426_ (_02946_, _06834_, _06006_);
  nand _25427_ (_02947_, _02946_, _06803_);
  or _25428_ (_02948_, _02946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25429_ (_02949_, _02948_, _06815_);
  and _25430_ (_02950_, _02949_, _02947_);
  nand _25431_ (_02951_, _06993_, _06841_);
  or _25432_ (_02952_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25433_ (_02953_, _02952_, _06012_);
  and _25434_ (_02954_, _02953_, _02951_);
  not _25435_ (_02955_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor _25436_ (_02956_, _06814_, _02955_);
  or _25437_ (_02957_, _02956_, rst);
  or _25438_ (_02958_, _02957_, _02954_);
  or _25439_ (_03162_, _02958_, _02950_);
  and _25440_ (_02959_, _02793_, _07105_);
  nand _25441_ (_02960_, _02959_, _06803_);
  or _25442_ (_02961_, _02959_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _25443_ (_02962_, _02961_, _06815_);
  and _25444_ (_02963_, _02962_, _02960_);
  nor _25445_ (_02964_, _02801_, _07945_);
  nor _25446_ (_02965_, _02800_, _13994_);
  or _25447_ (_02966_, _02965_, _02964_);
  and _25448_ (_02967_, _02966_, _06012_);
  nor _25449_ (_02968_, _06814_, _13994_);
  or _25450_ (_02969_, _02968_, rst);
  or _25451_ (_02970_, _02969_, _02967_);
  or _25452_ (_03245_, _02970_, _02963_);
  and _25453_ (_02971_, _02793_, _07754_);
  nand _25454_ (_02972_, _02971_, _06803_);
  or _25455_ (_02973_, _02971_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25456_ (_02974_, _02973_, _06815_);
  and _25457_ (_02975_, _02974_, _02972_);
  nor _25458_ (_02976_, _02801_, _06434_);
  and _25459_ (_02977_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25460_ (_02978_, _02977_, _02976_);
  and _25461_ (_02979_, _02978_, _06012_);
  and _25462_ (_02981_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25463_ (_02982_, _02981_, rst);
  or _25464_ (_02984_, _02982_, _02979_);
  or _25465_ (_03246_, _02984_, _02975_);
  and _25466_ (_02985_, _02793_, _06362_);
  nand _25467_ (_02986_, _02985_, _06803_);
  or _25468_ (_02987_, _02985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _25469_ (_02988_, _02987_, _06815_);
  and _25470_ (_02989_, _02988_, _02986_);
  nor _25471_ (_02990_, _02801_, _09037_);
  and _25472_ (_02991_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _25473_ (_02992_, _02991_, _02990_);
  and _25474_ (_02993_, _02992_, _06012_);
  and _25475_ (_02994_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _25476_ (_02995_, _02994_, rst);
  or _25477_ (_02996_, _02995_, _02993_);
  or _25478_ (_03261_, _02996_, _02989_);
  and _25479_ (_02997_, _02853_, _07754_);
  nand _25480_ (_02998_, _02997_, _06803_);
  or _25481_ (_02999_, _02997_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25482_ (_03000_, _02999_, _06815_);
  and _25483_ (_03001_, _03000_, _02998_);
  nor _25484_ (_03002_, _02860_, _06434_);
  and _25485_ (_03003_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25486_ (_03004_, _03003_, _03002_);
  and _25487_ (_03005_, _03004_, _06012_);
  and _25488_ (_03006_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _25489_ (_03007_, _03006_, rst);
  or _25490_ (_03008_, _03007_, _03005_);
  or _25491_ (_03263_, _03008_, _03001_);
  and _25492_ (_03009_, _02853_, _06362_);
  nand _25493_ (_03010_, _03009_, _06803_);
  or _25494_ (_03011_, _03009_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _25495_ (_03012_, _03011_, _06815_);
  and _25496_ (_03014_, _03012_, _03010_);
  nor _25497_ (_03015_, _02860_, _09037_);
  and _25498_ (_03016_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25499_ (_03017_, _03016_, _03015_);
  and _25500_ (_03018_, _03017_, _06012_);
  and _25501_ (_03019_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25502_ (_03020_, _03019_, rst);
  or _25503_ (_03021_, _03020_, _03018_);
  or _25504_ (_03264_, _03021_, _03014_);
  and _25505_ (_03022_, _02853_, _08801_);
  nand _25506_ (_03023_, _03022_, _06803_);
  or _25507_ (_03024_, _03022_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25508_ (_03025_, _03024_, _06815_);
  and _25509_ (_03026_, _03025_, _03023_);
  nor _25510_ (_03027_, _02860_, _09341_);
  not _25511_ (_03028_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor _25512_ (_03029_, _02859_, _03028_);
  or _25513_ (_03030_, _03029_, _03027_);
  and _25514_ (_03031_, _03030_, _06012_);
  nor _25515_ (_03032_, _06814_, _03028_);
  or _25516_ (_03033_, _03032_, rst);
  or _25517_ (_03034_, _03033_, _03031_);
  or _25518_ (_03270_, _03034_, _03026_);
  and _25519_ (_03035_, _06834_, _06383_);
  nand _25520_ (_03036_, _03035_, _06803_);
  or _25521_ (_03037_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _25522_ (_03038_, _03037_, _06815_);
  and _25523_ (_03039_, _03038_, _03036_);
  nand _25524_ (_03040_, _07977_, _06841_);
  and _25525_ (_03041_, _03037_, _06012_);
  and _25526_ (_03042_, _03041_, _03040_);
  nor _25527_ (_03043_, _06814_, _00222_);
  or _25528_ (_03044_, _03043_, rst);
  or _25529_ (_03045_, _03044_, _03042_);
  or _25530_ (_03285_, _03045_, _03039_);
  and _25531_ (_03046_, _06834_, _06032_);
  nand _25532_ (_03047_, _03046_, _06803_);
  or _25533_ (_03048_, _03046_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25534_ (_03049_, _03048_, _06815_);
  and _25535_ (_03050_, _03049_, _03047_);
  nand _25536_ (_03051_, _06841_, _06609_);
  or _25537_ (_03052_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25538_ (_03053_, _03052_, _06012_);
  and _25539_ (_03054_, _03053_, _03051_);
  not _25540_ (_03055_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor _25541_ (_03056_, _06814_, _03055_);
  or _25542_ (_03058_, _03056_, rst);
  or _25543_ (_03059_, _03058_, _03054_);
  or _25544_ (_03287_, _03059_, _03050_);
  and _25545_ (_03060_, _06834_, _07105_);
  nand _25546_ (_03061_, _03060_, _06803_);
  or _25547_ (_03062_, _03060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25548_ (_03063_, _03062_, _06815_);
  and _25549_ (_03064_, _03063_, _03061_);
  nand _25550_ (_03065_, _07945_, _06841_);
  or _25551_ (_03066_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25552_ (_03067_, _03066_, _06012_);
  and _25553_ (_03068_, _03067_, _03065_);
  nor _25554_ (_03069_, _06814_, _14003_);
  or _25555_ (_03070_, _03069_, rst);
  or _25556_ (_03071_, _03070_, _03068_);
  or _25557_ (_03289_, _03071_, _03064_);
  and _25558_ (_03072_, _02793_, _06383_);
  nand _25559_ (_03073_, _03072_, _06803_);
  or _25560_ (_03074_, _03072_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _25561_ (_03075_, _03074_, _06815_);
  and _25562_ (_03076_, _03075_, _03073_);
  and _25563_ (_03077_, _02800_, _07978_);
  nor _25564_ (_03078_, _02800_, _00211_);
  or _25565_ (_03079_, _03078_, _03077_);
  and _25566_ (_03080_, _03079_, _06012_);
  nor _25567_ (_03081_, _06814_, _00211_);
  or _25568_ (_03082_, _03081_, rst);
  or _25569_ (_03083_, _03082_, _03080_);
  or _25570_ (_03291_, _03083_, _03076_);
  and _25571_ (_03084_, _06810_, _06006_);
  nand _25572_ (_03085_, _03084_, _06803_);
  or _25573_ (_03086_, _03084_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25574_ (_03087_, _03086_, _06815_);
  and _25575_ (_03088_, _03087_, _03085_);
  nand _25576_ (_03089_, _06993_, _06822_);
  or _25577_ (_03090_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25578_ (_03091_, _03090_, _06012_);
  and _25579_ (_03092_, _03091_, _03089_);
  not _25580_ (_03093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor _25581_ (_03094_, _06814_, _03093_);
  or _25582_ (_03095_, _03094_, rst);
  or _25583_ (_03096_, _03095_, _03092_);
  or _25584_ (_03294_, _03096_, _03088_);
  and _25585_ (_03097_, _06810_, _07754_);
  nand _25586_ (_03098_, _03097_, _06803_);
  or _25587_ (_03099_, _03097_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25588_ (_03100_, _03099_, _06815_);
  and _25589_ (_03101_, _03100_, _03098_);
  nand _25590_ (_03102_, _06822_, _06434_);
  or _25591_ (_03103_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25592_ (_03104_, _03103_, _06012_);
  and _25593_ (_03105_, _03104_, _03102_);
  and _25594_ (_03106_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _25595_ (_03107_, _03106_, rst);
  or _25596_ (_03108_, _03107_, _03105_);
  or _25597_ (_03296_, _03108_, _03101_);
  nand _25598_ (_03109_, _02859_, _06803_);
  or _25599_ (_03110_, _02859_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _25600_ (_03111_, _03110_, _06815_);
  and _25601_ (_03112_, _03111_, _03109_);
  nand _25602_ (_03113_, _02859_, _07977_);
  and _25603_ (_03114_, _03113_, _06012_);
  and _25604_ (_03115_, _03114_, _03110_);
  nor _25605_ (_03116_, _06814_, _00216_);
  or _25606_ (_03117_, _03116_, rst);
  or _25607_ (_03118_, _03117_, _03115_);
  or _25608_ (_03298_, _03118_, _03112_);
  and _25609_ (_03120_, _02793_, _08801_);
  nand _25610_ (_03121_, _03120_, _06803_);
  or _25611_ (_03123_, _03120_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25612_ (_03125_, _03123_, _06815_);
  and _25613_ (_03126_, _03125_, _03121_);
  nor _25614_ (_03128_, _02801_, _09341_);
  not _25615_ (_03129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor _25616_ (_03130_, _02800_, _03129_);
  or _25617_ (_03131_, _03130_, _03128_);
  and _25618_ (_03132_, _03131_, _06012_);
  nor _25619_ (_03133_, _06814_, _03129_);
  or _25620_ (_03134_, _03133_, rst);
  or _25621_ (_03135_, _03134_, _03132_);
  or _25622_ (_03300_, _03135_, _03126_);
  and _25623_ (_03137_, _02853_, _06032_);
  nand _25624_ (_03138_, _03137_, _06803_);
  or _25625_ (_03139_, _03137_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25626_ (_03140_, _03139_, _06815_);
  and _25627_ (_03141_, _03140_, _03138_);
  nor _25628_ (_03142_, _02860_, _06609_);
  not _25629_ (_03143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor _25630_ (_03144_, _02859_, _03143_);
  or _25631_ (_03145_, _03144_, _03142_);
  and _25632_ (_03147_, _03145_, _06012_);
  nor _25633_ (_03149_, _06814_, _03143_);
  or _25634_ (_03150_, _03149_, rst);
  or _25635_ (_03152_, _03150_, _03147_);
  or _25636_ (_03303_, _03152_, _03141_);
  and _25637_ (_03154_, _02853_, _07105_);
  nand _25638_ (_03156_, _03154_, _06803_);
  or _25639_ (_03158_, _03154_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _25640_ (_03160_, _03158_, _06815_);
  and _25641_ (_03161_, _03160_, _03156_);
  nor _25642_ (_03163_, _02860_, _07945_);
  nor _25643_ (_03164_, _02859_, _13986_);
  or _25644_ (_03165_, _03164_, _03163_);
  and _25645_ (_03166_, _03165_, _06012_);
  nor _25646_ (_03167_, _06814_, _13986_);
  or _25647_ (_03168_, _03167_, rst);
  or _25648_ (_03169_, _03168_, _03166_);
  or _25649_ (_03305_, _03169_, _03161_);
  nor _25650_ (_03170_, _09037_, _06996_);
  and _25651_ (_03171_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or _25652_ (_03172_, _03171_, _06390_);
  or _25653_ (_03173_, _03172_, _03170_);
  or _25654_ (_03174_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _25655_ (_03175_, _03174_, _06071_);
  and _25656_ (_03317_, _03175_, _03173_);
  or _25657_ (_03176_, _08065_, _08032_);
  nor _25658_ (_03177_, _03176_, _07103_);
  nand _25659_ (_03178_, _03177_, _07751_);
  or _25660_ (_03179_, _03178_, _07609_);
  or _25661_ (_03180_, _03179_, _07365_);
  and _25662_ (_03181_, _03180_, _07344_);
  or _25663_ (_03182_, _06712_, _06710_);
  not _25664_ (_03183_, _06618_);
  nand _25665_ (_03184_, _06710_, _03183_);
  and _25666_ (_03185_, _03184_, _06615_);
  and _25667_ (_03186_, _03185_, _03182_);
  nand _25668_ (_03187_, _06747_, _06717_);
  and _25669_ (_03188_, _06748_, _06715_);
  and _25670_ (_03189_, _03188_, _03187_);
  and _25671_ (_03190_, _07454_, _07109_);
  and _25672_ (_03191_, _03190_, _07449_);
  nand _25673_ (_03192_, _03191_, _07108_);
  nand _25674_ (_03193_, _03192_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _25675_ (_03194_, _03193_, _03189_);
  nor _25676_ (_03195_, _03194_, _03186_);
  and _25677_ (_03196_, _03195_, _07684_);
  nand _25678_ (_03197_, _03196_, _07788_);
  or _25679_ (_03198_, _03197_, _03181_);
  nor _25680_ (_03199_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _25681_ (_03200_, _03199_, _10896_);
  and _25682_ (_03201_, _03200_, _03198_);
  and _25683_ (_03202_, _00274_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _25684_ (_03203_, _03202_, _00275_);
  nand _25685_ (_03204_, _03203_, _10896_);
  nand _25686_ (_03205_, _03204_, _08985_);
  or _25687_ (_03206_, _03205_, _03201_);
  nand _25688_ (_03207_, _08988_, _06434_);
  and _25689_ (_03208_, _03207_, _06071_);
  and _25690_ (_03322_, _03208_, _03206_);
  nand _25691_ (_03209_, _09037_, _07946_);
  or _25692_ (_03210_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _25693_ (_03211_, _03210_, _06071_);
  and _25694_ (_03330_, _03211_, _03209_);
  nor _25695_ (_03212_, _06967_, _06359_);
  and _25696_ (_03213_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _25697_ (_03214_, _03213_, _03212_);
  and _25698_ (_03344_, _03214_, _06071_);
  and _25699_ (_03347_, _08065_, _06071_);
  and _25700_ (_03215_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _25701_ (_03216_, _06530_, _05739_);
  or _25702_ (_03217_, _03216_, _03215_);
  and _25703_ (_03351_, _03217_, _06071_);
  and _25704_ (_03218_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _25705_ (_03219_, _06530_, _05716_);
  or _25706_ (_03220_, _03219_, _03218_);
  and _25707_ (_03353_, _03220_, _06071_);
  or _25708_ (_03221_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _25709_ (_03222_, _06530_, _05798_);
  and _25710_ (_03223_, _03222_, _06071_);
  and _25711_ (_03356_, _03223_, _03221_);
  and _25712_ (_03224_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _25713_ (_03225_, _06530_, _05782_);
  or _25714_ (_03226_, _03225_, _03224_);
  and _25715_ (_03358_, _03226_, _06071_);
  nor _25716_ (_03227_, _09341_, _06996_);
  and _25717_ (_03228_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _25718_ (_03229_, _03228_, _06390_);
  or _25719_ (_03230_, _03229_, _03227_);
  or _25720_ (_03231_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _25721_ (_03232_, _03231_, _06071_);
  and _25722_ (_03377_, _03232_, _03230_);
  and _25723_ (_03233_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _25724_ (_03234_, _06530_, _05749_);
  or _25725_ (_03235_, _03234_, _03233_);
  and _25726_ (_03424_, _03235_, _06071_);
  or _25727_ (_03236_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _25728_ (_03237_, _06530_, _05865_);
  and _25729_ (_03238_, _03237_, _06071_);
  and _25730_ (_03431_, _03238_, _03236_);
  and _25731_ (_03239_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _25732_ (_03240_, _06530_, _05737_);
  or _25733_ (_03241_, _03240_, _03239_);
  and _25734_ (_03440_, _03241_, _06071_);
  or _25735_ (_03242_, _09583_, _07893_);
  or _25736_ (_03243_, _09005_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _25737_ (_03244_, _03243_, _06071_);
  and _25738_ (_03444_, _03244_, _03242_);
  and _25739_ (_03450_, _07741_, _06071_);
  and _25740_ (_03247_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _25741_ (_03248_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _25742_ (_03249_, _03248_, _03247_);
  and _25743_ (_03472_, _03249_, _06071_);
  and _25744_ (_03250_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _25745_ (_03251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _25746_ (_03252_, _11290_, _03251_);
  and _25747_ (_03253_, _11290_, _03251_);
  nor _25748_ (_03254_, _03253_, _03252_);
  and _25749_ (_03255_, _03254_, _11297_);
  nor _25750_ (_03256_, _03254_, _11297_);
  or _25751_ (_03257_, _03256_, _03255_);
  or _25752_ (_03258_, _03257_, _09711_);
  or _25753_ (_03259_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _25754_ (_03260_, _03259_, _11270_);
  and _25755_ (_03262_, _03260_, _03258_);
  or _25756_ (_03479_, _03262_, _03250_);
  nor _25757_ (_03481_, _12052_, rst);
  nor _25758_ (_03265_, _06530_, _06528_);
  nor _25759_ (_03266_, _11370_, _11367_);
  nor _25760_ (_03267_, _03266_, _06528_);
  and _25761_ (_03268_, _03267_, _05694_);
  nor _25762_ (_03269_, _03267_, _05694_);
  nor _25763_ (_03271_, _03269_, _03268_);
  nor _25764_ (_03272_, _03271_, _03265_);
  and _25765_ (_03273_, _05699_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _25766_ (_03274_, _03273_, _03265_);
  nor _25767_ (_03275_, _03274_, _11234_);
  or _25768_ (_03276_, _03275_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _25769_ (_03277_, _03276_, _03272_);
  and _25770_ (_03485_, _03277_, _06071_);
  or _25771_ (_03278_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _25772_ (_03279_, _06530_, _05835_);
  and _25773_ (_03280_, _03279_, _06071_);
  and _25774_ (_03488_, _03280_, _03278_);
  and _25775_ (_03499_, _07604_, _06071_);
  and _25776_ (_03500_, _07680_, _06071_);
  nor _25777_ (_03521_, _11763_, rst);
  or _25778_ (_03281_, _01784_, _07564_);
  not _25779_ (_03282_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _25780_ (_03283_, _01784_, _03282_);
  and _25781_ (_03284_, _03283_, _06012_);
  and _25782_ (_03286_, _03284_, _03281_);
  nor _25783_ (_03288_, _06814_, _03282_);
  or _25784_ (_03290_, _01791_, _01632_);
  and _25785_ (_03292_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _25786_ (_03293_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _25787_ (_03295_, _03293_, _00275_);
  and _25788_ (_03297_, _03295_, _01783_);
  or _25789_ (_03299_, _03297_, _03292_);
  and _25790_ (_03301_, _03299_, _06815_);
  or _25791_ (_03302_, _03301_, _03288_);
  or _25792_ (_03304_, _03302_, _03286_);
  and _25793_ (_03554_, _03304_, _06071_);
  and _25794_ (_03306_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _25795_ (_03307_, _06530_, _10690_);
  or _25796_ (_03308_, _03307_, _03306_);
  and _25797_ (_03563_, _03308_, _06071_);
  or _25798_ (_03309_, _08535_, _05747_);
  or _25799_ (_03310_, _06526_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _25800_ (_03311_, _03310_, _06071_);
  and _25801_ (_03565_, _03311_, _03309_);
  and _25802_ (_03312_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _25803_ (_03313_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nand _25804_ (_03314_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _25805_ (_03315_, _03314_, _03313_);
  nand _25806_ (_03316_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand _25807_ (_03318_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _25808_ (_03319_, _03318_, _03316_);
  and _25809_ (_03320_, _03319_, _03315_);
  nand _25810_ (_03321_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand _25811_ (_03323_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _25812_ (_03324_, _03323_, _03321_);
  nand _25813_ (_03325_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand _25814_ (_03326_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _25815_ (_03327_, _03326_, _03325_);
  and _25816_ (_03328_, _03327_, _03324_);
  and _25817_ (_03329_, _03328_, _03320_);
  nand _25818_ (_03331_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand _25819_ (_03332_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _25820_ (_03333_, _03332_, _03331_);
  nand _25821_ (_03334_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand _25822_ (_03335_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _25823_ (_03336_, _03335_, _03334_);
  and _25824_ (_03337_, _03336_, _03333_);
  nand _25825_ (_03338_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nand _25826_ (_03339_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and _25827_ (_03340_, _03339_, _03338_);
  nand _25828_ (_03341_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _25829_ (_03342_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _25830_ (_03343_, _03342_, _03341_);
  and _25831_ (_03345_, _03343_, _03340_);
  and _25832_ (_03346_, _03345_, _03337_);
  and _25833_ (_03348_, _03346_, _03329_);
  nand _25834_ (_03349_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _25835_ (_03350_, _13897_, _12143_);
  and _25836_ (_03352_, _03350_, _03349_);
  nand _25837_ (_03354_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _25838_ (_03355_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _25839_ (_03357_, _03355_, _03354_);
  and _25840_ (_03359_, _03357_, _03352_);
  nor _25841_ (_03360_, _13983_, p1_in[5]);
  and _25842_ (_03361_, _13983_, _02892_);
  nor _25843_ (_03362_, _03361_, _03360_);
  nand _25844_ (_03363_, _03362_, _14007_);
  nor _25845_ (_03364_, _13983_, p0_in[5]);
  and _25846_ (_03365_, _13983_, _03055_);
  nor _25847_ (_03366_, _03365_, _03364_);
  nand _25848_ (_03367_, _03366_, _14000_);
  and _25849_ (_03368_, _03367_, _03363_);
  nor _25850_ (_03369_, _13983_, p3_in[5]);
  and _25851_ (_03370_, _13983_, _03143_);
  nor _25852_ (_03371_, _03370_, _03369_);
  nand _25853_ (_03372_, _03371_, _13966_);
  nor _25854_ (_03373_, _13983_, p2_in[5]);
  and _25855_ (_03374_, _13983_, _02803_);
  nor _25856_ (_03375_, _03374_, _03373_);
  nand _25857_ (_03376_, _03375_, _13991_);
  and _25858_ (_03378_, _03376_, _03372_);
  and _25859_ (_03379_, _03378_, _03368_);
  and _25860_ (_03380_, _03379_, _03359_);
  nand _25861_ (_03381_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _25862_ (_03382_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _25863_ (_03383_, _03382_, _03381_);
  and _25864_ (_03384_, _03383_, _03380_);
  nand _25865_ (_03385_, _03384_, _03348_);
  nand _25866_ (_03386_, _03385_, _13919_);
  nand _25867_ (_03387_, _03386_, _13925_);
  or _25868_ (_03388_, _03387_, _03312_);
  nand _25869_ (_03389_, _13924_, _07643_);
  and _25870_ (_03390_, _03389_, _06071_);
  and _25871_ (_03570_, _03390_, _03388_);
  and _25872_ (_03391_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor _25873_ (_03392_, _06967_, _06434_);
  or _25874_ (_03393_, _03392_, _03391_);
  and _25875_ (_03576_, _03393_, _06071_);
  or _25876_ (_03394_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _25877_ (_03395_, _06530_, _05793_);
  and _25878_ (_03396_, _03395_, _06071_);
  and _25879_ (_03579_, _03396_, _03394_);
  and _25880_ (_03585_, _07536_, _06071_);
  or _25881_ (_03397_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _25882_ (_03398_, _06530_, _05732_);
  and _25883_ (_03399_, _03398_, _06071_);
  and _25884_ (_03587_, _03399_, _03397_);
  or _25885_ (_03400_, _01784_, _00366_);
  not _25886_ (_03401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _25887_ (_03402_, _01784_, _03401_);
  and _25888_ (_03403_, _03402_, _06012_);
  and _25889_ (_03404_, _03403_, _03400_);
  nor _25890_ (_03405_, _06814_, _03401_);
  and _25891_ (_03406_, _01783_, _06032_);
  nand _25892_ (_03407_, _03406_, _06803_);
  or _25893_ (_03408_, _03406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _25894_ (_03409_, _03408_, _06815_);
  and _25895_ (_03410_, _03409_, _03407_);
  or _25896_ (_03411_, _03410_, _03405_);
  or _25897_ (_03412_, _03411_, _03404_);
  and _25898_ (_03592_, _03412_, _06071_);
  and _25899_ (_03413_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _25900_ (_03414_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _25901_ (_03415_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _25902_ (_03416_, _03415_, _03414_);
  nand _25903_ (_03417_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand _25904_ (_03418_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _25905_ (_03419_, _03418_, _03417_);
  and _25906_ (_03420_, _03419_, _03416_);
  nand _25907_ (_03421_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand _25908_ (_03422_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _25909_ (_03423_, _03422_, _03421_);
  nand _25910_ (_03425_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand _25911_ (_03426_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _25912_ (_03427_, _03426_, _03425_);
  and _25913_ (_03428_, _03427_, _03423_);
  and _25914_ (_03429_, _03428_, _03420_);
  nand _25915_ (_03430_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand _25916_ (_03432_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _25917_ (_03433_, _03432_, _03430_);
  nand _25918_ (_03434_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand _25919_ (_03435_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _25920_ (_03436_, _03435_, _03434_);
  and _25921_ (_03437_, _03436_, _03433_);
  nand _25922_ (_03438_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _25923_ (_03439_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _25924_ (_03441_, _03439_, _03438_);
  nand _25925_ (_03442_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _25926_ (_03443_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _25927_ (_03445_, _03443_, _03442_);
  and _25928_ (_03446_, _03445_, _03441_);
  and _25929_ (_03447_, _03446_, _03437_);
  and _25930_ (_03448_, _03447_, _03429_);
  nand _25931_ (_03449_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _25932_ (_03451_, _13897_, _12100_);
  and _25933_ (_03452_, _03451_, _03449_);
  nand _25934_ (_03453_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand _25935_ (_03454_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _25936_ (_03455_, _03454_, _03453_);
  and _25937_ (_03456_, _03455_, _03452_);
  nor _25938_ (_03457_, _13983_, p2_in[6]);
  and _25939_ (_03458_, _13983_, _03129_);
  nor _25940_ (_03459_, _03458_, _03457_);
  nand _25941_ (_03460_, _03459_, _13991_);
  nor _25942_ (_03461_, _13983_, p3_in[6]);
  and _25943_ (_03462_, _13983_, _03028_);
  nor _25944_ (_03463_, _03462_, _03461_);
  nand _25945_ (_03464_, _03463_, _13966_);
  and _25946_ (_03465_, _03464_, _03460_);
  nor _25947_ (_03466_, _13983_, p0_in[6]);
  and _25948_ (_03467_, _13983_, _02930_);
  nor _25949_ (_03468_, _03467_, _03466_);
  nand _25950_ (_03469_, _03468_, _14000_);
  nor _25951_ (_03470_, _13983_, p1_in[6]);
  and _25952_ (_03471_, _13983_, _02821_);
  nor _25953_ (_03473_, _03471_, _03470_);
  nand _25954_ (_03474_, _03473_, _14007_);
  and _25955_ (_03475_, _03474_, _03469_);
  and _25956_ (_03476_, _03475_, _03465_);
  and _25957_ (_03477_, _03476_, _03456_);
  nand _25958_ (_03478_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _25959_ (_03480_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _25960_ (_03482_, _03480_, _03478_);
  and _25961_ (_03484_, _03482_, _03477_);
  nand _25962_ (_03486_, _03484_, _03448_);
  nand _25963_ (_03487_, _03486_, _13919_);
  nand _25964_ (_03489_, _03487_, _13925_);
  or _25965_ (_03490_, _03489_, _03413_);
  nand _25966_ (_03491_, _13924_, _07426_);
  and _25967_ (_03492_, _03491_, _06071_);
  and _25968_ (_03614_, _03492_, _03490_);
  and _25969_ (_03617_, _11935_, _06071_);
  or _25970_ (_03493_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _25971_ (_03494_, _06530_, _05708_);
  and _25972_ (_03495_, _03494_, _06071_);
  and _25973_ (_03630_, _03495_, _03493_);
  and _25974_ (_03639_, _08062_, _06071_);
  nor _25975_ (_03645_, _12163_, rst);
  or _25976_ (_03496_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _25977_ (_03497_, _06530_, _05791_);
  and _25978_ (_03498_, _03497_, _06071_);
  and _25979_ (_03650_, _03498_, _03496_);
  nor _25980_ (_03652_, _12199_, rst);
  nor _25981_ (_03669_, _12021_, rst);
  nand _25982_ (_03671_, _12336_, _06071_);
  nor _25983_ (_03678_, _12420_, rst);
  and _25984_ (_03501_, _12524_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _25985_ (_03502_, _01721_, _11865_);
  and _25986_ (_03503_, _11396_, _13379_);
  and _25987_ (_03504_, _11874_, _11408_);
  and _25988_ (_03505_, _11400_, _11396_);
  or _25989_ (_03506_, _03505_, _03504_);
  or _25990_ (_03507_, _03506_, _03503_);
  and _25991_ (_03508_, _11404_, _11396_);
  or _25992_ (_03509_, _03508_, _11859_);
  or _25993_ (_03510_, _03509_, _03507_);
  or _25994_ (_03511_, _03510_, _03502_);
  and _25995_ (_03512_, _13639_, _11422_);
  or _25996_ (_03513_, _03512_, _11837_);
  and _25997_ (_03514_, _13379_, _08732_);
  and _25998_ (_03515_, _03514_, _11412_);
  and _25999_ (_03516_, _03514_, _11810_);
  or _26000_ (_03517_, _03516_, _03515_);
  and _26001_ (_03518_, _11401_, _08757_);
  and _26002_ (_03519_, _11410_, _08757_);
  or _26003_ (_03520_, _03519_, _03518_);
  or _26004_ (_03522_, _03520_, _03517_);
  or _26005_ (_03523_, _03522_, _03513_);
  and _26006_ (_03524_, _11810_, _11410_);
  and _26007_ (_03525_, _11415_, _11401_);
  or _26008_ (_03526_, _03525_, _03524_);
  and _26009_ (_03527_, _11404_, _08732_);
  and _26010_ (_03528_, _03527_, _08757_);
  and _26011_ (_03529_, _11414_, _08757_);
  or _26012_ (_03530_, _03529_, _03528_);
  and _26013_ (_03531_, _03514_, _11422_);
  and _26014_ (_03532_, _11404_, _11391_);
  or _26015_ (_03533_, _03532_, _03531_);
  or _26016_ (_03534_, _03533_, _03530_);
  or _26017_ (_03535_, _03534_, _03526_);
  or _26018_ (_03536_, _11803_, _11413_);
  and _26019_ (_03537_, _13632_, _11391_);
  and _26020_ (_03538_, _11889_, _11408_);
  or _26021_ (_03539_, _03538_, _13352_);
  or _26022_ (_03540_, _03539_, _03537_);
  or _26023_ (_03541_, _03540_, _03536_);
  and _26024_ (_03542_, _11415_, _03527_);
  or _26025_ (_03543_, _03542_, _03541_);
  or _26026_ (_03544_, _03543_, _03535_);
  or _26027_ (_03545_, _03544_, _03523_);
  or _26028_ (_03546_, _03545_, _03511_);
  and _26029_ (_03547_, _03546_, _08775_);
  or _26030_ (_03682_, _03547_, _03501_);
  or _26031_ (_03548_, _08535_, _05726_);
  or _26032_ (_03549_, _06526_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _26033_ (_03550_, _03549_, _06071_);
  and _26034_ (_03702_, _03550_, _03548_);
  and _26035_ (_03551_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _26036_ (_03552_, _06530_, _06962_);
  or _26037_ (_03553_, _03552_, _03551_);
  and _26038_ (_03713_, _03553_, _06071_);
  and _26039_ (_03555_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _26040_ (_03556_, _06530_, _06850_);
  or _26041_ (_03557_, _03556_, _03555_);
  and _26042_ (_03715_, _03557_, _06071_);
  and _26043_ (_03558_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _26044_ (_03725_, _03558_, _08603_);
  and _26045_ (_03559_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _26046_ (_03560_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand _26047_ (_03561_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _26048_ (_03562_, _03561_, _03560_);
  nand _26049_ (_03564_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _26050_ (_03566_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _26051_ (_03567_, _03566_, _03564_);
  and _26052_ (_03568_, _03567_, _03562_);
  nand _26053_ (_03569_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _26054_ (_03571_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _26055_ (_03572_, _03571_, _03569_);
  nand _26056_ (_03573_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _26057_ (_03574_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _26058_ (_03575_, _03574_, _03573_);
  and _26059_ (_03577_, _03575_, _03572_);
  and _26060_ (_03578_, _03577_, _03568_);
  nand _26061_ (_03580_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _26062_ (_03581_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _26063_ (_03582_, _03581_, _03580_);
  nand _26064_ (_03583_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand _26065_ (_03584_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _26066_ (_03586_, _03584_, _03583_);
  and _26067_ (_03588_, _03586_, _03582_);
  nand _26068_ (_03589_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand _26069_ (_03590_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _26070_ (_03591_, _03590_, _03589_);
  nand _26071_ (_03593_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _26072_ (_03594_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _26073_ (_03595_, _03594_, _03593_);
  and _26074_ (_03596_, _03595_, _03591_);
  and _26075_ (_03597_, _03596_, _03588_);
  and _26076_ (_03598_, _03597_, _03578_);
  nand _26077_ (_03599_, _13897_, _12213_);
  nand _26078_ (_03600_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _26079_ (_03601_, _03600_, _03599_);
  nand _26080_ (_03602_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _26081_ (_03603_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _26082_ (_03604_, _03603_, _03602_);
  and _26083_ (_03605_, _03604_, _03601_);
  nor _26084_ (_03606_, _13983_, p0_in[4]);
  and _26085_ (_03607_, _13983_, _02955_);
  nor _26086_ (_03608_, _03607_, _03606_);
  nand _26087_ (_03609_, _03608_, _14000_);
  nor _26088_ (_03610_, _13983_, p1_in[4]);
  and _26089_ (_03611_, _13983_, _03093_);
  nor _26090_ (_03612_, _03611_, _03610_);
  nand _26091_ (_03613_, _03612_, _14007_);
  and _26092_ (_03615_, _03613_, _03609_);
  nor _26093_ (_03616_, _13983_, p3_in[4]);
  and _26094_ (_03618_, _13983_, _02862_);
  nor _26095_ (_03619_, _03618_, _03616_);
  nand _26096_ (_03620_, _03619_, _13966_);
  nor _26097_ (_03621_, _13983_, p2_in[4]);
  and _26098_ (_03622_, _13983_, _02876_);
  nor _26099_ (_03623_, _03622_, _03621_);
  nand _26100_ (_03624_, _03623_, _13991_);
  and _26101_ (_03625_, _03624_, _03620_);
  and _26102_ (_03626_, _03625_, _03615_);
  and _26103_ (_03627_, _03626_, _03605_);
  nand _26104_ (_03628_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand _26105_ (_03629_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _26106_ (_03631_, _03629_, _03628_);
  and _26107_ (_03632_, _03631_, _03627_);
  nand _26108_ (_03633_, _03632_, _03598_);
  nand _26109_ (_03634_, _03633_, _13919_);
  nand _26110_ (_03635_, _03634_, _13925_);
  or _26111_ (_03636_, _03635_, _03559_);
  nand _26112_ (_03637_, _13924_, _07715_);
  and _26113_ (_03638_, _03637_, _06071_);
  and _26114_ (_03740_, _03638_, _03636_);
  or _26115_ (_03640_, _13975_, _13625_);
  or _26116_ (_03641_, _03640_, _01722_);
  not _26117_ (_03642_, _11861_);
  and _26118_ (_03643_, _08748_, _08732_);
  and _26119_ (_03644_, _03643_, _11412_);
  or _26120_ (_03646_, _03644_, _03642_);
  or _26121_ (_03647_, _11885_, _11413_);
  or _26122_ (_03648_, _11857_, _11847_);
  or _26123_ (_03649_, _03648_, _03647_);
  or _26124_ (_03651_, _03649_, _03646_);
  nand _26125_ (_03653_, _11842_, _11835_);
  or _26126_ (_03654_, _03653_, _03651_);
  or _26127_ (_03655_, _03654_, _03641_);
  and _26128_ (_03656_, _11889_, _08760_);
  or _26129_ (_03657_, _03656_, _11917_);
  or _26130_ (_03658_, _13627_, _11868_);
  or _26131_ (_03659_, _03658_, _03657_);
  or _26132_ (_03660_, _03659_, _03655_);
  and _26133_ (_03661_, _03660_, _06527_);
  and _26134_ (_03662_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26135_ (_03663_, _11403_, _11385_);
  or _26136_ (_03664_, _03663_, _13643_);
  or _26137_ (_03665_, _03664_, _03662_);
  or _26138_ (_03666_, _03665_, _03661_);
  and _26139_ (_03742_, _03666_, _06071_);
  and _26140_ (_03667_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _26141_ (_03668_, _06530_, _06532_);
  or _26142_ (_03670_, _03668_, _03667_);
  and _26143_ (_03748_, _03670_, _06071_);
  and _26144_ (_03672_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08003_);
  and _26145_ (_03673_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _26146_ (_03674_, _03673_, _03672_);
  and _26147_ (_03752_, _03674_, _06071_);
  or _26148_ (_03675_, _08535_, _05847_);
  or _26149_ (_03676_, _06526_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _26150_ (_03677_, _03676_, _06071_);
  and _26151_ (_03756_, _03677_, _03675_);
  nand _26152_ (_03679_, _02311_, _06359_);
  and _26153_ (_03680_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _26154_ (_03681_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _26155_ (_03683_, _03681_, _03680_);
  or _26156_ (_03684_, _03683_, _02311_);
  and _26157_ (_03685_, _03684_, _06071_);
  and _26158_ (_03780_, _03685_, _03679_);
  nand _26159_ (_03686_, _07946_, _06609_);
  or _26160_ (_03687_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _26161_ (_03688_, _03687_, _06071_);
  and _26162_ (_03813_, _03688_, _03686_);
  and _26163_ (_03689_, _12524_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and _26164_ (_03690_, _11840_, _08757_);
  or _26165_ (_03691_, _03529_, _03524_);
  or _26166_ (_03692_, _03691_, _03690_);
  and _26167_ (_03693_, _11396_, _11388_);
  and _26168_ (_03694_, _11391_, _11388_);
  or _26169_ (_03695_, _03694_, _03693_);
  or _26170_ (_03696_, _11876_, _03695_);
  or _26171_ (_03697_, _03696_, _01721_);
  or _26172_ (_03698_, _03697_, _03692_);
  and _26173_ (_03699_, _13967_, _11387_);
  or _26174_ (_03700_, _03699_, _11909_);
  or _26175_ (_03701_, _03700_, _13360_);
  or _26176_ (_03703_, _03701_, _13353_);
  or _26177_ (_03704_, _11856_, _12548_);
  or _26178_ (_03705_, _03528_, _03704_);
  or _26179_ (_03706_, _03705_, _03703_);
  or _26180_ (_03707_, _03706_, _03698_);
  or _26181_ (_03708_, _03707_, _03523_);
  and _26182_ (_03709_, _03708_, _08775_);
  or _26183_ (_03822_, _03709_, _03689_);
  and _26184_ (_03710_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _26185_ (_03711_, _07979_, _12197_);
  and _26186_ (_03712_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _26187_ (_03714_, _03712_, _07983_);
  or _26188_ (_03716_, _03714_, _03711_);
  or _26189_ (_03717_, _03716_, _03710_);
  and _26190_ (_03823_, _03717_, _06071_);
  and _26191_ (_03718_, _13346_, _08732_);
  and _26192_ (_03719_, _13360_, _08732_);
  or _26193_ (_03720_, _13337_, _11811_);
  or _26194_ (_03721_, _03720_, _08761_);
  or _26195_ (_03722_, _03721_, _03719_);
  and _26196_ (_03723_, _13360_, _08764_);
  or _26197_ (_03724_, _12542_, _11908_);
  or _26198_ (_03726_, _03724_, _13349_);
  or _26199_ (_03727_, _03726_, _03723_);
  or _26200_ (_03728_, _03727_, _03722_);
  or _26201_ (_03729_, _03728_, _03718_);
  not _26202_ (_03730_, _11836_);
  or _26203_ (_03731_, _12533_, _03730_);
  and _26204_ (_03732_, _11840_, _11415_);
  or _26205_ (_03733_, _03524_, _11844_);
  nor _26206_ (_03734_, _03733_, _03732_);
  nand _26207_ (_03735_, _03734_, _11804_);
  or _26208_ (_03736_, _11916_, _13978_);
  or _26209_ (_03737_, _03736_, _03735_);
  or _26210_ (_03738_, _03737_, _03731_);
  or _26211_ (_03739_, _03738_, _03729_);
  and _26212_ (_03741_, _03739_, _08775_);
  and _26213_ (_03743_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _26214_ (_03744_, _11811_, _11744_);
  or _26215_ (_03746_, _03744_, _03743_);
  and _26216_ (_03747_, _03746_, _06071_);
  or _26217_ (_03834_, _03747_, _03741_);
  and _26218_ (_03749_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _26219_ (_03750_, _07979_, _12019_);
  and _26220_ (_03751_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and _26221_ (_03753_, _03751_, _07983_);
  or _26222_ (_03754_, _03753_, _03750_);
  or _26223_ (_03755_, _03754_, _03749_);
  and _26224_ (_03837_, _03755_, _06071_);
  nand _26225_ (_03757_, _07946_, _06359_);
  or _26226_ (_03758_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _26227_ (_03759_, _03758_, _06071_);
  and _26228_ (_03847_, _03759_, _03757_);
  and _26229_ (_03760_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08003_);
  and _26230_ (_03761_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _26231_ (_03762_, _03761_, _03760_);
  and _26232_ (_03853_, _03762_, _06071_);
  and _26233_ (_03763_, _02793_, _06805_);
  nand _26234_ (_03764_, _03763_, _06803_);
  or _26235_ (_03765_, _03763_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _26236_ (_03766_, _03765_, _06815_);
  and _26237_ (_03767_, _03766_, _03764_);
  nor _26238_ (_03768_, _02801_, _06359_);
  and _26239_ (_03769_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _26240_ (_03770_, _03769_, _03768_);
  and _26241_ (_03771_, _03770_, _06012_);
  and _26242_ (_03773_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _26243_ (_03774_, _03773_, rst);
  or _26244_ (_03775_, _03774_, _03771_);
  or _26245_ (_03862_, _03775_, _03767_);
  and _26246_ (_03776_, _02853_, _06805_);
  nand _26247_ (_03777_, _03776_, _06803_);
  or _26248_ (_03778_, _03776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _26249_ (_03779_, _03778_, _06815_);
  and _26250_ (_03781_, _03779_, _03777_);
  nor _26251_ (_03782_, _02860_, _06359_);
  and _26252_ (_03783_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _26253_ (_03784_, _03783_, _03782_);
  and _26254_ (_03785_, _03784_, _06012_);
  and _26255_ (_03786_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _26256_ (_03787_, _03786_, rst);
  or _26257_ (_03788_, _03787_, _03785_);
  or _26258_ (_03867_, _03788_, _03781_);
  and _26259_ (_03880_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or _26260_ (_03789_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  nand _26261_ (_03790_, _06530_, _11005_);
  and _26262_ (_03791_, _03790_, _06071_);
  and _26263_ (_03889_, _03791_, _03789_);
  and _26264_ (_03891_, _00283_, _06071_);
  and _26265_ (_03792_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _26266_ (_03793_, _03792_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _26267_ (_03794_, _03792_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _26268_ (_03795_, _03794_, _03793_);
  and _26269_ (_03897_, _03795_, _06071_);
  or _26270_ (_03796_, _01784_, _07819_);
  not _26271_ (_03797_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _26272_ (_03798_, _01784_, _03797_);
  and _26273_ (_03799_, _03798_, _06012_);
  and _26274_ (_03800_, _03799_, _03796_);
  nor _26275_ (_03801_, _06814_, _03797_);
  and _26276_ (_03802_, _01783_, _06805_);
  nand _26277_ (_03803_, _03802_, _06803_);
  or _26278_ (_03804_, _03802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26279_ (_03805_, _03804_, _06815_);
  and _26280_ (_03806_, _03805_, _03803_);
  or _26281_ (_03807_, _03806_, _03801_);
  or _26282_ (_03808_, _03807_, _03800_);
  and _26283_ (_03903_, _03808_, _06071_);
  or _26284_ (_03809_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _26285_ (_03810_, _06530_, _05817_);
  and _26286_ (_03811_, _03810_, _06071_);
  and _26287_ (_03907_, _03811_, _03809_);
  nor _26288_ (_03812_, _02360_, _06359_);
  nor _26289_ (_03814_, _02313_, _02476_);
  and _26290_ (_03815_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor _26291_ (_03816_, _03815_, _03814_);
  nor _26292_ (_03817_, _03816_, _02315_);
  or _26293_ (_03818_, _03817_, _02323_);
  or _26294_ (_03819_, _03818_, _03812_);
  nand _26295_ (_03820_, _02323_, _02476_);
  and _26296_ (_03821_, _03820_, _06071_);
  and _26297_ (_03919_, _03821_, _03819_);
  nor _26298_ (_03824_, _06996_, _06359_);
  and _26299_ (_03825_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _26300_ (_03826_, _03825_, _06390_);
  or _26301_ (_03827_, _03826_, _03824_);
  or _26302_ (_03828_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _26303_ (_03829_, _03828_, _06071_);
  and _26304_ (_03924_, _03829_, _03827_);
  and _26305_ (_03929_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or _26306_ (_03830_, _08535_, _05829_);
  or _26307_ (_03831_, _06526_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _26308_ (_03832_, _03831_, _06071_);
  and _26309_ (_03936_, _03832_, _03830_);
  and _26310_ (_03833_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _26311_ (_03835_, _07979_, _12161_);
  and _26312_ (_03836_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and _26313_ (_03838_, _03836_, _07983_);
  or _26314_ (_03839_, _03838_, _03835_);
  or _26315_ (_03840_, _03839_, _03833_);
  and _26316_ (_03968_, _03840_, _06071_);
  or _26317_ (_03841_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _26318_ (_03842_, _06530_, _05789_);
  and _26319_ (_03843_, _03842_, _06071_);
  and _26320_ (_04006_, _03843_, _03841_);
  and _26321_ (_03844_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _26322_ (_03845_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _26323_ (_03846_, _03845_, _03844_);
  and _26324_ (_04040_, _03846_, _06071_);
  or _26325_ (_03848_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand _26326_ (_03849_, _06530_, _09701_);
  and _26327_ (_03850_, _03849_, _06071_);
  and _26328_ (_04050_, _03850_, _03848_);
  and _26329_ (_04054_, _00247_, _06071_);
  and _26330_ (_03851_, _11097_, _05860_);
  and _26331_ (_03852_, _11117_, _05849_);
  or _26332_ (_03854_, _03852_, _11202_);
  or _26333_ (_03855_, _03854_, _03851_);
  or _26334_ (_03856_, _11178_, _05851_);
  or _26335_ (_03857_, _03856_, _03855_);
  or _26336_ (_03858_, _03857_, _11125_);
  nand _26337_ (_03859_, _11138_, _11101_);
  nand _26338_ (_03860_, _11231_, _03859_);
  and _26339_ (_03861_, _11139_, _05850_);
  or _26340_ (_03863_, _11117_, _11171_);
  and _26341_ (_03864_, _03863_, _11101_);
  or _26342_ (_03865_, _03864_, _03861_);
  or _26343_ (_03866_, _03865_, _03860_);
  or _26344_ (_03868_, _03866_, _05885_);
  nand _26345_ (_03869_, _11136_, _11112_);
  or _26346_ (_03870_, _03869_, _03868_);
  or _26347_ (_03871_, _03870_, _03858_);
  and _26348_ (_03872_, _03871_, _08705_);
  nor _26349_ (_03873_, _05691_, _13383_);
  or _26350_ (_03874_, _03873_, rst);
  or _26351_ (_04056_, _03874_, _03872_);
  or _26352_ (_03875_, _13340_, _11845_);
  and _26353_ (_03876_, _11830_, _11391_);
  or _26354_ (_03877_, _03876_, _13976_);
  or _26355_ (_03878_, _03877_, _03875_);
  not _26356_ (_03879_, _11910_);
  or _26357_ (_03881_, _13344_, _03879_);
  or _26358_ (_03882_, _03881_, _03878_);
  and _26359_ (_03883_, _13354_, _11390_);
  or _26360_ (_03884_, _03883_, _03732_);
  or _26361_ (_03885_, _03884_, _12546_);
  or _26362_ (_03886_, _03885_, _03882_);
  and _26363_ (_03887_, _11884_, _11810_);
  or _26364_ (_03888_, _03647_, _03887_);
  or _26365_ (_03890_, _03888_, _03525_);
  or _26366_ (_03892_, _12549_, _11416_);
  or _26367_ (_03893_, _03892_, _03539_);
  and _26368_ (_03894_, _11830_, _11396_);
  and _26369_ (_03895_, _11414_, _08756_);
  or _26370_ (_03896_, _03895_, _13335_);
  or _26371_ (_03898_, _03896_, _03894_);
  nor _26372_ (_03899_, _03898_, _03893_);
  nand _26373_ (_03900_, _03899_, _13979_);
  or _26374_ (_03901_, _03900_, _03890_);
  or _26375_ (_03902_, _03901_, _03886_);
  and _26376_ (_03904_, _03902_, _06527_);
  and _26377_ (_03905_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26378_ (_03906_, _03905_, _11817_);
  or _26379_ (_03908_, _03906_, _03904_);
  and _26380_ (_04065_, _03908_, _06071_);
  nor _26381_ (_04070_, _11823_, rst);
  and _26382_ (_03909_, _11840_, _11810_);
  or _26383_ (_03910_, _13349_, _13340_);
  or _26384_ (_03911_, _03910_, _03909_);
  or _26385_ (_03912_, _03911_, _13346_);
  or _26386_ (_03913_, _12535_, _11868_);
  or _26387_ (_03914_, _03913_, _03644_);
  or _26388_ (_03915_, _11909_, _11811_);
  or _26389_ (_03916_, _03915_, _11738_);
  or _26390_ (_03917_, _03916_, _03914_);
  or _26391_ (_03918_, _13353_, _03894_);
  and _26392_ (_03920_, _11397_, _08749_);
  or _26393_ (_03921_, _03920_, _03918_);
  or _26394_ (_03922_, _03921_, _03917_);
  or _26395_ (_03923_, _13335_, _11812_);
  or _26396_ (_03925_, _03923_, _13355_);
  or _26397_ (_03926_, _03925_, _03892_);
  or _26398_ (_03927_, _11833_, _11806_);
  or _26399_ (_03928_, _11880_, _11853_);
  or _26400_ (_03930_, _03928_, _03927_);
  or _26401_ (_03931_, _03930_, _03926_);
  or _26402_ (_03932_, _03931_, _03922_);
  or _26403_ (_03933_, _03932_, _03912_);
  and _26404_ (_03934_, _03933_, _06527_);
  and _26405_ (_03935_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26406_ (_03937_, _13641_, _11744_);
  or _26407_ (_03938_, _13385_, _03937_);
  or _26408_ (_03939_, _03938_, _03935_);
  or _26409_ (_03940_, _03939_, _03934_);
  and _26410_ (_04077_, _03940_, _06071_);
  or _26411_ (_03941_, _13924_, rst);
  nor _26412_ (_04086_, _03941_, _13919_);
  and _26413_ (_04089_, _00427_, _06071_);
  or _26414_ (_03942_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  nand _26415_ (_03943_, _06530_, _10989_);
  and _26416_ (_03944_, _03943_, _06071_);
  and _26417_ (_04094_, _03944_, _03942_);
  nor _26418_ (_04107_, _00294_, rst);
  and _26419_ (_03945_, _11867_, _11422_);
  or _26420_ (_03946_, _03723_, _13629_);
  or _26421_ (_03947_, _03946_, _03945_);
  or _26422_ (_03948_, _03947_, _03722_);
  or _26423_ (_03949_, _03948_, _03926_);
  and _26424_ (_03950_, _11391_, _08748_);
  or _26425_ (_03951_, _03950_, _11909_);
  or _26426_ (_03952_, _03951_, _11738_);
  or _26427_ (_03953_, _13627_, _12533_);
  and _26428_ (_03954_, _11412_, _08750_);
  and _26429_ (_03955_, _11736_, _11810_);
  or _26430_ (_03956_, _03955_, _03954_);
  or _26431_ (_03957_, _03956_, _03953_);
  or _26432_ (_03958_, _03957_, _03952_);
  or _26433_ (_03959_, _03918_, _13625_);
  or _26434_ (_03960_, _03959_, _03958_);
  or _26435_ (_03961_, _03960_, _03912_);
  or _26436_ (_03962_, _03961_, _03949_);
  and _26437_ (_03963_, _03962_, _06527_);
  and _26438_ (_03964_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26439_ (_03965_, _03964_, _03938_);
  or _26440_ (_03966_, _03965_, _03963_);
  and _26441_ (_04111_, _03966_, _06071_);
  and _26442_ (_03967_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _26443_ (_03969_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _26444_ (_03970_, _03969_, _03967_);
  and _26445_ (_03971_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _26446_ (_03972_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _26447_ (_03973_, _03972_, _03971_);
  or _26448_ (_03974_, _03973_, _03970_);
  and _26449_ (_03975_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _26450_ (_03976_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _26451_ (_03977_, _03976_, _03975_);
  and _26452_ (_03978_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _26453_ (_03979_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _26454_ (_03980_, _03979_, _03978_);
  or _26455_ (_03981_, _03980_, _03977_);
  or _26456_ (_03982_, _03981_, _03974_);
  and _26457_ (_03983_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _26458_ (_03984_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _26459_ (_03985_, _03984_, _03983_);
  and _26460_ (_03986_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _26461_ (_03987_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _26462_ (_03988_, _03987_, _03986_);
  or _26463_ (_03989_, _03988_, _03985_);
  and _26464_ (_03990_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _26465_ (_03991_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _26466_ (_03992_, _03991_, _03990_);
  and _26467_ (_03993_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _26468_ (_03994_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _26469_ (_03995_, _03994_, _03993_);
  or _26470_ (_03996_, _03995_, _03992_);
  or _26471_ (_03997_, _03996_, _03989_);
  or _26472_ (_03998_, _03997_, _03982_);
  and _26473_ (_03999_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26474_ (_04000_, _13897_, _12076_);
  or _26475_ (_04001_, _04000_, _03999_);
  and _26476_ (_04002_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _26477_ (_04003_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _26478_ (_04004_, _04003_, _04002_);
  or _26479_ (_04005_, _04004_, _04001_);
  or _26480_ (_04007_, _13983_, p2_in[7]);
  or _26481_ (_04008_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _26482_ (_04009_, _04008_, _04007_);
  and _26483_ (_04010_, _04009_, _13991_);
  or _26484_ (_04011_, _13983_, p3_in[7]);
  or _26485_ (_04012_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _26486_ (_04013_, _04012_, _04011_);
  and _26487_ (_04014_, _04013_, _13966_);
  or _26488_ (_04015_, _04014_, _04010_);
  or _26489_ (_04016_, _13983_, p0_in[7]);
  or _26490_ (_04017_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _26491_ (_04018_, _04017_, _04016_);
  and _26492_ (_04019_, _04018_, _14000_);
  or _26493_ (_04020_, _13983_, p1_in[7]);
  or _26494_ (_04021_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _26495_ (_04022_, _04021_, _04020_);
  and _26496_ (_04023_, _04022_, _14007_);
  or _26497_ (_04024_, _04023_, _04019_);
  or _26498_ (_04025_, _04024_, _04015_);
  or _26499_ (_04026_, _04025_, _04005_);
  and _26500_ (_04027_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _26501_ (_04028_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _26502_ (_04029_, _04028_, _04027_);
  or _26503_ (_04030_, _04029_, _04026_);
  or _26504_ (_04031_, _04030_, _03998_);
  and _26505_ (_04032_, _04031_, _13919_);
  and _26506_ (_04033_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _26507_ (_04034_, _04033_, _04032_);
  or _26508_ (_04035_, _04034_, _13924_);
  or _26509_ (_04036_, _13925_, _07819_);
  and _26510_ (_04037_, _04036_, _06071_);
  and _26511_ (_04114_, _04037_, _04035_);
  not _26512_ (_04038_, _08774_);
  and _26513_ (_04039_, _04038_, _08771_);
  or _26514_ (_04041_, _08776_, _08761_);
  or _26515_ (_04122_, _04041_, _04039_);
  or _26516_ (_04042_, _08535_, _05768_);
  or _26517_ (_04043_, _06526_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _26518_ (_04044_, _04043_, _06071_);
  and _26519_ (_04144_, _04044_, _04042_);
  and _26520_ (_04045_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or _26521_ (_04046_, _12274_, _11735_);
  or _26522_ (_04047_, _04046_, _03690_);
  and _26523_ (_04048_, _11410_, _08756_);
  or _26524_ (_04049_, _04048_, _12549_);
  or _26525_ (_04051_, _04049_, _11841_);
  or _26526_ (_04052_, _04051_, _12269_);
  or _26527_ (_04053_, _04052_, _12532_);
  or _26528_ (_04055_, _04053_, _04047_);
  and _26529_ (_04057_, _04055_, _08775_);
  or _26530_ (_04146_, _04057_, _04045_);
  or _26531_ (_04058_, _03538_, _11908_);
  or _26532_ (_04059_, _04058_, _03732_);
  or _26533_ (_04060_, _12535_, _11803_);
  or _26534_ (_04061_, _04060_, _04059_);
  and _26535_ (_04062_, _04061_, _06527_);
  and _26536_ (_04063_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26537_ (_04064_, _04063_, _04062_);
  or _26538_ (_04066_, _04064_, _13642_);
  and _26539_ (_04154_, _04066_, _06071_);
  and _26540_ (_04067_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or _26541_ (_04068_, _03694_, _12548_);
  or _26542_ (_04069_, _04068_, _12547_);
  or _26543_ (_04071_, _03883_, _11912_);
  or _26544_ (_04072_, _04071_, _04069_);
  or _26545_ (_04073_, _04072_, _04060_);
  or _26546_ (_04074_, _04073_, _03890_);
  and _26547_ (_04075_, _04074_, _08775_);
  or _26548_ (_04157_, _04075_, _04067_);
  and _26549_ (_04076_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26550_ (_04078_, _13639_, _11412_);
  and _26551_ (_04079_, _04078_, _06527_);
  or _26552_ (_04080_, _04079_, _04076_);
  or _26553_ (_04081_, _04080_, _13642_);
  and _26554_ (_04159_, _04081_, _06071_);
  or _26555_ (_04083_, _13628_, _12532_);
  and _26556_ (_04084_, _04083_, _11421_);
  or _26557_ (_04085_, _04084_, _13385_);
  or _26558_ (_04087_, _13638_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26559_ (_04088_, _04087_, _04085_);
  or _26560_ (_04090_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05686_);
  and _26561_ (_04091_, _04090_, _06071_);
  and _26562_ (_04164_, _04091_, _04088_);
  and _26563_ (_04092_, _12524_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _26564_ (_04093_, _03538_, _11859_);
  or _26565_ (_04095_, _04093_, _03536_);
  or _26566_ (_04096_, _04048_, _03537_);
  or _26567_ (_04097_, _04096_, _03525_);
  or _26568_ (_04098_, _11876_, _11839_);
  or _26569_ (_04099_, _04098_, _03506_);
  or _26570_ (_04100_, _04099_, _04097_);
  or _26571_ (_04101_, _04100_, _04095_);
  and _26572_ (_04102_, _04101_, _08775_);
  or _26573_ (_04166_, _04102_, _04092_);
  and _26574_ (_04103_, _12524_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nor _26575_ (_04104_, _13332_, _11837_);
  nand _26576_ (_04105_, _04104_, _11846_);
  nor _26577_ (_04106_, _04105_, _12543_);
  nand _26578_ (_04108_, _04106_, _13977_);
  or _26579_ (_04109_, _04108_, _03890_);
  or _26580_ (_04110_, _13346_, _12528_);
  or _26581_ (_04112_, _04110_, _03884_);
  or _26582_ (_04113_, _04112_, _03731_);
  or _26583_ (_04115_, _04113_, _04109_);
  and _26584_ (_04116_, _04115_, _08775_);
  or _26585_ (_04168_, _04116_, _04103_);
  or _26586_ (_04117_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _26587_ (_04118_, _06530_, _05773_);
  and _26588_ (_04119_, _04118_, _06071_);
  and _26589_ (_04184_, _04119_, _04117_);
  and _26590_ (_04120_, _13884_, _12030_);
  or _26591_ (_04121_, _00303_, _13849_);
  or _26592_ (_04123_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _26593_ (_04124_, _04123_, _13818_);
  and _26594_ (_04125_, _04124_, _04121_);
  and _26595_ (_04126_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _26596_ (_04127_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _26597_ (_04128_, _04127_, _04126_);
  and _26598_ (_04129_, _04128_, _13849_);
  nor _26599_ (_04130_, _12426_, _10916_);
  and _26600_ (_04131_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _26601_ (_04132_, _04131_, _04130_);
  and _26602_ (_04133_, _04132_, _13828_);
  and _26603_ (_04134_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _26604_ (_04135_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26605_ (_04136_, _04135_, _04134_);
  and _26606_ (_04137_, _04136_, _12426_);
  or _26607_ (_04138_, _04137_, _04133_);
  or _26608_ (_04139_, _04138_, _04129_);
  or _26609_ (_04140_, _04139_, _04125_);
  and _26610_ (_04141_, _04140_, _04120_);
  and _26611_ (_04142_, _13847_, _12030_);
  and _26612_ (_04143_, _13874_, _12030_);
  nor _26613_ (_04145_, _04143_, _04142_);
  and _26614_ (_04147_, _13887_, _12030_);
  and _26615_ (_04148_, _04147_, _13816_);
  or _26616_ (_04149_, _13838_, _13819_);
  and _26617_ (_04150_, _04149_, _13837_);
  nor _26618_ (_04151_, _04150_, _04148_);
  and _26619_ (_04152_, _04151_, _04145_);
  not _26620_ (_04153_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _26621_ (_04155_, _04120_, _04153_);
  and _26622_ (_04156_, _13817_, _13819_);
  and _26623_ (_04158_, _04147_, _13883_);
  nor _26624_ (_04160_, _04158_, _04156_);
  and _26625_ (_04161_, _04160_, _04155_);
  and _26626_ (_04162_, _04161_, _04152_);
  and _26627_ (_04163_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _26628_ (_04165_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _26629_ (_04167_, _04165_, _04163_);
  and _26630_ (_04169_, _04167_, _13842_);
  or _26631_ (_04170_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _26632_ (_04171_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _26633_ (_04172_, _04171_, _13831_);
  and _26634_ (_04173_, _04172_, _04170_);
  nor _26635_ (_04174_, _12426_, _01916_);
  and _26636_ (_04175_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _26637_ (_04176_, _04175_, _04174_);
  and _26638_ (_04177_, _04176_, _13818_);
  nand _26639_ (_04178_, _12426_, _06056_);
  or _26640_ (_04179_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _26641_ (_04180_, _04179_, _13828_);
  and _26642_ (_04181_, _04180_, _04178_);
  or _26643_ (_04182_, _04181_, _04177_);
  or _26644_ (_04183_, _04182_, _04173_);
  or _26645_ (_04185_, _04183_, _04169_);
  and _26646_ (_04187_, _04185_, _04156_);
  or _26647_ (_04188_, _04187_, _04162_);
  and _26648_ (_04189_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _26649_ (_04190_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _26650_ (_04191_, _04190_, _04189_);
  and _26651_ (_04192_, _04191_, _13849_);
  nor _26652_ (_04193_, _12426_, _01786_);
  and _26653_ (_04195_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _26654_ (_04196_, _04195_, _04193_);
  and _26655_ (_04198_, _04196_, _13818_);
  nor _26656_ (_04200_, _12426_, _01815_);
  and _26657_ (_04202_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _26658_ (_04203_, _04202_, _04200_);
  and _26659_ (_04204_, _04203_, _13831_);
  or _26660_ (_04205_, _04204_, _04198_);
  and _26661_ (_04206_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _26662_ (_04207_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _26663_ (_04208_, _04207_, _04206_);
  and _26664_ (_04209_, _04208_, _12426_);
  or _26665_ (_04210_, _04209_, _04205_);
  or _26666_ (_04211_, _04210_, _04192_);
  and _26667_ (_04212_, _04211_, _04158_);
  and _26668_ (_04213_, _00070_, _13831_);
  and _26669_ (_04214_, _00229_, _13818_);
  or _26670_ (_04215_, _04214_, _04213_);
  and _26671_ (_04216_, _04215_, _12426_);
  or _26672_ (_04217_, _00005_, _13849_);
  or _26673_ (_04219_, _04022_, _12426_);
  and _26674_ (_04220_, _04219_, _13842_);
  and _26675_ (_04221_, _04220_, _04217_);
  or _26676_ (_04222_, _00139_, _13849_);
  or _26677_ (_04223_, _03362_, _12426_);
  and _26678_ (_04224_, _04223_, _13828_);
  and _26679_ (_04225_, _04224_, _04222_);
  or _26680_ (_04226_, _04225_, _04221_);
  and _26681_ (_04227_, _03473_, _13831_);
  and _26682_ (_04228_, _03612_, _13818_);
  or _26683_ (_04229_, _04228_, _04227_);
  and _26684_ (_04230_, _04229_, _13849_);
  or _26685_ (_04232_, _04230_, _04226_);
  or _26686_ (_04233_, _04232_, _04216_);
  and _26687_ (_04234_, _04233_, _04143_);
  or _26688_ (_04235_, _04234_, _04212_);
  and _26689_ (_04236_, _12432_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _26690_ (_04237_, _13839_, _12030_);
  and _26691_ (_04238_, _03366_, _13828_);
  and _26692_ (_04239_, _03608_, _13818_);
  or _26693_ (_04240_, _04239_, _04238_);
  and _26694_ (_04241_, _04240_, _13849_);
  and _26695_ (_04242_, _00135_, _13828_);
  and _26696_ (_04243_, _00224_, _13818_);
  or _26697_ (_04244_, _04243_, _04242_);
  and _26698_ (_04245_, _04244_, _12426_);
  or _26699_ (_04246_, _14005_, _13849_);
  or _26700_ (_04247_, _04018_, _12426_);
  and _26701_ (_04248_, _04247_, _13842_);
  and _26702_ (_04250_, _04248_, _04246_);
  or _26703_ (_04251_, _00066_, _13849_);
  or _26704_ (_04252_, _03468_, _12426_);
  and _26705_ (_04253_, _04252_, _13831_);
  and _26706_ (_04254_, _04253_, _04251_);
  or _26707_ (_04255_, _04254_, _04250_);
  or _26708_ (_04256_, _04255_, _04245_);
  or _26709_ (_04257_, _04256_, _04241_);
  and _26710_ (_04258_, _04257_, _04237_);
  or _26711_ (_04259_, _04258_, _04236_);
  or _26712_ (_04260_, _04259_, _04235_);
  or _26713_ (_04261_, _04260_, _04188_);
  and _26714_ (_04262_, _13988_, _13842_);
  and _26715_ (_04263_, _00218_, _13818_);
  or _26716_ (_04264_, _04263_, _04262_);
  and _26717_ (_04265_, _00148_, _13828_);
  and _26718_ (_04266_, _00075_, _13831_);
  or _26719_ (_04267_, _04266_, _04265_);
  or _26720_ (_04268_, _04267_, _04264_);
  and _26721_ (_04269_, _04268_, _13846_);
  and _26722_ (_04270_, _00144_, _13828_);
  and _26723_ (_04271_, _00079_, _13831_);
  or _26724_ (_04272_, _04271_, _04270_);
  and _26725_ (_04273_, _13997_, _13842_);
  and _26726_ (_04274_, _00213_, _13818_);
  or _26727_ (_04275_, _04274_, _04273_);
  or _26728_ (_04276_, _04275_, _04272_);
  and _26729_ (_04277_, _04276_, _12221_);
  or _26730_ (_04278_, _04277_, _04269_);
  and _26731_ (_04279_, _04278_, _12426_);
  and _26732_ (_04280_, _04009_, _13842_);
  and _26733_ (_04281_, _03623_, _13818_);
  or _26734_ (_04282_, _04281_, _04280_);
  and _26735_ (_04283_, _03375_, _13828_);
  and _26736_ (_04284_, _03459_, _13831_);
  or _26737_ (_04285_, _04284_, _04283_);
  or _26738_ (_04286_, _04285_, _04282_);
  and _26739_ (_04287_, _04286_, _12221_);
  and _26740_ (_04288_, _04013_, _13842_);
  and _26741_ (_04289_, _03619_, _13818_);
  or _26742_ (_04290_, _04289_, _04288_);
  and _26743_ (_04291_, _03371_, _13828_);
  and _26744_ (_04292_, _03463_, _13831_);
  or _26745_ (_04293_, _04292_, _04291_);
  or _26746_ (_04294_, _04293_, _04290_);
  and _26747_ (_04295_, _04294_, _13846_);
  or _26748_ (_04296_, _04295_, _04287_);
  and _26749_ (_04297_, _04296_, _13849_);
  or _26750_ (_04298_, _04297_, _04279_);
  and _26751_ (_04299_, _04298_, _04142_);
  nor _26752_ (_04300_, _12426_, _01030_);
  and _26753_ (_04301_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _26754_ (_04302_, _04301_, _04300_);
  and _26755_ (_04303_, _04302_, _13818_);
  or _26756_ (_04304_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _26757_ (_04305_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _26758_ (_04306_, _04305_, _13828_);
  and _26759_ (_04307_, _04306_, _04304_);
  or _26760_ (_04308_, _04307_, _04303_);
  nor _26761_ (_04309_, _12426_, _00764_);
  and _26762_ (_04310_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _26763_ (_04311_, _04310_, _04309_);
  and _26764_ (_04312_, _04311_, _13831_);
  or _26765_ (_04313_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _26766_ (_04314_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _26767_ (_04315_, _04314_, _13842_);
  and _26768_ (_04316_, _04315_, _04313_);
  or _26769_ (_04317_, _04316_, _04312_);
  or _26770_ (_04318_, _04317_, _04308_);
  and _26771_ (_04319_, _04318_, _13839_);
  nor _26772_ (_04320_, _12426_, _06464_);
  and _26773_ (_04321_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _26774_ (_04322_, _04321_, _04320_);
  and _26775_ (_04323_, _04322_, _13818_);
  or _26776_ (_04324_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _26777_ (_04325_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _26778_ (_04326_, _04325_, _13828_);
  and _26779_ (_04327_, _04326_, _04324_);
  or _26780_ (_04328_, _04327_, _04323_);
  and _26781_ (_04329_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _26782_ (_04330_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _26783_ (_04331_, _04330_, _04329_);
  and _26784_ (_04332_, _04331_, _13831_);
  or _26785_ (_04333_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _26786_ (_04334_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _26787_ (_04335_, _04334_, _13842_);
  and _26788_ (_04336_, _04335_, _04333_);
  or _26789_ (_04337_, _04336_, _04332_);
  or _26790_ (_04338_, _04337_, _04328_);
  and _26791_ (_04339_, _04338_, _13853_);
  or _26792_ (_04340_, _04339_, _04319_);
  and _26793_ (_04341_, _04340_, _13819_);
  and _26794_ (_04342_, _13848_, _13819_);
  nand _26795_ (_04343_, _12426_, _06495_);
  or _26796_ (_04344_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _26797_ (_04345_, _04344_, _13828_);
  and _26798_ (_04346_, _04345_, _04343_);
  nand _26799_ (_04347_, _12426_, _06489_);
  or _26800_ (_04348_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _26801_ (_04349_, _04348_, _13818_);
  and _26802_ (_04350_, _04349_, _04347_);
  or _26803_ (_04351_, _04350_, _04346_);
  or _26804_ (_04352_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand _26805_ (_04353_, _12426_, _06492_);
  and _26806_ (_04354_, _04353_, _13831_);
  and _26807_ (_04356_, _04354_, _04352_);
  or _26808_ (_04357_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand _26809_ (_04358_, _12426_, _06482_);
  and _26810_ (_04359_, _04358_, _13842_);
  and _26811_ (_04360_, _04359_, _04357_);
  or _26812_ (_04362_, _04360_, _04356_);
  or _26813_ (_04363_, _04362_, _04351_);
  and _26814_ (_04364_, _04363_, _04342_);
  and _26815_ (_04365_, _13874_, _13819_);
  nor _26816_ (_04366_, _12426_, _13703_);
  and _26817_ (_04367_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _26818_ (_04369_, _04367_, _04366_);
  and _26819_ (_04370_, _04369_, _13828_);
  nand _26820_ (_04372_, _12426_, _07907_);
  or _26821_ (_04374_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _26822_ (_04375_, _04374_, _13818_);
  and _26823_ (_04376_, _04375_, _04372_);
  or _26824_ (_04377_, _04376_, _04370_);
  or _26825_ (_04378_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _26826_ (_04379_, _12426_, _13746_);
  and _26827_ (_04380_, _04379_, _13842_);
  and _26828_ (_04381_, _04380_, _04378_);
  or _26829_ (_04382_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand _26830_ (_04383_, _12426_, _00435_);
  and _26831_ (_04384_, _04383_, _13831_);
  and _26832_ (_04385_, _04384_, _04382_);
  or _26833_ (_04386_, _04385_, _04381_);
  or _26834_ (_04387_, _04386_, _04377_);
  and _26835_ (_04388_, _04387_, _04365_);
  and _26836_ (_04389_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _26837_ (_04390_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _26838_ (_04391_, _04390_, _04389_);
  and _26839_ (_04392_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _26840_ (_04393_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _26841_ (_04394_, _04393_, _04392_);
  or _26842_ (_04395_, _04394_, _04391_);
  and _26843_ (_04396_, _04395_, _13849_);
  and _26844_ (_04397_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _26845_ (_04398_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _26846_ (_04399_, _04398_, _04397_);
  and _26847_ (_04400_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _26848_ (_04401_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _26849_ (_04402_, _04401_, _04400_);
  or _26850_ (_04403_, _04402_, _04399_);
  and _26851_ (_04404_, _04403_, _12426_);
  or _26852_ (_04405_, _04404_, _04396_);
  and _26853_ (_04406_, _04405_, _04148_);
  or _26854_ (_04407_, _04406_, _04388_);
  or _26855_ (_04408_, _04407_, _04364_);
  or _26856_ (_04409_, _04408_, _04341_);
  or _26857_ (_04410_, _04409_, _04299_);
  or _26858_ (_04411_, _04410_, _04261_);
  or _26859_ (_04412_, _04411_, _04141_);
  and _26860_ (_04413_, _04148_, _07766_);
  nor _26861_ (_04414_, _04413_, _12231_);
  nand _26862_ (_04415_, _04236_, _06803_);
  and _26863_ (_04416_, _04415_, _04414_);
  and _26864_ (_04417_, _04416_, _04412_);
  and _26865_ (_04418_, _13842_, _06360_);
  and _26866_ (_04419_, _13831_, _12120_);
  or _26867_ (_04420_, _04419_, _04418_);
  and _26868_ (_04421_, _04420_, _13849_);
  and _26869_ (_04422_, _13842_, _12019_);
  and _26870_ (_04423_, _13831_, _06435_);
  or _26871_ (_04424_, _04423_, _04422_);
  and _26872_ (_04425_, _04424_, _12426_);
  nor _26873_ (_04426_, _12426_, _06609_);
  and _26874_ (_04427_, _12426_, _11023_);
  or _26875_ (_04428_, _04427_, _04426_);
  and _26876_ (_04429_, _04428_, _13828_);
  nor _26877_ (_04430_, _12426_, _06993_);
  and _26878_ (_04431_, _12426_, _07978_);
  or _26879_ (_04432_, _04431_, _04430_);
  and _26880_ (_04433_, _04432_, _13818_);
  or _26881_ (_04434_, _04433_, _04429_);
  or _26882_ (_04435_, _04434_, _04425_);
  nor _26883_ (_04436_, _04435_, _04421_);
  nor _26884_ (_04438_, _04436_, _04414_);
  or _26885_ (_04439_, _04438_, _04417_);
  and _26886_ (_04186_, _04439_, _06071_);
  nor _26887_ (_04440_, _00426_, rst);
  or _26888_ (_04441_, _00425_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _26889_ (_04442_, _00425_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _26890_ (_04443_, _04442_, _04441_);
  and _26891_ (_04194_, _04443_, _04440_);
  or _26892_ (_04444_, _03703_, _13340_);
  and _26893_ (_04445_, _04444_, _06527_);
  nand _26894_ (_04446_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand _26895_ (_04447_, _04446_, _11819_);
  or _26896_ (_04448_, _04447_, _04445_);
  and _26897_ (_04197_, _04448_, _06071_);
  and _26898_ (_04449_, _11889_, _13378_);
  or _26899_ (_04450_, _04449_, _03950_);
  or _26900_ (_04451_, _04450_, _11917_);
  or _26901_ (_04452_, _04451_, _03883_);
  or _26902_ (_04453_, _04452_, _04058_);
  or _26903_ (_04454_, _03658_, _13976_);
  or _26904_ (_04455_, _04454_, _13630_);
  or _26905_ (_04456_, _04455_, _04453_);
  or _26906_ (_04457_, _04456_, _03655_);
  and _26907_ (_04458_, _04457_, _06527_);
  and _26908_ (_04459_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26909_ (_04460_, _04459_, _03664_);
  or _26910_ (_04461_, _04460_, _04458_);
  and _26911_ (_04201_, _04461_, _06071_);
  or _26912_ (_04463_, _04093_, _03883_);
  or _26913_ (_04465_, _04463_, _03898_);
  or _26914_ (_04466_, _13337_, _11868_);
  or _26915_ (_04467_, _13633_, _03876_);
  or _26916_ (_04468_, _04467_, _04466_);
  or _26917_ (_04469_, _03526_, _13345_);
  or _26918_ (_04470_, _04469_, _04468_);
  or _26919_ (_04471_, _11869_, _11837_);
  or _26920_ (_04472_, _03888_, _04471_);
  or _26921_ (_04473_, _04472_, _04470_);
  or _26922_ (_04474_, _04473_, _04465_);
  and _26923_ (_04475_, _04474_, _06527_);
  and _26924_ (_04476_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _26925_ (_04478_, _04476_, _11818_);
  or _26926_ (_04479_, _04478_, _04475_);
  and _26927_ (_04218_, _04479_, _06071_);
  or _26928_ (_04481_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _26929_ (_04482_, _03792_, rst);
  and _26930_ (_04231_, _04482_, _04481_);
  nand _26931_ (_04483_, _07759_, _07715_);
  or _26932_ (_04484_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _26933_ (_04485_, _04484_, _06071_);
  and _26934_ (_04249_, _04485_, _04483_);
  nand _26935_ (_04486_, _08988_, _06359_);
  and _26936_ (_04487_, _04486_, _06071_);
  and _26937_ (_04488_, _02646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _26938_ (_04489_, _04488_, _02647_);
  nand _26939_ (_04490_, _04489_, _09028_);
  nor _26940_ (_04491_, _12295_, _06803_);
  and _26941_ (_04492_, _12295_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _26942_ (_04493_, _04492_, _04491_);
  or _26943_ (_04494_, _04493_, _09028_);
  and _26944_ (_04495_, _04494_, _04490_);
  or _26945_ (_04496_, _04495_, _08988_);
  and _26946_ (_04355_, _04496_, _04487_);
  nor _26947_ (_04497_, _13738_, _13778_);
  and _26948_ (_04498_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _26949_ (_04499_, _04498_, _04497_);
  and _26950_ (_04500_, _04499_, _13798_);
  nand _26951_ (_04501_, _07885_, _06359_);
  nand _26952_ (_04502_, _09341_, _07902_);
  and _26953_ (_04503_, _04502_, _02727_);
  and _26954_ (_04504_, _04503_, _04501_);
  or _26955_ (_04361_, _04504_, _04500_);
  and _26956_ (_04505_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _26957_ (_04506_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _26958_ (_04507_, _04506_, _04505_);
  or _26959_ (_04508_, _04507_, _13744_);
  and _26960_ (_04509_, _04508_, _06071_);
  nand _26961_ (_04510_, _13759_, _06359_);
  and _26962_ (_04368_, _04510_, _04509_);
  and _26963_ (_04511_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _26964_ (_04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _26965_ (_04513_, pc_log_change, _04512_);
  or _26966_ (_04514_, _04513_, _04511_);
  and _26967_ (_04371_, _04514_, _06071_);
  nand _26968_ (_04515_, _13723_, _07977_);
  or _26969_ (_04516_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _26970_ (_04517_, _04516_, _06071_);
  and _26971_ (_04373_, _04517_, _04515_);
  not _26972_ (_04518_, _06054_);
  and _26973_ (_04519_, _06059_, _04518_);
  and _26974_ (_04520_, _04519_, _06036_);
  not _26975_ (_04521_, _04520_);
  or _26976_ (_04522_, _04521_, _06053_);
  or _26977_ (_04523_, _04520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _26978_ (_04524_, _04523_, _06071_);
  and _26979_ (_04437_, _04524_, _04522_);
  and _26980_ (_04525_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _26981_ (_04526_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _26982_ (_04527_, _04526_, _04525_);
  and _26983_ (_04528_, _04527_, _13798_);
  nand _26984_ (_04529_, _09037_, _07885_);
  nand _26985_ (_04530_, _07977_, _07902_);
  and _26986_ (_04531_, _04530_, _02727_);
  and _26987_ (_04532_, _04531_, _04529_);
  or _26988_ (_04462_, _04532_, _04528_);
  and _26989_ (_04533_, _13759_, _11023_);
  and _26990_ (_04534_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _26991_ (_04535_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _26992_ (_04536_, _04535_, _04534_);
  nor _26993_ (_04537_, _04536_, _13744_);
  and _26994_ (_04538_, _13753_, _06435_);
  or _26995_ (_04539_, _04538_, _04537_);
  or _26996_ (_04540_, _04539_, _04533_);
  and _26997_ (_04464_, _04540_, _06071_);
  nand _26998_ (_04541_, _13723_, _06609_);
  or _26999_ (_04542_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _27000_ (_04543_, _04542_, _06071_);
  and _27001_ (_04477_, _04543_, _04541_);
  nand _27002_ (_04544_, _13723_, _06993_);
  or _27003_ (_04545_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _27004_ (_04546_, _04545_, _06071_);
  and _27005_ (_04480_, _04546_, _04544_);
  and _27006_ (_04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27007_ (_04548_, _04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27008_ (_04549_, _04548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _27009_ (_04550_, _04549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _27010_ (_04551_, _04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _27011_ (_04552_, _04551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _27012_ (_04553_, _04552_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _27013_ (_04554_, _04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _27014_ (_04555_, _04554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _27015_ (_04556_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _27016_ (_04557_, _04556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _27017_ (_04558_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _27018_ (_04559_, _04558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _27019_ (_04560_, _04558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _27020_ (_04561_, _04560_, _04559_);
  and _27021_ (_04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _27022_ (_04563_, _04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27023_ (_04564_, _04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27024_ (_04565_, _04564_, _04563_);
  and _27025_ (_04566_, _02453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27026_ (_04567_, _04566_);
  nor _27027_ (_04568_, _04563_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27028_ (_04569_, _04563_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27029_ (_04570_, _04569_, _04568_);
  nor _27030_ (_04571_, _04570_, _08210_);
  and _27031_ (_04572_, _04570_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _27032_ (_04573_, _04572_, _04571_);
  or _27033_ (_04574_, _04573_, _04567_);
  nor _27034_ (_04575_, _04570_, _08176_);
  and _27035_ (_04576_, _04570_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _27036_ (_04577_, _04576_, _04575_);
  nor _27037_ (_04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27038_ (_04579_, _04578_);
  or _27039_ (_04580_, _04579_, _04577_);
  and _27040_ (_04581_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01884_);
  not _27041_ (_04582_, _04581_);
  nor _27042_ (_04583_, _04570_, _08240_);
  and _27043_ (_04584_, _04570_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _27044_ (_04585_, _04584_, _04583_);
  or _27045_ (_04586_, _04585_, _04582_);
  and _27046_ (_04587_, _04586_, _04580_);
  and _27047_ (_04588_, _04587_, _04574_);
  or _27048_ (_04589_, _04588_, _04565_);
  not _27049_ (_04590_, _04563_);
  not _27050_ (_04591_, _04570_);
  and _27051_ (_04592_, _04591_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27052_ (_04593_, _04570_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _27053_ (_04594_, _04593_, _04592_);
  or _27054_ (_04595_, _04594_, _04590_);
  not _27055_ (_04596_, _04565_);
  and _27056_ (_04597_, _04570_, _08228_);
  or _27057_ (_04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  nand _27058_ (_04599_, _04598_, _04581_);
  or _27059_ (_04600_, _04599_, _04597_);
  and _27060_ (_04601_, _04570_, _08233_);
  or _27061_ (_04602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nand _27062_ (_04603_, _04602_, _04562_);
  or _27063_ (_04604_, _04603_, _04601_);
  and _27064_ (_04605_, _04604_, _04600_);
  and _27065_ (_04606_, _04570_, _08215_);
  or _27066_ (_04607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _27067_ (_04608_, _04607_, _04578_);
  or _27068_ (_04609_, _04608_, _04606_);
  and _27069_ (_04610_, _04570_, _08203_);
  or _27070_ (_04611_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _27071_ (_04612_, _04611_, _04566_);
  or _27072_ (_04613_, _04612_, _04610_);
  and _27073_ (_04614_, _04613_, _04609_);
  and _27074_ (_04615_, _04614_, _04605_);
  or _27075_ (_04616_, _04615_, _04596_);
  and _27076_ (_04617_, _04616_, _04595_);
  and _27077_ (_04618_, _04617_, _04589_);
  and _27078_ (_04619_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _27079_ (_04620_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _27080_ (_04621_, _04620_, _04619_);
  and _27081_ (_04622_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _27082_ (_04623_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _27083_ (_04624_, _04623_, _04622_);
  and _27084_ (_04625_, _04624_, _04621_);
  and _27085_ (_04626_, _04625_, _04596_);
  and _27086_ (_04627_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _27087_ (_04628_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _27088_ (_04629_, _04628_, _04627_);
  and _27089_ (_04630_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _27090_ (_04631_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _27091_ (_04632_, _04631_, _04630_);
  and _27092_ (_04633_, _04632_, _04629_);
  and _27093_ (_04634_, _04633_, _04565_);
  or _27094_ (_04635_, _04634_, _04591_);
  nor _27095_ (_04636_, _04635_, _04626_);
  and _27096_ (_04637_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _27097_ (_04638_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor _27098_ (_04639_, _04638_, _04637_);
  and _27099_ (_04640_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _27100_ (_04641_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _27101_ (_04642_, _04641_, _04640_);
  and _27102_ (_04643_, _04642_, _04639_);
  nor _27103_ (_04644_, _04643_, _04565_);
  and _27104_ (_04645_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _27105_ (_04646_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _27106_ (_04647_, _04646_, _04645_);
  and _27107_ (_04648_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _27108_ (_04649_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _27109_ (_04650_, _04649_, _04648_);
  and _27110_ (_04651_, _04650_, _04647_);
  nor _27111_ (_04652_, _04651_, _04596_);
  or _27112_ (_04653_, _04652_, _04644_);
  and _27113_ (_04654_, _04653_, _04591_);
  nor _27114_ (_04655_, _04654_, _04636_);
  nor _27115_ (_04656_, _04655_, _04618_);
  nor _27116_ (_04657_, _04556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _27117_ (_04658_, _04657_, _04557_);
  and _27118_ (_04659_, _04658_, _04656_);
  and _27119_ (_04660_, _04659_, _02142_);
  nor _27120_ (_04661_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _27121_ (_04662_, _04661_, _04558_);
  and _27122_ (_04663_, _04662_, _04656_);
  nor _27123_ (_04664_, _04662_, _04656_);
  nor _27124_ (_04665_, _04664_, _04663_);
  nor _27125_ (_04666_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _27126_ (_04667_, _04666_, _04556_);
  and _27127_ (_04668_, _04667_, _04656_);
  nor _27128_ (_04669_, _04554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _27129_ (_04670_, _04669_, _04555_);
  and _27130_ (_04671_, _04670_, _04656_);
  nor _27131_ (_04672_, _04667_, _04656_);
  nor _27132_ (_04673_, _04672_, _04668_);
  nor _27133_ (_04674_, _04670_, _04656_);
  nor _27134_ (_04675_, _04674_, _04671_);
  not _27135_ (_04676_, _04675_);
  nor _27136_ (_04677_, _04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _27137_ (_04678_, _04677_, _04554_);
  and _27138_ (_04679_, _04678_, _04656_);
  nor _27139_ (_04680_, _04552_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _27140_ (_04681_, _04680_, _04553_);
  and _27141_ (_04682_, _04681_, _04656_);
  nor _27142_ (_04683_, _04678_, _04656_);
  nor _27143_ (_04684_, _04683_, _04679_);
  nor _27144_ (_04685_, _04551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _27145_ (_04686_, _04685_, _04552_);
  and _27146_ (_04687_, _04686_, _04656_);
  nor _27147_ (_04688_, _04686_, _04656_);
  and _27148_ (_04689_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _27149_ (_04690_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _27150_ (_04691_, _04690_, _04689_);
  and _27151_ (_04692_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _27152_ (_04693_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _27153_ (_04694_, _04693_, _04692_);
  and _27154_ (_04695_, _04694_, _04691_);
  nor _27155_ (_04696_, _04695_, _04565_);
  and _27156_ (_04697_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _27157_ (_04698_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _27158_ (_04699_, _04698_, _04697_);
  and _27159_ (_04700_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _27160_ (_04701_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _27161_ (_04702_, _04701_, _04700_);
  and _27162_ (_04703_, _04702_, _04699_);
  nor _27163_ (_04704_, _04703_, _04596_);
  or _27164_ (_04705_, _04704_, _04696_);
  and _27165_ (_04706_, _04705_, _04570_);
  and _27166_ (_04707_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _27167_ (_04708_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _27168_ (_04709_, _04708_, _04707_);
  and _27169_ (_04710_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _27170_ (_04711_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _27171_ (_04712_, _04711_, _04710_);
  and _27172_ (_04713_, _04712_, _04709_);
  nor _27173_ (_04714_, _04713_, _04565_);
  and _27174_ (_04715_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _27175_ (_04716_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _27176_ (_04717_, _04716_, _04715_);
  and _27177_ (_04718_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _27178_ (_04719_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _27179_ (_04720_, _04719_, _04718_);
  and _27180_ (_04721_, _04720_, _04717_);
  nor _27181_ (_04722_, _04721_, _04596_);
  or _27182_ (_04723_, _04722_, _04714_);
  and _27183_ (_04724_, _04723_, _04591_);
  nor _27184_ (_04725_, _04724_, _04706_);
  nor _27185_ (_04726_, _04725_, _04618_);
  nor _27186_ (_04727_, _04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _27187_ (_04728_, _04727_, _04551_);
  and _27188_ (_04729_, _04728_, _04726_);
  nor _27189_ (_04730_, _04728_, _04726_);
  nor _27190_ (_04731_, _04730_, _04729_);
  not _27191_ (_04732_, _04731_);
  and _27192_ (_04733_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _27193_ (_04734_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _27194_ (_04735_, _04734_, _04733_);
  and _27195_ (_04736_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _27196_ (_04737_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _27197_ (_04738_, _04737_, _04736_);
  and _27198_ (_04739_, _04738_, _04735_);
  and _27199_ (_04740_, _04739_, _04596_);
  and _27200_ (_04741_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _27201_ (_04742_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _27202_ (_04743_, _04742_, _04741_);
  and _27203_ (_04744_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _27204_ (_04745_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _27205_ (_04746_, _04745_, _04744_);
  and _27206_ (_04747_, _04746_, _04743_);
  and _27207_ (_04748_, _04747_, _04565_);
  or _27208_ (_04749_, _04748_, _04591_);
  nor _27209_ (_04750_, _04749_, _04740_);
  and _27210_ (_04751_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _27211_ (_04752_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _27212_ (_04753_, _04752_, _04751_);
  and _27213_ (_04754_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _27214_ (_04755_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _27215_ (_04756_, _04755_, _04754_);
  and _27216_ (_04757_, _04756_, _04753_);
  nor _27217_ (_04758_, _04757_, _04565_);
  and _27218_ (_04759_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _27219_ (_04760_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _27220_ (_04761_, _04760_, _04759_);
  and _27221_ (_04762_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _27222_ (_04763_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _27223_ (_04764_, _04763_, _04762_);
  and _27224_ (_04765_, _04764_, _04761_);
  nor _27225_ (_04766_, _04765_, _04596_);
  or _27226_ (_04767_, _04766_, _04758_);
  and _27227_ (_04768_, _04767_, _04591_);
  nor _27228_ (_04769_, _04768_, _04750_);
  nor _27229_ (_04770_, _04769_, _04618_);
  nor _27230_ (_04771_, _04549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _27231_ (_04772_, _04771_, _04550_);
  and _27232_ (_04773_, _04772_, _04770_);
  nor _27233_ (_04774_, _04772_, _04770_);
  nor _27234_ (_04775_, _04774_, _04773_);
  not _27235_ (_04776_, _04775_);
  and _27236_ (_04777_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _27237_ (_04778_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _27238_ (_04779_, _04778_, _04777_);
  and _27239_ (_04780_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _27240_ (_04781_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _27241_ (_04782_, _04781_, _04780_);
  and _27242_ (_04783_, _04782_, _04779_);
  and _27243_ (_04784_, _04783_, _04596_);
  and _27244_ (_04785_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _27245_ (_04786_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _27246_ (_04787_, _04786_, _04785_);
  and _27247_ (_04788_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _27248_ (_04789_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _27249_ (_04790_, _04789_, _04788_);
  and _27250_ (_04791_, _04790_, _04787_);
  and _27251_ (_04792_, _04791_, _04565_);
  or _27252_ (_04793_, _04792_, _04570_);
  nor _27253_ (_04794_, _04793_, _04784_);
  and _27254_ (_04795_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _27255_ (_04796_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _27256_ (_04797_, _04796_, _04795_);
  and _27257_ (_04798_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _27258_ (_04799_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _27259_ (_04800_, _04799_, _04798_);
  and _27260_ (_04801_, _04800_, _04797_);
  and _27261_ (_04802_, _04801_, _04596_);
  and _27262_ (_04803_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _27263_ (_04804_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _27264_ (_04805_, _04804_, _04803_);
  and _27265_ (_04806_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _27266_ (_04807_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _27267_ (_04808_, _04807_, _04806_);
  and _27268_ (_04809_, _04808_, _04805_);
  and _27269_ (_04810_, _04809_, _04565_);
  or _27270_ (_04811_, _04810_, _04591_);
  nor _27271_ (_04812_, _04811_, _04802_);
  nor _27272_ (_04813_, _04812_, _04794_);
  nor _27273_ (_04814_, _04813_, _04618_);
  nor _27274_ (_04815_, _04548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _27275_ (_04816_, _04815_, _04549_);
  and _27276_ (_04817_, _04816_, _04814_);
  and _27277_ (_04818_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _27278_ (_04819_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _27279_ (_04820_, _04819_, _04818_);
  and _27280_ (_04821_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _27281_ (_04822_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _27282_ (_04823_, _04822_, _04821_);
  and _27283_ (_04824_, _04823_, _04820_);
  and _27284_ (_04825_, _04824_, _04596_);
  and _27285_ (_04826_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _27286_ (_04827_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _27287_ (_04828_, _04827_, _04826_);
  and _27288_ (_04829_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _27289_ (_04830_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _27290_ (_04831_, _04830_, _04829_);
  and _27291_ (_04832_, _04831_, _04828_);
  and _27292_ (_04833_, _04832_, _04565_);
  or _27293_ (_04834_, _04833_, _04591_);
  nor _27294_ (_04835_, _04834_, _04825_);
  and _27295_ (_04836_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _27296_ (_04837_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _27297_ (_04838_, _04837_, _04836_);
  and _27298_ (_04839_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _27299_ (_04840_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _27300_ (_04841_, _04840_, _04839_);
  and _27301_ (_04842_, _04841_, _04838_);
  nor _27302_ (_04843_, _04842_, _04565_);
  and _27303_ (_04844_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _27304_ (_04845_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _27305_ (_04846_, _04845_, _04844_);
  and _27306_ (_04847_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _27307_ (_04848_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _27308_ (_04849_, _04848_, _04847_);
  and _27309_ (_04850_, _04849_, _04846_);
  nor _27310_ (_04851_, _04850_, _04596_);
  or _27311_ (_04852_, _04851_, _04843_);
  and _27312_ (_04853_, _04852_, _04591_);
  nor _27313_ (_04854_, _04853_, _04835_);
  nor _27314_ (_04855_, _04854_, _04618_);
  nor _27315_ (_04856_, _04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27316_ (_04857_, _04856_, _04548_);
  and _27317_ (_04858_, _04857_, _04855_);
  nor _27318_ (_04859_, _04857_, _04855_);
  and _27319_ (_04860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02461_);
  and _27320_ (_04861_, _01884_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27321_ (_04862_, _04861_, _04860_);
  not _27322_ (_04863_, _04862_);
  and _27323_ (_04864_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _27324_ (_04865_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _27325_ (_04866_, _04865_, _04864_);
  and _27326_ (_04867_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _27327_ (_04868_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _27328_ (_04869_, _04868_, _04867_);
  and _27329_ (_04870_, _04869_, _04866_);
  nor _27330_ (_04871_, _04870_, _04565_);
  and _27331_ (_04872_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _27332_ (_04873_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _27333_ (_04874_, _04873_, _04872_);
  and _27334_ (_04875_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _27335_ (_04876_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _27336_ (_04877_, _04876_, _04875_);
  and _27337_ (_04878_, _04877_, _04874_);
  nor _27338_ (_04879_, _04878_, _04596_);
  or _27339_ (_04880_, _04879_, _04871_);
  and _27340_ (_04881_, _04880_, _04570_);
  and _27341_ (_04882_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _27342_ (_04883_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _27343_ (_04884_, _04883_, _04882_);
  and _27344_ (_04885_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _27345_ (_04886_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _27346_ (_04887_, _04886_, _04885_);
  and _27347_ (_04888_, _04887_, _04884_);
  nor _27348_ (_04889_, _04888_, _04565_);
  and _27349_ (_04890_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _27350_ (_04891_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _27351_ (_04892_, _04891_, _04890_);
  and _27352_ (_04893_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _27353_ (_04894_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _27354_ (_04895_, _04894_, _04893_);
  and _27355_ (_04896_, _04895_, _04892_);
  nor _27356_ (_04897_, _04896_, _04596_);
  or _27357_ (_04898_, _04897_, _04889_);
  and _27358_ (_04899_, _04898_, _04591_);
  nor _27359_ (_04900_, _04899_, _04881_);
  nor _27360_ (_04901_, _04900_, _04618_);
  and _27361_ (_04902_, _04901_, _04863_);
  and _27362_ (_04903_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _27363_ (_04904_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _27364_ (_04905_, _04904_, _04903_);
  and _27365_ (_04906_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _27366_ (_04907_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _27367_ (_04908_, _04907_, _04906_);
  and _27368_ (_04909_, _04908_, _04905_);
  nor _27369_ (_04910_, _04909_, _04565_);
  and _27370_ (_04911_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _27371_ (_04912_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _27372_ (_04913_, _04912_, _04911_);
  and _27373_ (_04914_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _27374_ (_04915_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _27375_ (_04916_, _04915_, _04914_);
  and _27376_ (_04917_, _04916_, _04913_);
  nor _27377_ (_04918_, _04917_, _04596_);
  or _27378_ (_04919_, _04918_, _04910_);
  and _27379_ (_04920_, _04919_, _04591_);
  and _27380_ (_04921_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _27381_ (_04922_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _27382_ (_04923_, _04922_, _04921_);
  and _27383_ (_04924_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _27384_ (_04925_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _27385_ (_04926_, _04925_, _04924_);
  and _27386_ (_04927_, _04926_, _04923_);
  nor _27387_ (_04928_, _04927_, _04596_);
  and _27388_ (_04929_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _27389_ (_04930_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _27390_ (_04931_, _04930_, _04929_);
  and _27391_ (_04932_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _27392_ (_04933_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _27393_ (_04934_, _04933_, _04932_);
  and _27394_ (_04935_, _04934_, _04931_);
  nor _27395_ (_04936_, _04935_, _04565_);
  nor _27396_ (_04937_, _04936_, _04928_);
  nor _27397_ (_04938_, _04937_, _04591_);
  nor _27398_ (_04939_, _04938_, _04920_);
  nor _27399_ (_04940_, _04939_, _04618_);
  and _27400_ (_04941_, _04940_, _01884_);
  and _27401_ (_04942_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _27402_ (_04943_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _27403_ (_04944_, _04943_, _04942_);
  and _27404_ (_04945_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _27405_ (_04946_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _27406_ (_04947_, _04946_, _04945_);
  and _27407_ (_04948_, _04947_, _04944_);
  and _27408_ (_04949_, _04948_, _04596_);
  and _27409_ (_04950_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _27410_ (_04951_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor _27411_ (_04952_, _04951_, _04950_);
  and _27412_ (_04953_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _27413_ (_04954_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _27414_ (_04955_, _04954_, _04953_);
  and _27415_ (_04956_, _04955_, _04952_);
  and _27416_ (_04957_, _04956_, _04565_);
  or _27417_ (_04958_, _04957_, _04570_);
  nor _27418_ (_04959_, _04958_, _04949_);
  and _27419_ (_04960_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _27420_ (_04961_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _27421_ (_04962_, _04961_, _04960_);
  and _27422_ (_04963_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _27423_ (_04964_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _27424_ (_04965_, _04964_, _04963_);
  and _27425_ (_04966_, _04965_, _04962_);
  nor _27426_ (_04967_, _04966_, _04565_);
  and _27427_ (_04968_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _27428_ (_04969_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _27429_ (_04970_, _04969_, _04968_);
  and _27430_ (_04971_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _27431_ (_04972_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _27432_ (_04973_, _04972_, _04971_);
  and _27433_ (_04974_, _04973_, _04970_);
  nor _27434_ (_04975_, _04974_, _04596_);
  or _27435_ (_04976_, _04975_, _04967_);
  and _27436_ (_04977_, _04976_, _04570_);
  nor _27437_ (_04978_, _04977_, _04959_);
  nor _27438_ (_04979_, _04978_, _04618_);
  and _27439_ (_04980_, _04979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27440_ (_04981_, _04940_, _01884_);
  nor _27441_ (_04982_, _04981_, _04941_);
  and _27442_ (_04983_, _04982_, _04980_);
  nor _27443_ (_04984_, _04983_, _04941_);
  nor _27444_ (_04985_, _04901_, _04863_);
  nor _27445_ (_04986_, _04985_, _04902_);
  not _27446_ (_04987_, _04986_);
  nor _27447_ (_04988_, _04987_, _04984_);
  nor _27448_ (_04989_, _04988_, _04902_);
  nor _27449_ (_04990_, _04989_, _04859_);
  nor _27450_ (_04991_, _04990_, _04858_);
  nor _27451_ (_04992_, _04816_, _04814_);
  nor _27452_ (_04993_, _04992_, _04817_);
  not _27453_ (_04994_, _04993_);
  nor _27454_ (_04995_, _04994_, _04991_);
  nor _27455_ (_04996_, _04995_, _04817_);
  nor _27456_ (_04997_, _04996_, _04776_);
  nor _27457_ (_04998_, _04997_, _04773_);
  nor _27458_ (_04999_, _04998_, _04732_);
  nor _27459_ (_05000_, _04999_, _04729_);
  nor _27460_ (_05001_, _05000_, _04688_);
  or _27461_ (_05002_, _05001_, _04687_);
  nor _27462_ (_05003_, _04681_, _04656_);
  nor _27463_ (_05004_, _05003_, _04682_);
  and _27464_ (_05005_, _05004_, _05002_);
  and _27465_ (_05006_, _05005_, _04684_);
  or _27466_ (_05007_, _05006_, _04682_);
  nor _27467_ (_05008_, _05007_, _04679_);
  nor _27468_ (_05009_, _05008_, _04676_);
  and _27469_ (_05010_, _05009_, _04673_);
  or _27470_ (_05011_, _05010_, _04671_);
  nor _27471_ (_05012_, _05011_, _04668_);
  nor _27472_ (_05013_, _04658_, _04656_);
  nor _27473_ (_05014_, _05013_, _04659_);
  not _27474_ (_05015_, _05014_);
  nor _27475_ (_05016_, _05015_, _05012_);
  and _27476_ (_05017_, _05016_, _04665_);
  or _27477_ (_05018_, _05017_, _04663_);
  nor _27478_ (_05019_, _05018_, _04660_);
  and _27479_ (_05020_, _05019_, _04561_);
  not _27480_ (_05021_, _05020_);
  not _27481_ (_05022_, _04656_);
  nor _27482_ (_05023_, _05019_, _05022_);
  nor _27483_ (_05024_, _04656_, _04561_);
  nor _27484_ (_05025_, _05024_, cy_reg);
  not _27485_ (_05026_, _05025_);
  nor _27486_ (_05027_, _05026_, _05023_);
  and _27487_ (_05028_, _05027_, _05021_);
  nor _27488_ (_05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _27489_ (_05030_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  or _27490_ (_05031_, _05030_, _05029_);
  nand _27491_ (_05032_, _05031_, _04559_);
  or _27492_ (_05033_, _05031_, _04559_);
  and _27493_ (_05034_, _05033_, _05032_);
  nor _27494_ (_05035_, _05034_, _05028_);
  not _27495_ (_05036_, cy_reg);
  nor _27496_ (_05037_, _04662_, _05036_);
  nor _27497_ (_05038_, _05016_, _04659_);
  nor _27498_ (_05039_, _05038_, _04665_);
  and _27499_ (_05040_, _05038_, _04665_);
  or _27500_ (_05041_, _05040_, _05039_);
  nor _27501_ (_05042_, _05041_, cy_reg);
  nor _27502_ (_05043_, _05042_, _05037_);
  nor _27503_ (_05044_, _05043_, _02178_);
  and _27504_ (_05045_, _05034_, _05028_);
  or _27505_ (_05046_, _05045_, _05044_);
  or _27506_ (_05047_, _05046_, _05035_);
  and _27507_ (_05048_, _04561_, cy_reg);
  and _27508_ (_05049_, _04656_, _04561_);
  nor _27509_ (_05050_, _05049_, _05024_);
  nor _27510_ (_05051_, _05050_, _05019_);
  and _27511_ (_05052_, _05050_, _05019_);
  or _27512_ (_05053_, _05052_, _05051_);
  and _27513_ (_05054_, _05053_, _05036_);
  nor _27514_ (_05055_, _05054_, _05048_);
  and _27515_ (_05056_, _05055_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _27516_ (_05057_, _05055_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _27517_ (_05058_, _05043_, _02178_);
  nor _27518_ (_05059_, _04667_, _05036_);
  nor _27519_ (_05060_, _05009_, _04671_);
  nor _27520_ (_05061_, _05060_, _04673_);
  and _27521_ (_05062_, _05060_, _04673_);
  or _27522_ (_05063_, _05062_, _05061_);
  nor _27523_ (_05064_, _05063_, cy_reg);
  nor _27524_ (_05065_, _05064_, _05059_);
  and _27525_ (_05066_, _05065_, _01872_);
  nor _27526_ (_05067_, _05065_, _01872_);
  and _27527_ (_05068_, _04678_, cy_reg);
  nor _27528_ (_05069_, _05005_, _04682_);
  and _27529_ (_05070_, _05069_, _04684_);
  nor _27530_ (_05071_, _05069_, _04684_);
  nor _27531_ (_05072_, _05071_, _05070_);
  nor _27532_ (_05073_, _05072_, cy_reg);
  nor _27533_ (_05074_, _05073_, _05068_);
  nor _27534_ (_05075_, _05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _27535_ (_05076_, _05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _27536_ (_05077_, _04686_, cy_reg);
  nor _27537_ (_05078_, _04687_, _04688_);
  and _27538_ (_05079_, _05078_, _05000_);
  nor _27539_ (_05080_, _05078_, _05000_);
  or _27540_ (_05081_, _05080_, _05079_);
  and _27541_ (_05082_, _05081_, _05036_);
  or _27542_ (_05083_, _05082_, _05077_);
  and _27543_ (_05084_, _05083_, _01996_);
  nor _27544_ (_05085_, _05083_, _01996_);
  and _27545_ (_05086_, _04998_, _04732_);
  nor _27546_ (_05087_, _05086_, _04999_);
  nor _27547_ (_05088_, _05087_, cy_reg);
  nor _27548_ (_05089_, _04728_, _05036_);
  nor _27549_ (_05090_, _05089_, _05088_);
  and _27550_ (_05091_, _05090_, _02437_);
  nor _27551_ (_05092_, _05090_, _02437_);
  and _27552_ (_05093_, _04996_, _04776_);
  nor _27553_ (_05094_, _05093_, _04997_);
  nor _27554_ (_05095_, _05094_, cy_reg);
  nor _27555_ (_05096_, _04772_, _05036_);
  nor _27556_ (_05097_, _05096_, _05095_);
  and _27557_ (_05098_, _05097_, _02076_);
  nor _27558_ (_05099_, _05097_, _02076_);
  and _27559_ (_05100_, _04816_, cy_reg);
  and _27560_ (_05101_, _04994_, _04991_);
  nor _27561_ (_05102_, _05101_, _04995_);
  and _27562_ (_05103_, _05102_, _05036_);
  nor _27563_ (_05104_, _05103_, _05100_);
  and _27564_ (_05105_, _05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _27565_ (_05106_, _04857_, cy_reg);
  nor _27566_ (_05107_, _04859_, _04858_);
  not _27567_ (_05108_, _05107_);
  nor _27568_ (_05109_, _05108_, _04989_);
  and _27569_ (_05110_, _05108_, _04989_);
  nor _27570_ (_05111_, _05110_, _05109_);
  and _27571_ (_05112_, _05111_, _05036_);
  nor _27572_ (_05113_, _05112_, _05106_);
  nor _27573_ (_05114_, _05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27574_ (_05115_, _05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27575_ (_05116_, _04862_, _05036_);
  and _27576_ (_05117_, _04987_, _04984_);
  nor _27577_ (_05118_, _05117_, _04988_);
  and _27578_ (_05119_, _05118_, _05036_);
  nor _27579_ (_05120_, _05119_, _05116_);
  nor _27580_ (_05121_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27581_ (_05122_, _04979_, _05036_);
  nor _27582_ (_05123_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27583_ (_05124_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27584_ (_05125_, _05124_, _05123_);
  nand _27585_ (_05126_, _05125_, _05122_);
  or _27586_ (_05127_, _05125_, _05122_);
  and _27587_ (_05128_, _05127_, _05126_);
  nor _27588_ (_05129_, _04982_, _04980_);
  nor _27589_ (_05130_, _05129_, _04983_);
  nor _27590_ (_05131_, _05130_, cy_reg);
  and _27591_ (_05132_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _27592_ (_05133_, _05132_, _05131_);
  and _27593_ (_05134_, _05133_, _02433_);
  nor _27594_ (_05135_, _05133_, _02433_);
  or _27595_ (_05136_, _05135_, _05134_);
  or _27596_ (_05137_, _05136_, _05128_);
  and _27597_ (_05138_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27598_ (_05139_, _05138_, _05137_);
  or _27599_ (_05140_, _05139_, _05121_);
  or _27600_ (_05141_, _05140_, _05115_);
  or _27601_ (_05142_, _05141_, _05114_);
  nor _27602_ (_05143_, _05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _27603_ (_05144_, _05143_, _05142_);
  or _27604_ (_05145_, _05144_, _05105_);
  or _27605_ (_05146_, _05145_, _05099_);
  or _27606_ (_05147_, _05146_, _05098_);
  or _27607_ (_05148_, _05147_, _05092_);
  or _27608_ (_05149_, _05148_, _05091_);
  or _27609_ (_05150_, _05149_, _05085_);
  or _27610_ (_05151_, _05150_, _05084_);
  nor _27611_ (_05152_, _05004_, _05002_);
  nor _27612_ (_05153_, _05152_, _05005_);
  nor _27613_ (_05154_, _05153_, cy_reg);
  nor _27614_ (_05155_, _04681_, _05036_);
  nor _27615_ (_05156_, _05155_, _05154_);
  nor _27616_ (_05157_, _05156_, _01876_);
  and _27617_ (_05158_, _05156_, _01876_);
  or _27618_ (_05159_, _05158_, _05157_);
  or _27619_ (_05160_, _05159_, _05151_);
  or _27620_ (_05161_, _05160_, _05076_);
  or _27621_ (_05162_, _05161_, _05075_);
  and _27622_ (_05163_, _04670_, cy_reg);
  and _27623_ (_05164_, _05008_, _04676_);
  nor _27624_ (_05165_, _05164_, _05009_);
  and _27625_ (_05166_, _05165_, _05036_);
  nor _27626_ (_05167_, _05166_, _05163_);
  and _27627_ (_05168_, _05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor _27628_ (_05169_, _05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or _27629_ (_05170_, _05169_, _05168_);
  or _27630_ (_05171_, _05170_, _05162_);
  or _27631_ (_05172_, _05171_, _05067_);
  or _27632_ (_05173_, _05172_, _05066_);
  and _27633_ (_05174_, _04658_, cy_reg);
  and _27634_ (_05175_, _05015_, _05012_);
  nor _27635_ (_05176_, _05175_, _05016_);
  and _27636_ (_05177_, _05176_, _05036_);
  nor _27637_ (_05178_, _05177_, _05174_);
  and _27638_ (_05179_, _05178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor _27639_ (_05180_, _05178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or _27640_ (_05181_, _05180_, _05179_);
  or _27641_ (_05182_, _05181_, _05173_);
  or _27642_ (_05183_, _05182_, _05058_);
  or _27643_ (_05184_, _05183_, _05057_);
  or _27644_ (_05185_, _05184_, _05056_);
  or _27645_ (_05186_, _05185_, _05047_);
  and _27646_ (_05187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27647_ (_05188_, _05187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _27648_ (_05189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27649_ (_05190_, _05189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _27650_ (_05191_, _05190_, _05188_);
  not _27651_ (_05192_, _05191_);
  nor _27652_ (_05193_, _05188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27653_ (_05194_, _05188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27654_ (_05195_, _05194_, _05193_);
  or _27655_ (_05196_, _05195_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand _27656_ (_05197_, _05195_, _08925_);
  and _27657_ (_05198_, _05197_, _05196_);
  and _27658_ (_05199_, _05198_, _05192_);
  or _27659_ (_05200_, _05195_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _27660_ (_05201_, _05195_, _08203_);
  and _27661_ (_05202_, _05201_, _05191_);
  and _27662_ (_05203_, _05202_, _05200_);
  or _27663_ (_05204_, _05203_, _05199_);
  or _27664_ (_05205_, _05204_, _02433_);
  or _27665_ (_05206_, _02000_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27666_ (_05207_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27667_ (_05208_, _05207_, _05187_);
  and _27668_ (_05209_, _05208_, _05206_);
  and _27669_ (_05210_, _02429_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27670_ (_05211_, _02000_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _27671_ (_05212_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [13]);
  or _27672_ (_05213_, _05212_, _05211_);
  and _27673_ (_05214_, _05213_, _05210_);
  or _27674_ (_05215_, _05214_, _05209_);
  nor _27675_ (_05216_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _27676_ (_05217_, _05216_, _02429_);
  nor _27677_ (_05218_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27678_ (_05219_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _27679_ (_05220_, _05219_, _05218_);
  and _27680_ (_05221_, _05220_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _27681_ (_05222_, _05216_, _02429_);
  nor _27682_ (_05223_, _05222_, _05217_);
  or _27683_ (_05224_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _08819_);
  nand _27684_ (_05225_, _05224_, _05223_);
  or _27685_ (_05226_, _05225_, _05221_);
  and _27686_ (_05227_, _05226_, _02433_);
  nor _27687_ (_05228_, _05220_, _08210_);
  and _27688_ (_05229_, _05220_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _27689_ (_05230_, _05229_, _05228_);
  or _27690_ (_05231_, _05230_, _05223_);
  and _27691_ (_05232_, _05231_, _05227_);
  or _27692_ (_05233_, _05232_, _05215_);
  and _27693_ (_05234_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _27694_ (_05235_, _02000_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _27695_ (_05236_, _05235_, _05234_);
  and _27696_ (_05237_, _05236_, _02429_);
  and _27697_ (_05238_, _02000_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _27698_ (_05239_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27699_ (_05240_, _05239_, _05238_);
  and _27700_ (_05241_, _05240_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27701_ (_05242_, _05241_, _05237_);
  or _27702_ (_05243_, _05242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27703_ (_05244_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and _27704_ (_05245_, _02000_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _27705_ (_05246_, _05245_, _02429_);
  or _27706_ (_05247_, _05246_, _05244_);
  or _27707_ (_05248_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27708_ (_05249_, _02000_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _27709_ (_05250_, _05249_, _05248_);
  or _27710_ (_05251_, _05250_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27711_ (_05252_, _05251_, _05247_);
  or _27712_ (_05253_, _05252_, _02433_);
  and _27713_ (_05254_, _05253_, _02004_);
  and _27714_ (_05255_, _05254_, _05243_);
  and _27715_ (_05256_, _05210_, _05240_);
  or _27716_ (_05257_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _27717_ (_05258_, _02000_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27718_ (_05259_, _05258_, _05187_);
  and _27719_ (_05260_, _05259_, _05257_);
  or _27720_ (_05261_, _05260_, _05256_);
  and _27721_ (_05262_, _05252_, _02433_);
  or _27722_ (_05263_, _05262_, _05261_);
  and _27723_ (_05264_, _05263_, _05255_);
  nor _27724_ (_05265_, _05195_, _08176_);
  and _27725_ (_05266_, _05195_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _27726_ (_05267_, _05266_, _05265_);
  and _27727_ (_05268_, _05267_, _05192_);
  or _27728_ (_05269_, _05195_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand _27729_ (_05270_, _05195_, _08215_);
  and _27730_ (_05271_, _05270_, _05191_);
  and _27731_ (_05272_, _05271_, _05269_);
  or _27732_ (_05273_, _05272_, _05268_);
  or _27733_ (_05274_, _05273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27734_ (_05275_, _05274_, _05264_);
  and _27735_ (_05276_, _05275_, _05233_);
  and _27736_ (_05277_, _05276_, _05205_);
  or _27737_ (_05278_, _02433_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _27738_ (_05279_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _27739_ (_05280_, _05279_, _05278_);
  nand _27740_ (_05281_, _05280_, _05220_);
  or _27741_ (_05282_, _02433_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _27742_ (_05283_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27743_ (_05284_, _05283_, _05282_);
  or _27744_ (_05285_, _05284_, _05220_);
  and _27745_ (_05286_, _05285_, _05281_);
  or _27746_ (_05287_, _05286_, _05223_);
  or _27747_ (_05288_, _05195_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand _27748_ (_05289_, _05195_, _08246_);
  and _27749_ (_05290_, _05289_, _05192_);
  and _27750_ (_05291_, _05290_, _05288_);
  nand _27751_ (_05292_, _05195_, _08233_);
  or _27752_ (_05293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _27753_ (_05294_, _05293_, _05191_);
  and _27754_ (_05295_, _05294_, _05292_);
  or _27755_ (_05296_, _05295_, _02433_);
  or _27756_ (_05297_, _05296_, _05291_);
  nand _27757_ (_05298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _27758_ (_05299_, _05298_, _05224_);
  and _27759_ (_05300_, _05299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _27760_ (_05301_, _02000_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _27761_ (_05302_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _27762_ (_05303_, _05302_, _02429_);
  and _27763_ (_05304_, _05303_, _05301_);
  or _27764_ (_05305_, _05304_, _05300_);
  and _27765_ (_05306_, _05305_, _05189_);
  and _27766_ (_05307_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02433_);
  or _27767_ (_05308_, _05213_, _02429_);
  or _27768_ (_05309_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _27769_ (_05310_, _02000_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _27770_ (_05311_, _05310_, _05309_);
  or _27771_ (_05312_, _05311_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27772_ (_05313_, _05312_, _05308_);
  and _27773_ (_05314_, _05313_, _05307_);
  or _27774_ (_05315_, _05314_, _05306_);
  and _27775_ (_05316_, _05305_, _02433_);
  or _27776_ (_05317_, _05316_, _05215_);
  and _27777_ (_05318_, _05317_, _05315_);
  and _27778_ (_05319_, _05318_, _05297_);
  and _27779_ (_05320_, _05319_, _05287_);
  nand _27780_ (_05321_, _05195_, _08228_);
  or _27781_ (_05322_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _27782_ (_05323_, _05322_, _05321_);
  or _27783_ (_05324_, _05323_, _05192_);
  or _27784_ (_05325_, _05195_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _27785_ (_05326_, _05195_, _08886_);
  and _27786_ (_05327_, _05326_, _05325_);
  or _27787_ (_05328_, _05327_, _05191_);
  and _27788_ (_05329_, _05328_, _05324_);
  or _27789_ (_05330_, _05329_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27790_ (_05331_, _05220_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _27791_ (_05332_, _05245_, _02433_);
  or _27792_ (_05333_, _05332_, _05331_);
  and _27793_ (_05334_, _05220_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _27794_ (_05335_, _05238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _27795_ (_05336_, _05335_, _05334_);
  nand _27796_ (_05337_, _05336_, _05333_);
  nand _27797_ (_05338_, _05337_, _05223_);
  and _27798_ (_05339_, _05338_, _05330_);
  and _27799_ (_05340_, _05339_, _05320_);
  or _27800_ (_05341_, _05340_, _05277_);
  nor _27801_ (_05342_, _04578_, _02461_);
  nor _27802_ (_05343_, _05342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27803_ (_05344_, _05342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27804_ (_05345_, _05344_, _05343_);
  nand _27805_ (_05346_, _05345_, _08233_);
  nor _27806_ (_05347_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27807_ (_05348_, _05347_, _02453_);
  nor _27808_ (_05349_, _05348_, _05342_);
  and _27809_ (_05350_, _05349_, _04602_);
  and _27810_ (_05351_, _05350_, _05346_);
  or _27811_ (_05352_, _05345_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not _27812_ (_05353_, _05349_);
  nand _27813_ (_05354_, _05345_, _08246_);
  and _27814_ (_05355_, _05354_, _05353_);
  and _27815_ (_05356_, _05355_, _05352_);
  or _27816_ (_05357_, _05356_, _05351_);
  and _27817_ (_05358_, _05357_, _04581_);
  nand _27818_ (_05359_, _05345_, _08215_);
  and _27819_ (_05360_, _05349_, _04607_);
  and _27820_ (_05361_, _05360_, _05359_);
  and _27821_ (_05362_, _05345_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _27822_ (_05363_, _05345_, _08176_);
  or _27823_ (_05364_, _05363_, _05362_);
  and _27824_ (_05365_, _05364_, _05353_);
  or _27825_ (_05366_, _05365_, _05361_);
  and _27826_ (_05367_, _05366_, _04566_);
  or _27827_ (_05368_, _05367_, _05358_);
  nand _27828_ (_05369_, _05345_, _08228_);
  and _27829_ (_05370_, _05349_, _04598_);
  and _27830_ (_05371_, _05370_, _05369_);
  and _27831_ (_05372_, _05345_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _27832_ (_05373_, _05345_, _08240_);
  or _27833_ (_05374_, _05373_, _05372_);
  and _27834_ (_05375_, _05374_, _05353_);
  or _27835_ (_05376_, _05375_, _05371_);
  and _27836_ (_05377_, _05376_, _04562_);
  nand _27837_ (_05378_, _05345_, _08203_);
  and _27838_ (_05379_, _05349_, _04611_);
  and _27839_ (_05380_, _05379_, _05378_);
  and _27840_ (_05381_, _05345_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _27841_ (_05382_, _05345_, _08210_);
  or _27842_ (_05383_, _05382_, _05381_);
  and _27843_ (_05384_, _05383_, _05353_);
  or _27844_ (_05385_, _05384_, _05380_);
  and _27845_ (_05386_, _05385_, _04578_);
  or _27846_ (_05387_, _05386_, _05377_);
  or _27847_ (_05388_, _05387_, _05368_);
  nor _27848_ (_05389_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _27849_ (_05390_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _27850_ (_05391_, _05390_, _05389_);
  or _27851_ (_05392_, _05391_, _04579_);
  nor _27852_ (_05393_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _27853_ (_05394_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand _27854_ (_05395_, _05394_, _05393_);
  nand _27855_ (_05396_, _05395_, _04562_);
  and _27856_ (_05397_, _05396_, _05392_);
  nor _27857_ (_05398_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _27858_ (_05399_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _27859_ (_05400_, _05399_, _05398_);
  nand _27860_ (_05401_, _05400_, _04566_);
  nor _27861_ (_05402_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _27862_ (_05403_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand _27863_ (_05404_, _05403_, _05402_);
  nand _27864_ (_05405_, _05404_, _04581_);
  and _27865_ (_05406_, _05405_, _05401_);
  and _27866_ (_05407_, _05406_, _05397_);
  nand _27867_ (_05408_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _27868_ (_05409_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _27869_ (_05410_, _05409_, _05408_);
  nand _27870_ (_05411_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand _27871_ (_05412_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _27872_ (_05413_, _05412_, _05411_);
  and _27873_ (_05414_, _05413_, _05410_);
  nand _27874_ (_05415_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _27875_ (_05416_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _27876_ (_05417_, _05416_, _05415_);
  nand _27877_ (_05418_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _27878_ (_05419_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _27879_ (_05420_, _05419_, _05418_);
  and _27880_ (_05421_, _05420_, _05417_);
  and _27881_ (_05422_, _05421_, _05414_);
  and _27882_ (_05423_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _27883_ (_05424_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or _27884_ (_05425_, _05424_, _05423_);
  and _27885_ (_05426_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _27886_ (_05427_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or _27887_ (_05428_, _05427_, _05426_);
  or _27888_ (_05429_, _05428_, _05425_);
  and _27889_ (_05430_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _27890_ (_05431_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _27891_ (_05432_, _05431_, _05430_);
  and _27892_ (_05433_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _27893_ (_05434_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _27894_ (_05435_, _05434_, _05433_);
  or _27895_ (_05436_, _05435_, _05432_);
  and _27896_ (_05437_, _05436_, _05429_);
  and _27897_ (_05438_, _05437_, _05422_);
  and _27898_ (_05439_, _05438_, _05407_);
  or _27899_ (_05440_, _05439_, _02461_);
  nor _27900_ (_05441_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _27901_ (_05442_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _27902_ (_05443_, _05442_, _05441_);
  or _27903_ (_05444_, _05443_, _04579_);
  or _27904_ (_05445_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand _27905_ (_05446_, _05445_, _04562_);
  or _27906_ (_05447_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand _27907_ (_05448_, _05447_, _04562_);
  and _27908_ (_05449_, _05448_, _05446_);
  and _27909_ (_05450_, _05449_, _05444_);
  nor _27910_ (_05451_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _27911_ (_05452_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _27912_ (_05453_, _05452_, _05451_);
  nand _27913_ (_05454_, _05453_, _04581_);
  nor _27914_ (_05455_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _27915_ (_05456_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _27916_ (_05457_, _05456_, _05455_);
  nand _27917_ (_05458_, _05457_, _04566_);
  and _27918_ (_05459_, _05458_, _05454_);
  and _27919_ (_05460_, _05459_, _05450_);
  nand _27920_ (_05461_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _27921_ (_05462_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _27922_ (_05463_, _05462_, _05461_);
  nand _27923_ (_05464_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _27924_ (_05465_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _27925_ (_05466_, _05465_, _05464_);
  and _27926_ (_05467_, _05466_, _05463_);
  nand _27927_ (_05468_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nand _27928_ (_05469_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _27929_ (_05470_, _05469_, _05468_);
  nand _27930_ (_05471_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nand _27931_ (_05472_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _27932_ (_05473_, _05472_, _05471_);
  and _27933_ (_05474_, _05473_, _05470_);
  and _27934_ (_05475_, _05474_, _05467_);
  and _27935_ (_05476_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _27936_ (_05477_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or _27937_ (_05478_, _05477_, _05476_);
  and _27938_ (_05479_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _27939_ (_05480_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or _27940_ (_05481_, _05480_, _05479_);
  or _27941_ (_05482_, _05481_, _05478_);
  and _27942_ (_05483_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _27943_ (_05484_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or _27944_ (_05485_, _05484_, _05483_);
  and _27945_ (_05486_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _27946_ (_05487_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or _27947_ (_05488_, _05487_, _05486_);
  or _27948_ (_05489_, _05488_, _05485_);
  and _27949_ (_05490_, _05489_, _05482_);
  and _27950_ (_05491_, _05490_, _05475_);
  and _27951_ (_05492_, _05491_, _05460_);
  or _27952_ (_05493_, _05492_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27953_ (_05494_, _05493_, _05440_);
  or _27954_ (_05495_, _05494_, _02457_);
  and _27955_ (_05496_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _27956_ (_05497_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or _27957_ (_05498_, _05497_, _05496_);
  and _27958_ (_05499_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _27959_ (_05500_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or _27960_ (_05501_, _05500_, _05499_);
  or _27961_ (_05502_, _05501_, _05498_);
  and _27962_ (_05503_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _27963_ (_05504_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _27964_ (_05505_, _05504_, _05503_);
  and _27965_ (_05506_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _27966_ (_05507_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or _27967_ (_05508_, _05507_, _05506_);
  or _27968_ (_05509_, _05508_, _05505_);
  or _27969_ (_05510_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _27970_ (_05511_, _05510_, _04578_);
  or _27971_ (_05512_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand _27972_ (_05513_, _05512_, _04562_);
  or _27973_ (_05514_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _27974_ (_05515_, _05514_, _04581_);
  and _27975_ (_05516_, _05515_, _05513_);
  and _27976_ (_05517_, _05516_, _05511_);
  and _27977_ (_05518_, _05517_, _05509_);
  and _27978_ (_05519_, _05518_, _05502_);
  or _27979_ (_05520_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand _27980_ (_05521_, _05520_, _04562_);
  and _27981_ (_05522_, _05521_, _02461_);
  nand _27982_ (_05523_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or _27983_ (_05524_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _27984_ (_05525_, _05524_, _04566_);
  and _27985_ (_05526_, _05525_, _05523_);
  nand _27986_ (_05527_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand _27987_ (_05528_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _27988_ (_05529_, _05528_, _05527_);
  and _27989_ (_05530_, _05529_, _05526_);
  and _27990_ (_05531_, _05530_, _05522_);
  nand _27991_ (_05532_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _27992_ (_05533_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _27993_ (_05534_, _05533_, _05532_);
  nand _27994_ (_05535_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _27995_ (_05536_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _27996_ (_05537_, _05536_, _05535_);
  and _27997_ (_05538_, _05537_, _05534_);
  nand _27998_ (_05539_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or _27999_ (_05540_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand _28000_ (_05541_, _05540_, _04566_);
  and _28001_ (_05542_, _05541_, _05539_);
  or _28002_ (_05543_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _28003_ (_05544_, _05543_, _04581_);
  or _28004_ (_05545_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand _28005_ (_05546_, _05545_, _04578_);
  and _28006_ (_05547_, _05546_, _05544_);
  and _28007_ (_05548_, _05547_, _05542_);
  and _28008_ (_05549_, _05548_, _05538_);
  and _28009_ (_05550_, _05549_, _05531_);
  and _28010_ (_05551_, _05550_, _05519_);
  and _28011_ (_05552_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _28012_ (_05553_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or _28013_ (_05554_, _05553_, _05552_);
  and _28014_ (_05555_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _28015_ (_05556_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _28016_ (_05557_, _05556_, _05555_);
  or _28017_ (_05558_, _05557_, _05554_);
  and _28018_ (_05559_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _28019_ (_05560_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or _28020_ (_05561_, _05560_, _05559_);
  and _28021_ (_05562_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _28022_ (_05563_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or _28023_ (_05564_, _05563_, _05562_);
  or _28024_ (_05565_, _05564_, _05561_);
  or _28025_ (_05566_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _28026_ (_05567_, _05566_, _04578_);
  or _28027_ (_05568_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand _28028_ (_05569_, _05568_, _04562_);
  or _28029_ (_05570_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _28030_ (_05571_, _05570_, _04581_);
  and _28031_ (_05572_, _05571_, _05569_);
  and _28032_ (_05573_, _05572_, _05567_);
  and _28033_ (_05574_, _05573_, _05565_);
  and _28034_ (_05575_, _05574_, _05558_);
  nand _28035_ (_05576_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _28036_ (_05577_, _05576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand _28037_ (_05578_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _28038_ (_05579_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _28039_ (_05580_, _05579_, _05578_);
  or _28040_ (_05581_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand _28041_ (_05582_, _05581_, _04562_);
  or _28042_ (_05583_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand _28043_ (_05584_, _05583_, _04581_);
  and _28044_ (_05585_, _05584_, _05582_);
  and _28045_ (_05586_, _05585_, _05580_);
  and _28046_ (_05587_, _05586_, _05577_);
  nand _28047_ (_05588_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nand _28048_ (_05589_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _28049_ (_05590_, _05589_, _05588_);
  nand _28050_ (_05591_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or _28051_ (_05592_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand _28052_ (_05593_, _05592_, _04578_);
  and _28053_ (_05594_, _05593_, _05591_);
  and _28054_ (_05595_, _05594_, _05590_);
  nand _28055_ (_05596_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or _28056_ (_05597_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand _28057_ (_05598_, _05597_, _04566_);
  and _28058_ (_05599_, _05598_, _05596_);
  nand _28059_ (_05600_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or _28060_ (_05601_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _28061_ (_05602_, _05601_, _04566_);
  and _28062_ (_05603_, _05602_, _05600_);
  and _28063_ (_05604_, _05603_, _05599_);
  and _28064_ (_05605_, _05604_, _05595_);
  and _28065_ (_05606_, _05605_, _05587_);
  and _28066_ (_05607_, _05606_, _05575_);
  or _28067_ (_05608_, _05607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28068_ (_05609_, _05608_, _05551_);
  or _28069_ (_05610_, _02457_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _28070_ (_05611_, _04611_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _28071_ (_05612_, _05611_, _05610_);
  or _28072_ (_05613_, _02457_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _28073_ (_05614_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _28074_ (_05615_, _05614_, _02461_);
  and _28075_ (_05616_, _05615_, _05613_);
  or _28076_ (_05617_, _05616_, _05612_);
  and _28077_ (_05618_, _05617_, _01884_);
  or _28078_ (_05619_, _02457_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _28079_ (_05620_, _05619_, _04607_);
  and _28080_ (_05621_, _05620_, _04860_);
  or _28081_ (_05622_, _02457_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _28082_ (_05623_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _28083_ (_05624_, _05623_, _04547_);
  and _28084_ (_05625_, _05624_, _05622_);
  or _28085_ (_05626_, _05625_, _05621_);
  or _28086_ (_05627_, _05626_, _05618_);
  and _28087_ (_05628_, _05627_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _28088_ (_05629_, _02457_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _28089_ (_05630_, _04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _28090_ (_05631_, _05630_, _05629_);
  or _28091_ (_05632_, _02457_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _28092_ (_05633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and _28093_ (_05634_, _05633_, _02461_);
  and _28094_ (_05635_, _05634_, _05632_);
  or _28095_ (_05636_, _05635_, _05631_);
  and _28096_ (_05637_, _05636_, _04578_);
  and _28097_ (_05638_, _04566_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _28098_ (_05639_, _02457_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _28099_ (_05640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _28100_ (_05641_, _05640_, _05639_);
  and _28101_ (_05642_, _05641_, _05638_);
  or _28102_ (_05643_, _02457_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _28103_ (_05644_, _05643_, _04602_);
  and _28104_ (_05645_, _04860_, _02453_);
  and _28105_ (_05646_, _05645_, _05644_);
  or _28106_ (_05647_, _05646_, _05642_);
  or _28107_ (_05648_, _05647_, _05637_);
  or _28108_ (_05649_, _05648_, _05628_);
  and _28109_ (_05650_, _05617_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _28110_ (_05651_, _05620_, _04861_);
  or _28111_ (_05652_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _28112_ (_05653_, _02457_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _28113_ (_05654_, _05653_, _05652_);
  and _28114_ (_05655_, _05654_, _05347_);
  or _28115_ (_05656_, _05655_, _02453_);
  or _28116_ (_05657_, _05656_, _05651_);
  or _28117_ (_05658_, _05657_, _05650_);
  and _28118_ (_05659_, _05636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _28119_ (_05660_, _05644_, _04861_);
  and _28120_ (_05661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _28121_ (_05662_, _02457_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _28122_ (_05663_, _05662_, _05661_);
  and _28123_ (_05664_, _05663_, _05347_);
  or _28124_ (_05665_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _28125_ (_05666_, _05665_, _05660_);
  or _28126_ (_05667_, _05666_, _05659_);
  nor _28127_ (_05668_, _02472_, first_instr);
  and _28128_ (_05669_, _05668_, _05667_);
  and _28129_ (_05670_, _05669_, _05658_);
  and _28130_ (_05671_, _05670_, _05649_);
  and _28131_ (_05672_, _05671_, _05609_);
  nand _28132_ (_05673_, _05672_, _05495_);
  nor _28133_ (_05674_, _05673_, _04618_);
  and _28134_ (_05675_, _05674_, _05388_);
  and _28135_ (_05676_, _05675_, _05341_);
  and _28136_ (property_invalid_jnc, _05676_, _05186_);
  or _28137_ (_05677_, pc_log_change_r, _05036_);
  nand _28138_ (_05678_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _28139_ (_00000_, _05678_, _05677_);
  and _28140_ (_05679_, _02472_, first_instr);
  or _28141_ (_00001_, _05679_, rst);
  dff _28142_ (cy_reg, _00000_, clk);
  dff _28143_ (pc_log_change_r, pc_log_change, clk);
  dff _28144_ (first_instr, _00001_, clk);
  dff _28145_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _10170_, clk);
  dff _28146_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _10174_, clk);
  dff _28147_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _10176_, clk);
  dff _28148_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _10180_, clk);
  dff _28149_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _10184_, clk);
  dff _28150_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _10187_, clk);
  dff _28151_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _10190_, clk);
  dff _28152_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _14025_, clk);
  dff _28153_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _10077_, clk);
  dff _28154_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _10081_, clk);
  dff _28155_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _10086_, clk);
  dff _28156_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _10091_, clk);
  dff _28157_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _10094_, clk);
  dff _28158_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _10099_, clk);
  dff _28159_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _10104_, clk);
  dff _28160_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _10106_, clk);
  dff _28161_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _14024_, clk);
  dff _28162_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _09985_, clk);
  dff _28163_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _09989_, clk);
  dff _28164_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _09994_, clk);
  dff _28165_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _09996_, clk);
  dff _28166_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _10001_, clk);
  dff _28167_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _10005_, clk);
  dff _28168_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _10009_, clk);
  dff _28169_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _09885_, clk);
  dff _28170_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _09889_, clk);
  dff _28171_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _09892_, clk);
  dff _28172_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _09895_, clk);
  dff _28173_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _09898_, clk);
  dff _28174_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _09902_, clk);
  dff _28175_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _09905_, clk);
  dff _28176_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _09907_, clk);
  dff _28177_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _14016_, clk);
  dff _28178_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _14017_, clk);
  dff _28179_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _14018_, clk);
  dff _28180_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _14019_, clk);
  dff _28181_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _14020_, clk);
  dff _28182_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _14021_, clk);
  dff _28183_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _14022_, clk);
  dff _28184_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _14023_, clk);
  dff _28185_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _14008_, clk);
  dff _28186_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _14009_, clk);
  dff _28187_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _14010_, clk);
  dff _28188_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _14011_, clk);
  dff _28189_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _14012_, clk);
  dff _28190_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _14013_, clk);
  dff _28191_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _14014_, clk);
  dff _28192_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _14015_, clk);
  dff _28193_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _14046_, clk);
  dff _28194_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _14047_, clk);
  dff _28195_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _14048_, clk);
  dff _28196_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _14049_, clk);
  dff _28197_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _14050_, clk);
  dff _28198_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _14051_, clk);
  dff _28199_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _14052_, clk);
  dff _28200_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _14053_, clk);
  dff _28201_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _09547_, clk);
  dff _28202_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _09551_, clk);
  dff _28203_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _14040_, clk);
  dff _28204_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _14041_, clk);
  dff _28205_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _14042_, clk);
  dff _28206_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _14043_, clk);
  dff _28207_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _14044_, clk);
  dff _28208_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _14045_, clk);
  dff _28209_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _14032_, clk);
  dff _28210_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _14033_, clk);
  dff _28211_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _14034_, clk);
  dff _28212_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _14035_, clk);
  dff _28213_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _14036_, clk);
  dff _28214_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _14037_, clk);
  dff _28215_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _14038_, clk);
  dff _28216_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _14039_, clk);
  dff _28217_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _09356_, clk);
  dff _28218_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _09360_, clk);
  dff _28219_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _09363_, clk);
  dff _28220_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _09366_, clk);
  dff _28221_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _09371_, clk);
  dff _28222_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _09373_, clk);
  dff _28223_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _09376_, clk);
  dff _28224_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _09379_, clk);
  dff _28225_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _09253_, clk);
  dff _28226_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _09257_, clk);
  dff _28227_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _09261_, clk);
  dff _28228_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _09266_, clk);
  dff _28229_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _09270_, clk);
  dff _28230_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _09274_, clk);
  dff _28231_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _09278_, clk);
  dff _28232_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _09281_, clk);
  dff _28233_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _08846_, clk);
  dff _28234_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _08850_, clk);
  dff _28235_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _08855_, clk);
  dff _28236_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _08860_, clk);
  dff _28237_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _08863_, clk);
  dff _28238_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _08868_, clk);
  dff _28239_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _08872_, clk);
  dff _28240_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _08875_, clk);
  dff _28241_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _08738_, clk);
  dff _28242_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _08743_, clk);
  dff _28243_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _08747_, clk);
  dff _28244_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _08751_, clk);
  dff _28245_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _08755_, clk);
  dff _28246_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _08759_, clk);
  dff _28247_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _08763_, clk);
  dff _28248_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _08766_, clk);
  dff _28249_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _14027_, clk);
  dff _28250_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _09055_, clk);
  dff _28251_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _09058_, clk);
  dff _28252_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _09060_, clk);
  dff _28253_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _09065_, clk);
  dff _28254_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _09069_, clk);
  dff _28255_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _09074_, clk);
  dff _28256_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _09077_, clk);
  dff _28257_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _08960_, clk);
  dff _28258_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _08965_, clk);
  dff _28259_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _08969_, clk);
  dff _28260_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _08972_, clk);
  dff _28261_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _08976_, clk);
  dff _28262_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _14026_, clk);
  dff _28263_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _08981_, clk);
  dff _28264_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _08983_, clk);
  dff _28265_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _09161_, clk);
  dff _28266_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _09164_, clk);
  dff _28267_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _14028_, clk);
  dff _28268_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _14029_, clk);
  dff _28269_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _14030_, clk);
  dff _28270_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _14031_, clk);
  dff _28271_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _09176_, clk);
  dff _28272_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _09179_, clk);
  dff _28273_ (\oc8051_symbolic_cxrom1.regvalid [0], _07408_, clk);
  dff _28274_ (\oc8051_symbolic_cxrom1.regvalid [1], _07436_, clk);
  dff _28275_ (\oc8051_symbolic_cxrom1.regvalid [2], _07476_, clk);
  dff _28276_ (\oc8051_symbolic_cxrom1.regvalid [3], _07529_, clk);
  dff _28277_ (\oc8051_symbolic_cxrom1.regvalid [4], _07582_, clk);
  dff _28278_ (\oc8051_symbolic_cxrom1.regvalid [5], _07640_, clk);
  dff _28279_ (\oc8051_symbolic_cxrom1.regvalid [6], _07708_, clk);
  dff _28280_ (\oc8051_symbolic_cxrom1.regvalid [7], _07780_, clk);
  dff _28281_ (\oc8051_symbolic_cxrom1.regvalid [8], _07842_, clk);
  dff _28282_ (\oc8051_symbolic_cxrom1.regvalid [9], _07921_, clk);
  dff _28283_ (\oc8051_symbolic_cxrom1.regvalid [10], _07995_, clk);
  dff _28284_ (\oc8051_symbolic_cxrom1.regvalid [11], _08055_, clk);
  dff _28285_ (\oc8051_symbolic_cxrom1.regvalid [12], _08149_, clk);
  dff _28286_ (\oc8051_symbolic_cxrom1.regvalid [13], _08265_, clk);
  dff _28287_ (\oc8051_symbolic_cxrom1.regvalid [14], _08385_, clk);
  dff _28288_ (\oc8051_symbolic_cxrom1.regvalid [15], _07359_, clk);
  dff _28289_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13520_, clk);
  dff _28290_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11175_, clk);
  dff _28291_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _01851_, clk);
  dff _28292_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _13787_, clk);
  dff _28293_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03880_, clk);
  dff _28294_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _03929_, clk);
  dff _28295_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04231_, clk);
  dff _28296_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _03897_, clk);
  dff _28297_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _00186_, clk);
  dff _28298_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03639_, clk);
  dff _28299_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03585_, clk);
  dff _28300_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03521_, clk);
  dff _28301_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03500_, clk);
  dff _28302_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03499_, clk);
  dff _28303_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _00014_, clk);
  dff _28304_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00359_, clk);
  dff _28305_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07052_, clk);
  dff _28306_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _01317_, clk);
  dff _28307_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _06617_, clk);
  dff _28308_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _06606_, clk);
  dff _28309_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _06604_, clk);
  dff _28310_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _06589_, clk);
  dff _28311_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03450_, clk);
  dff _28312_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _05682_, clk);
  dff _28313_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _01763_, clk);
  dff _28314_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _02490_, clk);
  dff _28315_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _03013_, clk);
  dff _28316_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _03347_, clk);
  dff _28317_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _05974_, clk);
  dff _28318_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _06092_, clk);
  dff _28319_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _06074_, clk);
  dff _28320_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _06060_, clk);
  dff _28321_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _07066_, clk);
  dff _28322_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _07069_, clk);
  dff _28323_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _07072_, clk);
  dff _28324_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _07074_, clk);
  dff _28325_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _07077_, clk);
  dff _28326_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _07080_, clk);
  dff _28327_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _07082_, clk);
  dff _28328_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06950_, clk);
  dff _28329_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _12290_, clk);
  dff _28330_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _12300_, clk);
  dff _28331_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12907_, clk);
  dff _28332_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _02980_, clk);
  dff _28333_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04070_, clk);
  dff _28334_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _02983_, clk);
  dff _28335_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _07649_, clk);
  dff _28336_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04122_, clk);
  dff _28337_ (\oc8051_top_1.oc8051_decoder1.state [0], _00393_, clk);
  dff _28338_ (\oc8051_top_1.oc8051_decoder1.state [1], _04056_, clk);
  dff _28339_ (\oc8051_top_1.oc8051_decoder1.op [0], _07568_, clk);
  dff _28340_ (\oc8051_top_1.oc8051_decoder1.op [1], _07382_, clk);
  dff _28341_ (\oc8051_top_1.oc8051_decoder1.op [2], _03936_, clk);
  dff _28342_ (\oc8051_top_1.oc8051_decoder1.op [3], _03756_, clk);
  dff _28343_ (\oc8051_top_1.oc8051_decoder1.op [4], _07485_, clk);
  dff _28344_ (\oc8051_top_1.oc8051_decoder1.op [5], _03702_, clk);
  dff _28345_ (\oc8051_top_1.oc8051_decoder1.op [6], _03565_, clk);
  dff _28346_ (\oc8051_top_1.oc8051_decoder1.op [7], _04144_, clk);
  dff _28347_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04146_, clk);
  dff _28348_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _11599_, clk);
  dff _28349_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04154_, clk);
  dff _28350_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _11499_, clk);
  dff _28351_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04157_, clk);
  dff _28352_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03742_, clk);
  dff _28353_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _11988_, clk);
  dff _28354_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04159_, clk);
  dff _28355_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _04111_, clk);
  dff _28356_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _04077_, clk);
  dff _28357_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04164_, clk);
  dff _28358_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03682_, clk);
  dff _28359_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04166_, clk);
  dff _28360_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03834_, clk);
  dff _28361_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _04065_, clk);
  dff _28362_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _04218_, clk);
  dff _28363_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04168_, clk);
  dff _28364_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03822_, clk);
  dff _28365_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04197_, clk);
  dff _28366_ (\oc8051_top_1.oc8051_decoder1.wr , _04201_, clk);
  dff _28367_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _00388_, clk);
  dff _28368_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _00872_, clk);
  dff _28369_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _03330_, clk);
  dff _28370_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _08716_, clk);
  dff _28371_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _06658_, clk);
  dff _28372_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _02255_, clk);
  dff _28373_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03813_, clk);
  dff _28374_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _01442_, clk);
  dff _28375_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _03847_, clk);
  dff _28376_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _02041_, clk);
  dff _28377_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _03317_, clk);
  dff _28378_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _05935_, clk);
  dff _28379_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _02074_, clk);
  dff _28380_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _11489_, clk);
  dff _28381_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _07111_, clk);
  dff _28382_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _03377_, clk);
  dff _28383_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _03924_, clk);
  dff _28384_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _02499_, clk);
  dff _28385_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _13801_, clk);
  dff _28386_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _12048_, clk);
  dff _28387_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00781_, clk);
  dff _28388_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _06811_, clk);
  dff _28389_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _02186_, clk);
  dff _28390_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12624_, clk);
  dff _28391_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _00826_, clk);
  dff _28392_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _13436_, clk);
  dff _28393_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _01189_, clk);
  dff _28394_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _01236_, clk);
  dff _28395_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _07982_, clk);
  dff _28396_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _01914_, clk);
  dff _28397_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _11544_, clk);
  dff _28398_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _09983_, clk);
  dff _28399_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02175_, clk);
  dff _28400_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _06778_, clk);
  dff _28401_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _01902_, clk);
  dff _28402_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _12997_, clk);
  dff _28403_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _03837_, clk);
  dff _28404_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _03823_, clk);
  dff _28405_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _03968_, clk);
  dff _28406_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _11892_, clk);
  dff _28407_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _10178_, clk);
  dff _28408_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _13487_, clk);
  dff _28409_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _12018_, clk);
  dff _28410_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _13371_, clk);
  dff _28411_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _13605_, clk);
  dff _28412_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _11820_, clk);
  dff _28413_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _12012_, clk);
  dff _28414_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _13686_, clk);
  dff _28415_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _09300_, clk);
  dff _28416_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _11767_, clk);
  dff _28417_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _12099_, clk);
  dff _28418_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _03576_, clk);
  dff _28419_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _12101_, clk);
  dff _28420_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _05750_, clk);
  dff _28421_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _08866_, clk);
  dff _28422_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _08890_, clk);
  dff _28423_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _03344_, clk);
  dff _28424_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _09087_, clk);
  dff _28425_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _11072_, clk);
  dff _28426_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _08870_, clk);
  dff _28427_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _08894_, clk);
  dff _28428_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _09193_, clk);
  dff _28429_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _00264_, clk);
  dff _28430_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _01835_, clk);
  dff _28431_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _12917_, clk);
  dff _28432_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _12170_, clk);
  dff _28433_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _11443_, clk);
  dff _28434_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _00531_, clk);
  dff _28435_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _00864_, clk);
  dff _28436_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _08157_, clk);
  dff _28437_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01059_, clk);
  dff _28438_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01648_, clk);
  dff _28439_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01642_, clk);
  dff _28440_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _01056_, clk);
  dff _28441_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _01152_, clk);
  dff _28442_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01658_, clk);
  dff _28443_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _01651_, clk);
  dff _28444_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _01052_, clk);
  dff _28445_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _01673_, clk);
  dff _28446_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _01663_, clk);
  dff _28447_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _01045_, clk);
  dff _28448_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _01145_, clk);
  dff _28449_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01180_, clk);
  dff _28450_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01202_, clk);
  dff _28451_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01679_, clk);
  dff _28452_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _00725_, clk);
  dff _28453_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01716_, clk);
  dff _28454_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01009_, clk);
  dff _28455_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _01730_, clk);
  dff _28456_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01719_, clk);
  dff _28457_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01006_, clk);
  dff _28458_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _01138_, clk);
  dff _28459_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _01734_, clk);
  dff _28460_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _01732_, clk);
  dff _28461_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _01002_, clk);
  dff _28462_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _01743_, clk);
  dff _28463_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _01736_, clk);
  dff _28464_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _00999_, clk);
  dff _28465_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _01135_, clk);
  dff _28466_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _01175_, clk);
  dff _28467_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _01199_, clk);
  dff _28468_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _04371_, clk);
  dff _28469_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04184_, clk);
  dff _28470_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04006_, clk);
  dff _28471_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _03907_, clk);
  dff _28472_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03488_, clk);
  dff _28473_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _03431_, clk);
  dff _28474_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _12214_, clk);
  dff _28475_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11440_, clk);
  dff _28476_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11720_, clk);
  dff _28477_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _11898_, clk);
  dff _28478_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _01247_, clk);
  dff _28479_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _07987_, clk);
  dff _28480_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _13610_, clk);
  dff _28481_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _11809_, clk);
  dff _28482_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _11494_, clk);
  dff _28483_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _11285_, clk);
  dff _28484_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _12254_, clk);
  dff _28485_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03889_, clk);
  dff _28486_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _12217_, clk);
  dff _28487_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _10032_, clk);
  dff _28488_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _08447_, clk);
  dff _28489_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _04050_, clk);
  dff _28490_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04040_, clk);
  dff _28491_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _12229_, clk);
  dff _28492_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _11437_, clk);
  dff _28493_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05684_, clk);
  dff _28494_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _02080_, clk);
  dff _28495_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _04094_, clk);
  dff _28496_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _12261_, clk);
  dff _28497_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05683_, clk);
  dff _28498_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00572_, clk);
  dff _28499_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05681_, clk);
  dff _28500_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03472_, clk);
  dff _28501_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _13941_, clk);
  dff _28502_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _12281_, clk);
  dff _28503_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _11432_, clk);
  dff _28504_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03678_, clk);
  dff _28505_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03669_, clk);
  dff _28506_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03652_, clk);
  dff _28507_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03645_, clk);
  dff _28508_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _12287_, clk);
  dff _28509_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03481_, clk);
  dff _28510_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03136_, clk);
  dff _28511_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _02688_, clk);
  dff _28512_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00574_, clk);
  dff _28513_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _01299_, clk);
  dff _28514_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _13110_, clk);
  dff _28515_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _13098_, clk);
  dff _28516_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _13085_, clk);
  dff _28517_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _13056_, clk);
  dff _28518_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _13034_, clk);
  dff _28519_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12334_, clk);
  dff _28520_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _13281_, clk);
  dff _28521_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _13359_, clk);
  dff _28522_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _13328_, clk);
  dff _28523_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _13289_, clk);
  dff _28524_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12327_, clk);
  dff _28525_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _11409_, clk);
  dff _28526_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _12526_, clk);
  dff _28527_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _12496_, clk);
  dff _28528_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _12490_, clk);
  dff _28529_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _02545_, clk);
  dff _28530_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _11941_, clk);
  dff _28531_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _11832_, clk);
  dff _28532_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _12345_, clk);
  dff _28533_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _12293_, clk);
  dff _28534_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _12089_, clk);
  dff _28535_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _12220_, clk);
  dff _28536_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _12175_, clk);
  dff _28537_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _12141_, clk);
  dff _28538_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _12111_, clk);
  dff _28539_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _12342_, clk);
  dff _28540_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11402_, clk);
  dff _28541_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11291_, clk);
  dff _28542_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _11181_, clk);
  dff _28543_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _11223_, clk);
  dff _28544_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _11220_, clk);
  dff _28545_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03479_, clk);
  dff _28546_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _11502_, clk);
  dff _28547_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _02025_, clk);
  dff _28548_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _04199_, clk);
  dff _28549_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _10459_, clk);
  dff _28550_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _10449_, clk);
  dff _28551_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10430_, clk);
  dff _28552_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12361_, clk);
  dff _28553_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _11034_, clk);
  dff _28554_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _10901_, clk);
  dff _28555_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _11033_, clk);
  dff _28556_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05942_, clk);
  dff _28557_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _12358_, clk);
  dff _28558_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11393_, clk);
  dff _28559_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03485_, clk);
  dff _28560_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _11712_, clk);
  dff _28561_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _11389_, clk);
  dff _28562_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _11692_, clk);
  dff _28563_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _11871_, clk);
  dff _28564_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _09186_, clk);
  dff _28565_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _01829_, clk);
  dff _28566_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _02239_, clk);
  dff _28567_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _12367_, clk);
  dff _28568_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _11373_, clk);
  dff _28569_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _01278_, clk);
  dff _28570_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _00563_, clk);
  dff _28571_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _12179_, clk);
  dff _28572_ (\oc8051_top_1.oc8051_memory_interface1.reti , _02547_, clk);
  dff _28573_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11677_, clk);
  dff _28574_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _06953_, clk);
  dff _28575_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00728_, clk);
  dff _28576_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00592_, clk);
  dff _28577_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _07131_, clk);
  dff _28578_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12392_, clk);
  dff _28579_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _03853_, clk);
  dff _28580_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03752_, clk);
  dff _28581_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _03772_, clk);
  dff _28582_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10975_, clk);
  dff _28583_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _07589_, clk);
  dff _28584_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _07524_, clk);
  dff _28585_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _07125_, clk);
  dff _28586_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03483_, clk);
  dff _28587_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _02874_, clk);
  dff _28588_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _02792_, clk);
  dff _28589_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _02908_, clk);
  dff _28590_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _02895_, clk);
  dff _28591_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11004_, clk);
  dff _28592_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _03353_, clk);
  dff _28593_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _03351_, clk);
  dff _28594_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _10999_, clk);
  dff _28595_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _03358_, clk);
  dff _28596_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _03356_, clk);
  dff _28597_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _10996_, clk);
  dff _28598_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11205_, clk);
  dff _28599_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11306_, clk);
  dff _28600_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11339_, clk);
  dff _28601_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _03440_, clk);
  dff _28602_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _03424_, clk);
  dff _28603_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _10993_, clk);
  dff _28604_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _03579_, clk);
  dff _28605_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _03563_, clk);
  dff _28606_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _10991_, clk);
  dff _28607_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11188_, clk);
  dff _28608_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _03630_, clk);
  dff _28609_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _03587_, clk);
  dff _28610_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _10986_, clk);
  dff _28611_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _03713_, clk);
  dff _28612_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _03650_, clk);
  dff _28613_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _10983_, clk);
  dff _28614_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11184_, clk);
  dff _28615_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11303_, clk);
  dff _28616_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _03748_, clk);
  dff _28617_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _03715_, clk);
  dff _28618_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _01816_, clk);
  dff _28619_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _02261_, clk);
  dff _28620_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _02149_, clk);
  dff _28621_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _02274_, clk);
  dff _28622_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11886_, clk);
  dff _28623_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _10909_, clk);
  dff _28624_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11159_, clk);
  dff _28625_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _12694_, clk);
  dff _28626_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _02427_, clk);
  dff _28627_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _28628_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _28629_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _28630_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _28631_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _28632_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _28633_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _28634_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _28635_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _28636_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _28637_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _28638_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _28639_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _28640_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _28641_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _28642_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _28643_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _28644_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _28645_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _28646_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _28647_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _28648_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _28649_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _28650_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _28651_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _28652_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _28653_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _28654_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _28655_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _28656_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _28657_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _28658_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _28659_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _04089_, clk);
  dff _28660_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _12448_, clk);
  dff _28661_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _12440_, clk);
  dff _28662_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12415_, clk);
  dff _28663_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04194_, clk);
  dff _28664_ (\oc8051_top_1.oc8051_sfr1.bit_out , _04186_, clk);
  dff _28665_ (\oc8051_top_1.oc8051_sfr1.wait_data , _04086_, clk);
  dff _28666_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _12265_, clk);
  dff _28667_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _12235_, clk);
  dff _28668_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _12232_, clk);
  dff _28669_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _12226_, clk);
  dff _28670_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03740_, clk);
  dff _28671_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03570_, clk);
  dff _28672_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03614_, clk);
  dff _28673_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04114_, clk);
  dff _28674_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08089_, clk);
  dff _28675_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _02537_, clk);
  dff _28676_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03891_, clk);
  dff _28677_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _04107_, clk);
  dff _28678_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _04054_, clk);
  dff _28679_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08085_, clk);
  dff _28680_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _07736_, clk);
  dff _28681_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _06199_, clk);
  dff _28682_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _00897_, clk);
  dff _28683_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00886_, clk);
  dff _28684_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _03554_, clk);
  dff _28685_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _00621_, clk);
  dff _28686_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00618_, clk);
  dff _28687_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _03592_, clk);
  dff _28688_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _00641_, clk);
  dff _28689_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03903_, clk);
  dff _28690_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07258_, clk);
  dff _28691_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07260_, clk);
  dff _28692_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _06049_, clk);
  dff _28693_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _02104_, clk);
  dff _28694_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _06063_, clk);
  dff _28695_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _06052_, clk);
  dff _28696_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _06034_, clk);
  dff _28697_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13246_, clk);
  dff _28698_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07234_, clk);
  dff _28699_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07238_, clk);
  dff _28700_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _06096_, clk);
  dff _28701_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _02094_, clk);
  dff _28702_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _04249_, clk);
  dff _28703_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _06130_, clk);
  dff _28704_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _02099_, clk);
  dff _28705_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13206_, clk);
  dff _28706_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _09235_, clk);
  dff _28707_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _01461_, clk);
  dff _28708_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _13581_, clk);
  dff _28709_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _13565_, clk);
  dff _28710_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _13573_, clk);
  dff _28711_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _13568_, clk);
  dff _28712_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _02794_, clk);
  dff _28713_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _13601_, clk);
  dff _28714_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _13596_, clk);
  dff _28715_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _02506_, clk);
  dff _28716_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _13517_, clk);
  dff _28717_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _01890_, clk);
  dff _28718_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _00503_, clk);
  dff _28719_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _13536_, clk);
  dff _28720_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _13542_, clk);
  dff _28721_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _00316_, clk);
  dff _28722_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _13478_, clk);
  dff _28723_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _13475_, clk);
  dff _28724_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13324_, clk);
  dff _28725_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _02813_, clk);
  dff _28726_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _02810_, clk);
  dff _28727_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _00433_, clk);
  dff _28728_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _00430_, clk);
  dff _28729_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08858_, clk);
  dff _28730_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _00475_, clk);
  dff _28731_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _13441_, clk);
  dff _28732_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _02825_, clk);
  dff _28733_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02549_, clk);
  dff _28734_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10482_, clk);
  dff _28735_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _13841_, clk);
  dff _28736_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _13834_, clk);
  dff _28737_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _02737_, clk);
  dff _28738_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _13868_, clk);
  dff _28739_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _13862_, clk);
  dff _28740_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _13859_, clk);
  dff _28741_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _13855_, clk);
  dff _28742_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10480_, clk);
  dff _28743_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _02741_, clk);
  dff _28744_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _02551_, clk);
  dff _28745_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _13775_, clk);
  dff _28746_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _13773_, clk);
  dff _28747_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _13768_, clk);
  dff _28748_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _02752_, clk);
  dff _28749_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _13795_, clk);
  dff _28750_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _00470_, clk);
  dff _28751_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _03285_, clk);
  dff _28752_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _03159_, clk);
  dff _28753_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03127_, clk);
  dff _28754_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _03289_, clk);
  dff _28755_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03162_, clk);
  dff _28756_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _03287_, clk);
  dff _28757_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03157_, clk);
  dff _28758_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _05680_, clk);
  dff _28759_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _03153_, clk);
  dff _28760_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03124_, clk);
  dff _28761_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _03296_, clk);
  dff _28762_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03155_, clk);
  dff _28763_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03294_, clk);
  dff _28764_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03151_, clk);
  dff _28765_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _03122_, clk);
  dff _28766_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _03745_, clk);
  dff _28767_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03291_, clk);
  dff _28768_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _03261_, clk);
  dff _28769_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03246_, clk);
  dff _28770_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03245_, clk);
  dff _28771_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03148_, clk);
  dff _28772_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _03119_, clk);
  dff _28773_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03300_, clk);
  dff _28774_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _03862_, clk);
  dff _28775_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _03298_, clk);
  dff _28776_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _03264_, clk);
  dff _28777_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03263_, clk);
  dff _28778_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _03305_, clk);
  dff _28779_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03146_, clk);
  dff _28780_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _03303_, clk);
  dff _28781_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03270_, clk);
  dff _28782_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03867_, clk);
  dff _28783_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _08610_, clk);
  dff _28784_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03322_, clk);
  dff _28785_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10419_, clk);
  dff _28786_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10433_, clk);
  dff _28787_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10427_, clk);
  dff _28788_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10424_, clk);
  dff _28789_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _04355_, clk);
  dff _28790_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03617_, clk);
  dff _28791_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _03671_, clk);
  dff _28792_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _14001_, clk);
  dff _28793_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _13965_, clk);
  dff _28794_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _13995_, clk);
  dff _28795_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _13992_, clk);
  dff _28796_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _13989_, clk);
  dff _28797_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _13984_, clk);
  dff _28798_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _00321_, clk);
  dff _28799_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01067_, clk);
  dff _28800_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01078_, clk);
  dff _28801_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _13388_, clk);
  dff _28802_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _13392_, clk);
  dff _28803_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _13369_, clk);
  dff _28804_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _13366_, clk);
  dff _28805_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _13363_, clk);
  dff _28806_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _13374_, clk);
  dff _28807_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _13336_, clk);
  dff _28808_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01071_, clk);
  dff _28809_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _13413_, clk);
  dff _28810_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13416_, clk);
  dff _28811_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _13433_, clk);
  dff _28812_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13424_, clk);
  dff _28813_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13430_, clk);
  dff _28814_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13427_, clk);
  dff _28815_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13497_, clk);
  dff _28816_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _01075_, clk);
  dff _28817_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _01073_, clk);
  dff _28818_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _01024_, clk);
  dff _28819_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13439_, clk);
  dff _28820_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13457_, clk);
  dff _28821_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13464_, clk);
  dff _28822_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13461_, clk);
  dff _28823_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13508_, clk);
  dff _28824_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13502_, clk);
  dff _28825_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13505_, clk);
  dff _28826_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _01028_, clk);
  dff _28827_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13591_, clk);
  dff _28828_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13561_, clk);
  dff _28829_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13563_, clk);
  dff _28830_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13571_, clk);
  dff _28831_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13575_, clk);
  dff _28832_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13548_, clk);
  dff _28833_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13545_, clk);
  dff _28834_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01026_, clk);
  dff _28835_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _01049_, clk);
  dff _28836_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13600_, clk);
  dff _28837_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13615_, clk);
  dff _28838_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13607_, clk);
  dff _28839_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13612_, clk);
  dff _28840_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13626_, clk);
  dff _28841_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13622_, clk);
  dff _28842_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13624_, clk);
  dff _28843_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _01039_, clk);
  dff _28844_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01705_, clk);
  dff _28845_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08853_, clk);
  dff _28846_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _04082_, clk);
  dff _28847_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _00258_, clk);
  dff _28848_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _01624_, clk);
  dff _28849_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01620_, clk);
  dff _28850_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _01618_, clk);
  dff _28851_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _01616_, clk);
  dff _28852_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _01580_, clk);
  dff _28853_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _01575_, clk);
  dff _28854_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _01572_, clk);
  dff _28855_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _03919_, clk);
  dff _28856_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _01520_, clk);
  dff _28857_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _01501_, clk);
  dff _28858_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _01517_, clk);
  dff _28859_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _01515_, clk);
  dff _28860_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01512_, clk);
  dff _28861_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _01505_, clk);
  dff _28862_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _01464_, clk);
  dff _28863_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _03780_, clk);
  dff _28864_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _04437_, clk);
  dff _28865_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01367_, clk);
  dff _28866_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _01328_, clk);
  dff _28867_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _01359_, clk);
  dff _28868_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _01348_, clk);
  dff _28869_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _01292_, clk);
  dff _28870_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _01275_, clk);
  dff _28871_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _01289_, clk);
  dff _28872_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01739_, clk);
  dff _28873_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _01224_, clk);
  dff _28874_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _01196_, clk);
  dff _28875_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _01191_, clk);
  dff _28876_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01162_, clk);
  dff _28877_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _01157_, clk);
  dff _28878_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _01154_, clk);
  dff _28879_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _01149_, clk);
  dff _28880_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01048_, clk);
  dff _28881_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _05877_, clk);
  dff _28882_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _01086_, clk);
  dff _28883_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _01083_, clk);
  dff _28884_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _01042_, clk);
  dff _28885_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _01036_, clk);
  dff _28886_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _01019_, clk);
  dff _28887_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _01015_, clk);
  dff _28888_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _01013_, clk);
  dff _28889_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _02561_, clk);
  dff _28890_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _07629_, clk);
  dff _28891_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07620_, clk);
  dff _28892_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07539_, clk);
  dff _28893_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07472_, clk);
  dff _28894_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07522_, clk);
  dff _28895_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07513_, clk);
  dff _28896_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07510_, clk);
  dff _28897_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07482_, clk);
  dff _28898_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _06783_, clk);
  dff _28899_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _06379_, clk);
  dff _28900_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _06679_, clk);
  dff _28901_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02754_, clk);
  dff _28902_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _06346_, clk);
  dff _28903_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _12554_, clk);
  dff _28904_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12396_, clk);
  dff _28905_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _01408_, clk);
  dff _28906_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _08216_, clk);
  dff _28907_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02559_, clk);
  dff _28908_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _08226_, clk);
  dff _28909_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _03444_, clk);
  dff _28910_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01870_, clk);
  dff _28911_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _09148_, clk);
  dff _28912_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _10877_, clk);
  dff _28913_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01306_, clk);
  dff _28914_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01756_, clk);
  dff _28915_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _03725_, clk);
  dff _28916_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _02197_, clk);
  dff _28917_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _02466_, clk);
  dff _28918_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02555_, clk);
  dff _28919_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _06909_, clk);
  dff _28920_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _02765_, clk);
  dff _28921_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02674_, clk);
  dff _28922_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02769_, clk);
  dff _28923_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02673_, clk);
  dff _28924_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02707_, clk);
  dff _28925_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _03057_, clk);
  dff _28926_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _12211_, clk);
  dff _28927_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _12373_, clk);
  dff _28928_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02782_, clk);
  dff _28929_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _12206_, clk);
  dff _28930_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04462_, clk);
  dff _28931_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04464_, clk);
  dff _28932_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _12203_, clk);
  dff _28933_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _12331_, clk);
  dff _28934_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _12471_, clk);
  dff _28935_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _12560_, clk);
  dff _28936_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04361_, clk);
  dff _28937_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04368_, clk);
  dff _28938_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _12200_, clk);
  dff _28939_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02780_, clk);
  dff _28940_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _04373_, clk);
  dff _28941_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _12193_, clk);
  dff _28942_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _12315_, clk);
  dff _28943_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12468_, clk);
  dff _28944_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _04480_, clk);
  dff _28945_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _04477_, clk);
  dff _28946_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _12190_, clk);
  dff _28947_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02665_, clk);
  dff _28948_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _12181_, clk);
  dff _28949_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12303_, clk);
  dff _28950_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12461_, clk);
  dff _28951_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12557_, clk);
  dff _28952_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _12600_, clk);
  dff _28953_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _02398_, clk);
  dff _28954_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _02400_, clk);
  dff _28955_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02786_, clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
