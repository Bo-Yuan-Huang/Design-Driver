
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jnc, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jnc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_05685_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_05686_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_05687_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor (_05688_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_05689_, _05688_, _05687_);
  and (_05690_, _05689_, _05686_);
  and (_05691_, _05690_, _05685_);
  nor (_05692_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05693_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_05694_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_05695_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_05696_, _05695_, _05694_);
  or (_05697_, _05696_, _05693_);
  not (_05698_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_05699_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05698_);
  nand (_05700_, _05699_, _05694_);
  not (_05701_, _05700_);
  nand (_05702_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_05703_, _05702_, _05697_);
  nand (_05704_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_05705_, _05704_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_05706_, _05705_);
  nand (_05707_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not (_05708_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  not (_05709_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_05710_, _05694_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nand (_05711_, _05710_, _05709_);
  or (_05712_, _05711_, _05708_);
  and (_05713_, _05712_, _05707_);
  and (_05714_, _05695_, _05694_);
  nand (_05715_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_05716_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_05717_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  or (_05718_, _05717_, _05694_);
  or (_05719_, _05718_, _05716_);
  and (_05720_, _05719_, _05715_);
  and (_05721_, _05720_, _05713_);
  nand (_05722_, _05721_, _05703_);
  nand (_05723_, _05722_, _05692_);
  and (_05724_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05725_, _05724_);
  nand (_05726_, _05725_, _05723_);
  not (_05727_, _05726_);
  or (_05728_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.cdone );
  nand (_05729_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_05730_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_05731_, _05730_, _05729_);
  not (_05732_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_05733_, _05711_, _05732_);
  not (_05734_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_05735_, _05700_, _05734_);
  and (_05736_, _05735_, _05733_);
  not (_05737_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_05738_, _05696_, _05737_);
  not (_05739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_05740_, _05718_, _05739_);
  and (_05741_, _05740_, _05738_);
  and (_05742_, _05741_, _05736_);
  and (_05743_, _05742_, _05731_);
  or (_05744_, _05743_, _05728_);
  and (_05745_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05746_, _05745_);
  nand (_05747_, _05746_, _05744_);
  not (_05748_, _05747_);
  not (_05749_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_05751_, _05696_, _05749_);
  nand (_05752_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_05753_, _05752_, _05751_);
  not (_05754_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_05755_, _05705_, _05754_);
  not (_05756_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_05757_, _05711_, _05756_);
  and (_05758_, _05757_, _05755_);
  nand (_05759_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not (_05760_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_05761_, _05718_, _05760_);
  and (_05762_, _05761_, _05759_);
  and (_05763_, _05762_, _05758_);
  and (_05764_, _05763_, _05753_);
  or (_05765_, _05764_, _05728_);
  and (_05766_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05767_, _05766_);
  nand (_05768_, _05767_, _05765_);
  and (_05769_, _05768_, _05748_);
  and (_05770_, _05769_, _05727_);
  and (_05771_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05772_, _05771_);
  not (_05773_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_05774_, _05718_, _05773_);
  nand (_05775_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_05776_, _05775_, _05774_);
  nand (_05777_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not (_05778_, _05711_);
  nand (_05779_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_05780_, _05779_, _05777_);
  and (_05781_, _05780_, _05776_);
  not (_05782_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_05783_, _05696_, _05782_);
  nand (_05784_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_05785_, _05784_, _05783_);
  and (_05786_, _05785_, _05781_);
  or (_05787_, _05786_, _05728_);
  nand (_05788_, _05787_, _05772_);
  not (_05789_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_05790_, _05718_, _05789_);
  not (_05791_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_05792_, _05705_, _05791_);
  not (_05793_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_05794_, _05711_, _05793_);
  and (_05795_, _05794_, _05792_);
  and (_05796_, _05795_, _05790_);
  nand (_05797_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  not (_05798_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_05799_, _05700_, _05798_);
  and (_05800_, _05799_, _05797_);
  not (_05801_, _05696_);
  and (_05802_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_05803_, _05802_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_05804_, _05803_, _05800_);
  nand (_05805_, _05804_, _05796_);
  or (_05806_, _05805_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05807_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05808_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not (_05809_, _05808_);
  and (_05810_, _05809_, _05806_);
  not (_05811_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_05812_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nand (_05813_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_05814_, _05813_, _05812_);
  not (_05815_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_05816_, _05696_, _05815_);
  not (_05817_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_05818_, _05718_, _05817_);
  and (_05819_, _05818_, _05816_);
  nand (_05820_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_05821_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_05822_, _05821_, _05820_);
  and (_05823_, _05822_, _05819_);
  nand (_05824_, _05823_, _05814_);
  nand (_05825_, _05824_, _05811_);
  nand (_05826_, _05825_, _05807_);
  nor (_05827_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _05807_);
  not (_05828_, _05827_);
  and (_05829_, _05828_, _05826_);
  nand (_05830_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand (_05831_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_05832_, _05831_, _05830_);
  not (_05833_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_05834_, _05696_, _05833_);
  not (_05835_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_05836_, _05718_, _05835_);
  and (_05837_, _05836_, _05834_);
  nand (_05838_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_05839_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_05840_, _05839_, _05838_);
  and (_05841_, _05840_, _05837_);
  nand (_05842_, _05841_, _05832_);
  nand (_05843_, _05842_, _05811_);
  nand (_05844_, _05843_, _05807_);
  nor (_05845_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not (_05846_, _05845_);
  and (_05847_, _05846_, _05844_);
  nor (_05848_, _05847_, _05829_);
  and (_05849_, _05848_, _05810_);
  and (_05850_, _05849_, _05788_);
  and (_05851_, _05850_, _05770_);
  not (_05852_, _05788_);
  and (_05853_, _05849_, _05852_);
  nor (_05854_, _05768_, _05747_);
  and (_05855_, _05854_, _05726_);
  and (_05856_, _05855_, _05853_);
  not (_05857_, _05847_);
  not (_05858_, _05810_);
  and (_05859_, _05829_, _05858_);
  and (_05860_, _05859_, _05857_);
  and (_05861_, _05860_, _05852_);
  not (_05862_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_05863_, _05696_, _05862_);
  and (_05864_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  not (_05865_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_05866_, _05718_, _05865_);
  and (_05867_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_05868_, _05867_, _05866_);
  nand (_05869_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nand (_05870_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_05871_, _05870_, _05869_);
  nand (_05872_, _05871_, _05868_);
  or (_05873_, _05872_, _05864_);
  or (_05874_, _05873_, _05863_);
  or (_05875_, _05874_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_05876_, _05875_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05878_, _05807_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not (_05879_, _05878_);
  and (_05880_, _05879_, _05876_);
  not (_05881_, _05880_);
  and (_05882_, _05881_, _05769_);
  and (_05883_, _05882_, _05861_);
  or (_05884_, _05883_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_05885_, _05884_, _05856_);
  or (_05886_, _05885_, _05851_);
  and (_05887_, _05886_, _05691_);
  nor (_05888_, _05690_, _05685_);
  or (_05889_, _05888_, rst);
  or (_00393_, _05889_, _05887_);
  and (_05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_05891_, _05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_05892_, _05891_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_05893_, _05892_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_05894_, _05893_);
  not (_05895_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05896_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05686_);
  and (_05897_, _05896_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_05898_, _05897_, _05895_);
  not (_05899_, _05898_);
  nor (_05900_, _05892_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_05901_, _05900_, _05899_);
  and (_05902_, _05901_, _05894_);
  not (_05903_, _05902_);
  nor (_05904_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor (_05905_, _05904_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_05906_, _05905_, _05896_);
  and (_05907_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  not (_05908_, _05907_);
  and (_05909_, _05897_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05910_, _05904_, _05896_);
  and (_05911_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_05912_, _05911_, _05909_);
  and (_05913_, _05912_, _05908_);
  not (_05914_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_05915_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05686_);
  and (_05916_, _05915_, _05914_);
  and (_05917_, _05916_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_05918_, _05917_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_05919_, _05916_, _05895_);
  and (_05920_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  nor (_05921_, _05920_, _05918_);
  and (_05922_, _05921_, _05913_);
  and (_05923_, _05922_, _05903_);
  and (_05924_, _05893_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_05925_, _05924_);
  nor (_05926_, _05893_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_05927_, _05926_, _05899_);
  and (_05928_, _05927_, _05925_);
  not (_05929_, _05928_);
  and (_05930_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_05931_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_05932_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or (_05933_, _05932_, _05931_);
  or (_05934_, _05933_, _05909_);
  nor (_05936_, _05934_, _05930_);
  and (_05937_, _05936_, _05929_);
  and (_05938_, _05937_, _05923_);
  and (_05939_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_05940_, _05939_);
  nor (_05941_, _05924_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_05943_, _05941_, _05899_);
  and (_05944_, _05943_, _05940_);
  not (_05945_, _05944_);
  and (_05946_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  not (_05947_, _05946_);
  and (_05948_, _05919_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_05949_, _05948_);
  and (_05950_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nor (_05951_, _05950_, _05909_);
  and (_05952_, _05951_, _05949_);
  and (_05953_, _05952_, _05947_);
  and (_05954_, _05953_, _05945_);
  not (_05955_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_05956_, _05939_, _05955_);
  and (_05957_, _05939_, _05955_);
  nor (_05958_, _05957_, _05956_);
  nor (_05959_, _05958_, _05899_);
  not (_05960_, _05959_);
  and (_05961_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_05962_, _05917_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and (_05963_, _05919_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or (_05964_, _05963_, _05962_);
  or (_05965_, _05964_, _05909_);
  nor (_05966_, _05965_, _05961_);
  and (_05967_, _05966_, _05960_);
  nor (_05968_, _05967_, _05954_);
  and (_05969_, _05968_, _05938_);
  nor (_05970_, _05890_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_05971_, _05970_, _05891_);
  and (_05972_, _05971_, _05898_);
  and (_05973_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_05975_, _05973_, _05972_);
  and (_05976_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_05977_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_05978_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_05979_, _05978_, _05977_);
  nor (_05980_, _05979_, _05976_);
  and (_05981_, _05980_, _05975_);
  not (_05982_, _05981_);
  nor (_05983_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_05984_, _05983_, _05890_);
  and (_05985_, _05984_, _05898_);
  and (_05986_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_05987_, _05986_, _05985_);
  and (_05988_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_05989_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_05990_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_05991_, _05990_, _05989_);
  nor (_05992_, _05991_, _05988_);
  and (_05993_, _05992_, _05987_);
  and (_05994_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_05995_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_05996_, _05995_, _05994_);
  not (_05997_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_05998_, _05898_, _05997_);
  not (_05999_, _05998_);
  and (_06000_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_06001_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_06002_, _06001_, _06000_);
  and (_06003_, _06002_, _05999_);
  and (_06004_, _06003_, _05996_);
  and (_06005_, _06004_, _05993_);
  and (_06006_, _06005_, _05982_);
  and (_06007_, _05896_, _05895_);
  not (_06008_, _06007_);
  not (_06009_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_06010_, \oc8051_top_1.oc8051_decoder1.wr , _05686_);
  and (_06011_, _06010_, _06009_);
  and (_06012_, _06011_, _06008_);
  not (_06013_, _06012_);
  not (_06014_, _05892_);
  nor (_06015_, _05891_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_06016_, _06015_, _05899_);
  and (_06017_, _06016_, _06014_);
  not (_06018_, _06017_);
  and (_06019_, _05917_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_06020_, _05910_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_06021_, _06020_, _06019_);
  and (_06022_, _05919_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_06023_, _05906_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_06024_, _06023_, _06022_);
  and (_06025_, _06024_, _06021_);
  and (_06026_, _06025_, _06018_);
  nor (_06027_, _06026_, _06013_);
  and (_06028_, _06027_, _06006_);
  and (_06029_, _06028_, _05969_);
  not (_06030_, _06004_);
  and (_06031_, _06030_, _05993_);
  and (_06032_, _06031_, _05982_);
  and (_06033_, _06027_, _05969_);
  and (_06035_, _06033_, _06032_);
  nor (_06036_, _06035_, _06029_);
  and (_06037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_06038_, _06037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_06039_, _06038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_06040_, _06039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_06041_, _06040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_06042_, _06041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_06043_, _06042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_06044_, _06043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_06045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_06046_, _06045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_06047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_06048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_06050_, _06048_, _06047_);
  and (_06051_, _06050_, _06046_);
  and (_06053_, _06051_, _06044_);
  nor (_06054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_06055_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_06056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_06057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _06056_);
  and (_06058_, _06057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_06059_, _06058_, _06055_);
  not (_06061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_06062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_06064_, _06062_, _06054_);
  and (_06065_, _06064_, _06061_);
  not (_06066_, _06065_);
  and (_06067_, _06066_, _06059_);
  and (_06068_, _06067_, _06054_);
  nand (_06069_, _06068_, _06053_);
  nand (_06070_, _06069_, _06036_);
  not (_06071_, rst);
  or (_06072_, _06036_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_06073_, _06072_, _06071_);
  and (_05877_, _06073_, _06070_);
  not (_06075_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  not (_06076_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06077_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06076_);
  or (_06078_, _06077_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06079_, _06078_, _06075_);
  not (_06080_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  not (_06081_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_06082_, _06081_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06083_, _06082_, _06076_);
  or (_06084_, _06083_, _06080_);
  and (_06085_, _06084_, _06079_);
  not (_06086_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_06087_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06088_, _06087_, _06081_);
  or (_06089_, _06088_, _06086_);
  not (_06090_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_06091_, _06077_, _06081_);
  or (_06093_, _06091_, _06090_);
  and (_06094_, _06093_, _06089_);
  and (_06095_, _06094_, _06085_);
  or (_06097_, _06087_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_06098_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_06099_, _06098_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06100_, _06099_, ABINPUT[8]);
  nand (_06101_, _06098_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06102_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_06103_, _06102_, _06100_);
  or (_06104_, _06103_, _06097_);
  not (_06105_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_06106_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_06107_, _06106_, _06081_);
  or (_06108_, _06107_, _06105_);
  and (_06109_, _06106_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06110_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_06111_, _06110_, _06108_);
  and (_06112_, _06111_, _06104_);
  and (_06113_, _06112_, _06095_);
  and (_06114_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_06115_, _06114_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor (_06116_, _06099_, ABINPUT[0]);
  nor (_06117_, _06101_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_06118_, _06117_, _06116_);
  nor (_06119_, _06118_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_06120_, _06119_, _06115_);
  and (_06121_, _06120_, _06113_);
  not (_06122_, _06121_);
  and (_06123_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05686_);
  and (_06124_, _06123_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06125_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05686_);
  and (_06126_, _06125_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06127_, _06126_, _06124_);
  not (_06128_, _06127_);
  or (_06129_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06131_, _06129_, _06103_);
  nand (_06132_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06133_, _06132_, _06075_);
  not (_06134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_06135_, _06134_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06136_, _06135_, _06105_);
  and (_06137_, _06136_, _06133_);
  and (_06138_, _06137_, _06131_);
  not (_06139_, _06138_);
  nor (_06140_, _06139_, _06120_);
  nor (_06141_, _06140_, _06128_);
  and (_06142_, _06141_, _06122_);
  not (_06143_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06144_, _06123_, _06143_);
  and (_06145_, _06144_, _06126_);
  not (_06146_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  or (_06147_, _06078_, _06146_);
  not (_06148_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or (_06149_, _06083_, _06148_);
  and (_06150_, _06149_, _06147_);
  not (_06151_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_06152_, _06088_, _06151_);
  not (_06153_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_06154_, _06091_, _06153_);
  and (_06155_, _06154_, _06152_);
  and (_06156_, _06155_, _06150_);
  or (_06157_, _06099_, ABINPUT[5]);
  or (_06158_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_06159_, _06158_, _06157_);
  or (_06160_, _06159_, _06097_);
  not (_06161_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_06162_, _06107_, _06161_);
  nand (_06163_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_06164_, _06163_, _06162_);
  and (_06165_, _06164_, _06160_);
  and (_06166_, _06165_, _06156_);
  not (_06167_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  or (_06168_, _06083_, _06167_);
  not (_06169_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  or (_06170_, _06078_, _06169_);
  and (_06171_, _06170_, _06168_);
  not (_06172_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_06173_, _06088_, _06172_);
  not (_06174_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_06175_, _06091_, _06174_);
  and (_06176_, _06175_, _06173_);
  and (_06177_, _06176_, _06171_);
  or (_06178_, _06099_, ABINPUT[4]);
  or (_06179_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_06180_, _06179_, _06178_);
  or (_06181_, _06180_, _06097_);
  nand (_06182_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not (_06183_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06184_, _06107_, _06183_);
  and (_06185_, _06184_, _06182_);
  and (_06186_, _06185_, _06181_);
  and (_06187_, _06186_, _06177_);
  not (_06188_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  or (_06189_, _06078_, _06188_);
  not (_06190_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  or (_06191_, _06083_, _06190_);
  and (_06192_, _06191_, _06189_);
  not (_06193_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_06194_, _06088_, _06193_);
  not (_06195_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_06196_, _06091_, _06195_);
  nor (_06197_, _06196_, _06194_);
  and (_06198_, _06197_, _06192_);
  or (_06200_, _06099_, ABINPUT[1]);
  or (_06201_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_06202_, _06201_, _06200_);
  or (_06203_, _06202_, _06097_);
  not (_06204_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_06205_, _06107_, _06204_);
  and (_06206_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_06207_, _06206_, _06205_);
  and (_06208_, _06207_, _06203_);
  and (_06209_, _06208_, _06198_);
  not (_06210_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_06211_, _06088_, _06210_);
  nand (_06212_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_06213_, _06212_, _06211_);
  not (_06214_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or (_06215_, _06083_, _06214_);
  not (_06216_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_06217_, _06091_, _06216_);
  and (_06218_, _06217_, _06215_);
  and (_06219_, _06218_, _06213_);
  or (_06220_, _06099_, ABINPUT[2]);
  or (_06221_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_06222_, _06221_, _06220_);
  or (_06223_, _06222_, _06097_);
  not (_06224_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  or (_06225_, _06078_, _06224_);
  not (_06226_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_06227_, _06107_, _06226_);
  and (_06228_, _06227_, _06225_);
  and (_06229_, _06228_, _06223_);
  nand (_06230_, _06229_, _06219_);
  not (_06231_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or (_06232_, _06083_, _06231_);
  not (_06233_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  or (_06234_, _06078_, _06233_);
  and (_06235_, _06234_, _06232_);
  nand (_06236_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not (_06237_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06238_, _06107_, _06237_);
  and (_06239_, _06238_, _06236_);
  and (_06240_, _06239_, _06235_);
  not (_06241_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_06242_, _06091_, _06241_);
  not (_06243_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_06244_, _06088_, _06243_);
  and (_06245_, _06244_, _06242_);
  or (_06246_, _06099_, ABINPUT[3]);
  or (_06247_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_06248_, _06247_, _06246_);
  or (_06249_, _06248_, _06097_);
  and (_06250_, _06249_, _06245_);
  nand (_06251_, _06250_, _06240_);
  nor (_06252_, _06251_, _06230_);
  and (_06253_, _06252_, _06209_);
  and (_06254_, _06253_, _06187_);
  and (_06255_, _06254_, _06166_);
  not (_06256_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_06257_, _06078_, _06256_);
  not (_06258_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  or (_06259_, _06083_, _06258_);
  and (_06260_, _06259_, _06257_);
  not (_06261_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_06262_, _06088_, _06261_);
  not (_06263_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_06264_, _06091_, _06263_);
  and (_06265_, _06264_, _06262_);
  and (_06266_, _06265_, _06260_);
  or (_06267_, _06099_, ABINPUT[7]);
  or (_06268_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_06269_, _06268_, _06267_);
  or (_06270_, _06269_, _06097_);
  not (_06271_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06272_, _06107_, _06271_);
  nand (_06273_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_06274_, _06273_, _06272_);
  and (_06275_, _06274_, _06270_);
  and (_06276_, _06275_, _06266_);
  not (_06277_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  or (_06278_, _06083_, _06277_);
  not (_06279_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  or (_06280_, _06078_, _06279_);
  and (_06281_, _06280_, _06278_);
  not (_06282_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_06283_, _06091_, _06282_);
  not (_06284_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_06285_, _06088_, _06284_);
  and (_06286_, _06285_, _06283_);
  and (_06287_, _06286_, _06281_);
  or (_06288_, _06099_, ABINPUT[6]);
  or (_06289_, _06101_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_06290_, _06289_, _06288_);
  or (_06291_, _06290_, _06097_);
  not (_06292_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_06293_, _06107_, _06292_);
  nand (_06294_, _06109_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_06295_, _06294_, _06293_);
  and (_06296_, _06295_, _06291_);
  nand (_06297_, _06296_, _06287_);
  not (_06298_, _06297_);
  and (_06299_, _06298_, _06276_);
  and (_06300_, _06299_, _06255_);
  nor (_06301_, _06300_, _06120_);
  not (_06302_, _06120_);
  not (_06303_, _06276_);
  not (_06304_, _06166_);
  not (_06305_, _06187_);
  not (_06306_, _06209_);
  and (_06307_, _06230_, _06306_);
  and (_06308_, _06251_, _06307_);
  and (_06309_, _06308_, _06305_);
  and (_06310_, _06309_, _06304_);
  and (_06311_, _06297_, _06310_);
  and (_06312_, _06311_, _06303_);
  nor (_06313_, _06312_, _06302_);
  or (_06314_, _06313_, _06301_);
  and (_06315_, _06314_, _06113_);
  nor (_06316_, _06314_, _06113_);
  nor (_06317_, _06316_, _06315_);
  and (_06318_, _06317_, _06145_);
  nor (_06319_, _06318_, _06142_);
  and (_06320_, _05686_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  nor (_06321_, _06320_, _06123_);
  not (_06322_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06323_, _06125_, _06322_);
  and (_06324_, _06323_, _06321_);
  and (_06325_, _06138_, _06113_);
  nor (_06326_, _06138_, _06113_);
  nor (_06327_, _06326_, _06325_);
  and (_06328_, _06327_, _06324_);
  not (_06329_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06330_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05686_);
  and (_06331_, _06330_, _06329_);
  and (_06332_, _06331_, _06124_);
  and (_06333_, _06332_, _06326_);
  not (_06334_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_06335_, _06320_, _06334_);
  and (_06336_, _06335_, _06323_);
  not (_06337_, _06336_);
  nor (_06338_, _06337_, _06325_);
  and (_06339_, _06331_, _06144_);
  and (_06340_, _06339_, _06113_);
  or (_06341_, _06340_, _06338_);
  or (_06342_, _06341_, _06333_);
  nor (_06343_, _06342_, _06328_);
  nor (_06344_, _06330_, _06125_);
  and (_06345_, _06344_, _06320_);
  and (_06347_, _06331_, _06334_);
  nor (_06348_, _06347_, _06345_);
  and (_06349_, _06344_, _06321_);
  and (_06350_, _06126_, _06334_);
  nor (_06351_, _06350_, _06349_);
  and (_06352_, _06323_, _06123_);
  not (_06353_, _06352_);
  and (_06354_, _06353_, _06351_);
  and (_06355_, _06354_, _06348_);
  nor (_06356_, _06355_, _06113_);
  not (_06357_, _06356_);
  and (_06358_, _06357_, _06343_);
  and (_06359_, _06358_, _06319_);
  not (_06360_, _06359_);
  and (_06361_, _05993_, _05981_);
  and (_06362_, _06361_, _06030_);
  and (_06363_, _06362_, _06026_);
  not (_06364_, _05923_);
  and (_06365_, _05937_, _06364_);
  and (_06366_, _05967_, _05954_);
  and (_06367_, _06366_, _06365_);
  and (_06368_, _06367_, _06363_);
  and (_06369_, _06368_, _06011_);
  and (_06370_, _06369_, _06360_);
  and (_06371_, _06026_, _05981_);
  and (_06372_, _06371_, _06005_);
  and (_06373_, _06366_, _05938_);
  and (_06374_, _06373_, _06372_);
  and (_06375_, _06373_, _06363_);
  nor (_06376_, _06375_, _06374_);
  and (_06377_, _06372_, _06367_);
  not (_06378_, _06026_);
  and (_06380_, _06362_, _06378_);
  and (_06381_, _06380_, _06373_);
  nor (_06382_, _06381_, _06377_);
  and (_06383_, _06005_, _05981_);
  and (_06384_, _06383_, _06378_);
  and (_06385_, _06384_, _06373_);
  not (_06386_, _06385_);
  and (_06387_, _06386_, _06382_);
  and (_06388_, _06387_, _06376_);
  not (_06389_, _06388_);
  not (_06390_, _06011_);
  or (_06391_, _06377_, _06368_);
  and (_06392_, _06373_, _06361_);
  nor (_06393_, _06392_, _06391_);
  or (_06394_, _06393_, _06390_);
  or (_06395_, _06394_, _06389_);
  and (_06396_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or (_06397_, _06396_, _06370_);
  and (_09300_, _06397_, _06071_);
  and (_06398_, _06380_, _06367_);
  and (_06399_, _06398_, _06011_);
  not (_06400_, _06399_);
  and (_06401_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_06402_, _06400_, _06359_);
  or (_06403_, _06402_, _06401_);
  and (_12917_, _06403_, _06071_);
  or (_06404_, _06248_, _06129_);
  or (_06405_, _06132_, _06233_);
  or (_06406_, _06135_, _06237_);
  and (_06407_, _06406_, _06405_);
  nand (_06408_, _06407_, _06404_);
  and (_06409_, _06408_, _06127_);
  nor (_06410_, _06209_, _06120_);
  nor (_06411_, _06230_, _06120_);
  nor (_06412_, _06411_, _06307_);
  nor (_06413_, _06412_, _06410_);
  and (_06414_, _06413_, _06251_);
  nor (_06415_, _06413_, _06251_);
  nor (_06416_, _06415_, _06414_);
  and (_06417_, _06416_, _06145_);
  nor (_06418_, _06417_, _06409_);
  nor (_06419_, _06408_, _06251_);
  nor (_06420_, _06419_, _06337_);
  and (_06421_, _06408_, _06251_);
  nor (_06422_, _06421_, _06419_);
  and (_06423_, _06422_, _06324_);
  nor (_06424_, _06423_, _06420_);
  and (_06425_, _06421_, _06332_);
  not (_06426_, _06339_);
  nor (_06427_, _06426_, _06251_);
  nor (_06428_, _06427_, _06425_);
  not (_06429_, _06251_);
  nor (_06430_, _06355_, _06429_);
  not (_06431_, _06430_);
  and (_06432_, _06431_, _06428_);
  and (_06433_, _06432_, _06424_);
  and (_06434_, _06433_, _06418_);
  not (_06435_, _06434_);
  and (_06436_, _06435_, _06377_);
  not (_06437_, _06392_);
  nor (_06438_, _06388_, _06390_);
  nand (_06439_, _06438_, _06437_);
  and (_06440_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_06441_, _06440_, _06436_);
  or (_06442_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_06443_, _06442_, _06071_);
  and (_12997_, _06443_, _06441_);
  not (_06444_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _06445_);
  and (_06447_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_06448_, _06447_, _06446_);
  and (_06449_, _06448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_06450_, _06449_, _06444_);
  and (_06451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_06452_, _06451_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_06453_, _06452_);
  and (_06454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_06455_, _06454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_06457_, _06456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor (_06458_, _06457_, _06455_);
  and (_06459_, _06458_, _06453_);
  nor (_06460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  not (_06461_, _06460_);
  and (_06462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_06463_, _06462_, _06461_);
  not (_06464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_06465_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_06466_, _06465_, _06464_);
  and (_06467_, _06466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor (_06468_, _06467_, _06463_);
  and (_06469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_06470_, _06469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_06471_, _06470_);
  and (_06472_, _06471_, _06468_);
  and (_06473_, _06472_, _06459_);
  nor (_06474_, _06473_, _06450_);
  and (_06475_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _06444_);
  not (_06476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_06477_, _06476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_06478_, _06477_, _06461_);
  not (_06479_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_06480_, _06466_, _06479_);
  nor (_06481_, _06480_, _06478_);
  not (_06482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_06483_, _06469_, _06482_);
  not (_06484_, _06483_);
  nand (_06485_, _06484_, _06481_);
  and (_06486_, _06485_, _06475_);
  or (_06487_, _06486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not (_06488_, _06475_);
  not (_06489_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_06490_, _06451_, _06489_);
  not (_06491_, _06490_);
  not (_06492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_06493_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_06494_, _06493_, _06492_);
  not (_06495_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06496_, _06454_, _06495_);
  nor (_06497_, _06496_, _06494_);
  and (_06498_, _06497_, _06491_);
  or (_06499_, _06498_, _06488_);
  or (_06500_, _06499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06501_, _06500_, _06487_);
  or (_06502_, _06501_, _06474_);
  not (_06503_, _06472_);
  or (_06504_, _06459_, _06450_);
  or (_06505_, _06504_, _06503_);
  and (_06506_, _06505_, _06445_);
  or (_06507_, _06506_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_06508_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_06509_, _06508_);
  and (_06510_, _06509_, _06504_);
  nor (_06511_, _06508_, _06445_);
  or (_06512_, _06511_, _06510_);
  and (_06513_, _06512_, _06507_);
  and (_06514_, _06513_, _06502_);
  and (_06515_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_06516_, _06515_, _06514_);
  and (_00316_, _06516_, _06071_);
  and (_06517_, _06498_, _06484_);
  nand (_06518_, _06517_, _06481_);
  and (_06519_, _06518_, _06475_);
  nand (_06520_, _06473_, _06444_);
  or (_06521_, _06520_, _06519_);
  nor (_06522_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06445_);
  nand (_06523_, _06522_, _06508_);
  and (_06524_, _06523_, _06071_);
  and (_00503_, _06524_, _06521_);
  and (_06525_, _05704_, _05694_);
  nor (_06526_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_06527_, _06526_, _05686_);
  not (_06528_, _06527_);
  nor (_06529_, _06528_, _06525_);
  nor (_06530_, _06529_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_06531_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not (_06532_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_06533_, _06530_, _06532_);
  and (_06534_, _06533_, _06071_);
  and (_00572_, _06534_, _06531_);
  and (_06535_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_06536_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_06537_, _06059_, _06044_);
  and (_06538_, _06537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_06539_, _06046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_06540_, _06539_, _06538_);
  and (_06541_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_06542_, _06541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_06543_, _06540_, _06047_);
  and (_06544_, _06543_, _06542_);
  and (_06545_, _06054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_06546_, _06545_);
  and (_06547_, _06546_, _06053_);
  and (_06548_, _06547_, _06059_);
  and (_06549_, _06548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_06550_, _06549_, _06065_);
  or (_06551_, _06550_, _06544_);
  and (_06552_, _06551_, _06536_);
  and (_06553_, _06552_, _06036_);
  or (_06554_, _06553_, _06535_);
  not (_06555_, _06035_);
  nor (_06556_, _06359_, _06555_);
  or (_06557_, _06556_, _06554_);
  and (_01048_, _06557_, _06071_);
  nor (_06558_, rst, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_06559_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_06560_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_06561_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_01756_, _06561_, _06559_);
  nor (_06562_, _06519_, _06474_);
  and (_06563_, _06562_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_06564_, _06474_);
  and (_06565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06445_);
  nor (_06566_, _06565_, _06522_);
  nor (_06567_, _06566_, _06564_);
  or (_06568_, _06567_, _06508_);
  or (_06569_, _06568_, _06563_);
  or (_06570_, _06566_, _06509_);
  and (_06571_, _06570_, _06071_);
  and (_01890_, _06571_, _06569_);
  and (_06572_, _06297_, _06120_);
  or (_06573_, _06290_, _06129_);
  or (_06574_, _06132_, _06279_);
  or (_06575_, _06135_, _06292_);
  and (_06576_, _06575_, _06574_);
  and (_06577_, _06576_, _06573_);
  nor (_06578_, _06577_, _06120_);
  or (_06579_, _06578_, _06572_);
  and (_06580_, _06579_, _06127_);
  and (_06581_, _06310_, _06120_);
  and (_06582_, _06255_, _06302_);
  nor (_06583_, _06582_, _06581_);
  and (_06584_, _06583_, _06298_);
  not (_06585_, _06145_);
  nor (_06586_, _06583_, _06298_);
  or (_06587_, _06586_, _06585_);
  nor (_06588_, _06587_, _06584_);
  nor (_06590_, _06588_, _06580_);
  nor (_06591_, _06355_, _06298_);
  not (_06592_, _06591_);
  nand (_06593_, _06576_, _06573_);
  and (_06594_, _06593_, _06297_);
  nor (_06595_, _06593_, _06297_);
  nor (_06596_, _06595_, _06594_);
  and (_06597_, _06596_, _06324_);
  not (_06598_, _06597_);
  nor (_06599_, _06595_, _06337_);
  not (_06600_, _06599_);
  and (_06601_, _06594_, _06332_);
  nor (_06602_, _06426_, _06297_);
  nor (_06603_, _06602_, _06601_);
  and (_06605_, _06603_, _06600_);
  and (_06607_, _06605_, _06598_);
  and (_06608_, _06607_, _06592_);
  and (_06609_, _06608_, _06590_);
  and (_06610_, _06385_, _06011_);
  not (_06611_, _06610_);
  nor (_06612_, _06611_, _06609_);
  and (_06613_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_06614_, _06613_, _06612_);
  and (_02186_, _06614_, _06071_);
  and (_06615_, _06344_, _06144_);
  not (_06616_, _06615_);
  and (_06618_, _06139_, _06113_);
  or (_06619_, _06269_, _06129_);
  or (_06620_, _06132_, _06256_);
  or (_06621_, _06135_, _06271_);
  and (_06622_, _06621_, _06620_);
  nand (_06623_, _06622_, _06619_);
  nor (_06624_, _06623_, _06276_);
  not (_06625_, _06623_);
  nor (_06626_, _06625_, _06276_);
  and (_06627_, _06625_, _06276_);
  nor (_06628_, _06627_, _06626_);
  and (_06629_, _06577_, _06297_);
  or (_06630_, _06159_, _06129_);
  or (_06631_, _06132_, _06146_);
  or (_06632_, _06135_, _06161_);
  and (_06633_, _06632_, _06631_);
  nand (_06634_, _06633_, _06630_);
  and (_06635_, _06634_, _06166_);
  nor (_06636_, _06635_, _06596_);
  nor (_06637_, _06636_, _06629_);
  nor (_06638_, _06637_, _06628_);
  nor (_06639_, _06638_, _06624_);
  and (_06640_, _06637_, _06628_);
  nor (_06641_, _06640_, _06638_);
  not (_06642_, _06641_);
  and (_06643_, _06635_, _06596_);
  nor (_06644_, _06643_, _06636_);
  not (_06645_, _06644_);
  and (_06646_, _06633_, _06630_);
  nor (_06647_, _06646_, _06166_);
  and (_06648_, _06646_, _06166_);
  nor (_06649_, _06648_, _06647_);
  not (_06650_, _06649_);
  or (_06651_, _06180_, _06129_);
  or (_06652_, _06132_, _06169_);
  or (_06653_, _06135_, _06183_);
  and (_06654_, _06653_, _06652_);
  and (_06655_, _06654_, _06651_);
  and (_06656_, _06655_, _06187_);
  nor (_06657_, _06655_, _06187_);
  nor (_06659_, _06657_, _06656_);
  and (_06660_, _06407_, _06404_);
  and (_06661_, _06660_, _06251_);
  or (_06662_, _06222_, _06129_);
  or (_06663_, _06132_, _06224_);
  or (_06664_, _06135_, _06226_);
  and (_06665_, _06664_, _06663_);
  nand (_06666_, _06665_, _06662_);
  and (_06667_, _06666_, _06230_);
  nor (_06668_, _06666_, _06230_);
  nor (_06669_, _06668_, _06667_);
  or (_06670_, _06202_, _06129_);
  or (_06671_, _06132_, _06188_);
  or (_06672_, _06135_, _06204_);
  and (_06673_, _06672_, _06671_);
  nand (_06674_, _06673_, _06670_);
  and (_06675_, _06674_, _06209_);
  nor (_06676_, _06675_, _06669_);
  and (_06677_, _06665_, _06662_);
  and (_06678_, _06677_, _06230_);
  nor (_06680_, _06678_, _06676_);
  nor (_06681_, _06680_, _06422_);
  nor (_06682_, _06681_, _06661_);
  nor (_06683_, _06682_, _06659_);
  and (_06684_, _06682_, _06659_);
  nor (_06685_, _06684_, _06683_);
  and (_06686_, _06680_, _06422_);
  nor (_06687_, _06686_, _06681_);
  and (_06688_, _06675_, _06669_);
  nor (_06689_, _06688_, _06676_);
  and (_06690_, _06673_, _06670_);
  nor (_06691_, _06690_, _06209_);
  and (_06692_, _06690_, _06209_);
  nor (_06693_, _06692_, _06691_);
  nor (_06694_, _06693_, _06120_);
  not (_06695_, _06694_);
  nor (_06696_, _06695_, _06689_);
  not (_06697_, _06696_);
  nor (_06698_, _06697_, _06687_);
  not (_06699_, _06698_);
  nor (_06700_, _06699_, _06685_);
  nand (_06701_, _06654_, _06651_);
  or (_06702_, _06701_, _06187_);
  and (_06703_, _06701_, _06187_);
  or (_06704_, _06682_, _06703_);
  and (_06705_, _06704_, _06702_);
  or (_06706_, _06705_, _06700_);
  and (_06707_, _06706_, _06650_);
  and (_06708_, _06707_, _06645_);
  and (_06709_, _06708_, _06642_);
  nor (_06710_, _06709_, _06639_);
  nor (_06711_, _06710_, _06327_);
  nor (_06712_, _06711_, _06618_);
  nor (_06713_, _06712_, _06616_);
  not (_06714_, _06713_);
  and (_06715_, _06344_, _06335_);
  not (_06716_, _06715_);
  not (_06717_, _06326_);
  not (_06718_, _06422_);
  and (_06719_, _06691_, _06669_);
  nor (_06720_, _06719_, _06667_);
  nor (_06721_, _06720_, _06718_);
  nor (_06722_, _06721_, _06421_);
  nor (_06723_, _06722_, _06659_);
  and (_06724_, _06722_, _06659_);
  nor (_06725_, _06724_, _06723_);
  and (_06726_, _06693_, _06302_);
  and (_06727_, _06726_, _06669_);
  and (_06728_, _06720_, _06718_);
  nor (_06729_, _06728_, _06721_);
  and (_06730_, _06729_, _06727_);
  not (_06731_, _06730_);
  nor (_06732_, _06731_, _06725_);
  nor (_06733_, _06722_, _06656_);
  or (_06734_, _06733_, _06657_);
  or (_06735_, _06734_, _06732_);
  and (_06736_, _06735_, _06649_);
  and (_06737_, _06736_, _06596_);
  not (_06738_, _06628_);
  and (_06739_, _06647_, _06596_);
  nor (_06740_, _06739_, _06594_);
  nor (_06741_, _06740_, _06738_);
  and (_06742_, _06740_, _06738_);
  nor (_06743_, _06742_, _06741_);
  and (_06744_, _06743_, _06737_);
  not (_06745_, _06744_);
  nor (_06746_, _06741_, _06626_);
  and (_06747_, _06746_, _06745_);
  or (_06748_, _06747_, _06325_);
  and (_06749_, _06748_, _06717_);
  nor (_06750_, _06749_, _06716_);
  and (_06751_, _06335_, _06331_);
  nor (_06752_, _06252_, _06187_);
  and (_06753_, _06752_, _06751_);
  and (_06754_, _06753_, _06304_);
  nor (_06755_, _06754_, _06297_);
  and (_06756_, _06276_, _06120_);
  and (_06757_, _06756_, _06755_);
  nor (_06758_, _06757_, _06121_);
  not (_06759_, _06751_);
  and (_06760_, _06755_, _06276_);
  nor (_06761_, _06120_, _06113_);
  not (_06762_, _06761_);
  nor (_06763_, _06762_, _06760_);
  nor (_06764_, _06763_, _06759_);
  and (_06765_, _06764_, _06758_);
  not (_06766_, _06118_);
  nor (_06767_, _06753_, _06302_);
  and (_06768_, _06767_, _06766_);
  nor (_06769_, _06115_, _06766_);
  not (_06770_, _06324_);
  nor (_06771_, _06770_, _06769_);
  nor (_06772_, _06771_, _06336_);
  not (_06773_, _06772_);
  nor (_06774_, _06773_, _06753_);
  nor (_06775_, _06774_, _06768_);
  not (_06776_, _06113_);
  and (_06777_, _06323_, _06124_);
  and (_06779_, _06777_, _06776_);
  and (_06780_, _06115_, _06118_);
  and (_06781_, _06323_, _06144_);
  and (_06782_, _06332_, _06118_);
  nor (_06784_, _06782_, _06781_);
  nor (_06785_, _06784_, _06780_);
  nor (_06786_, _06785_, _06779_);
  and (_06787_, _06335_, _06126_);
  and (_06788_, _06787_, _06306_);
  and (_06789_, _06321_, _06126_);
  and (_06790_, _06789_, _06766_);
  nor (_06791_, _06790_, _06349_);
  and (_06792_, _06791_, _06302_);
  and (_06793_, _06426_, _06120_);
  nor (_06794_, _06793_, _06792_);
  nor (_06795_, _06794_, _06788_);
  and (_06796_, _06795_, _06786_);
  not (_06797_, _06796_);
  nor (_06798_, _06797_, _06775_);
  not (_06799_, _06798_);
  nor (_06800_, _06799_, _06765_);
  not (_06801_, _06800_);
  nor (_06802_, _06801_, _06750_);
  and (_06803_, _06802_, _06714_);
  nor (_06804_, _06004_, _05993_);
  and (_06805_, _06804_, _05982_);
  and (_06806_, _05954_, _05937_);
  not (_06807_, _05967_);
  nor (_06808_, _06378_, _05923_);
  and (_06809_, _06808_, _06807_);
  and (_06810_, _06809_, _06806_);
  and (_06812_, _06810_, _06805_);
  nand (_06813_, _06812_, _06803_);
  and (_06814_, _06010_, _06008_);
  and (_06815_, _06814_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  or (_06816_, _06812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06817_, _06816_, _06815_);
  and (_06818_, _06817_, _06813_);
  not (_06819_, _05954_);
  nor (_06820_, _05967_, _06819_);
  and (_06821_, _06820_, _06365_);
  and (_06822_, _06821_, _06372_);
  nand (_06823_, _06822_, _06359_);
  or (_06824_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_06825_, _06824_, _06012_);
  and (_06826_, _06825_, _06823_);
  not (_06827_, _06814_);
  and (_06828_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_06829_, _06828_, rst);
  or (_06830_, _06829_, _06826_);
  or (_03745_, _06830_, _06818_);
  nor (_06831_, t2ex_i, rst);
  and (_04082_, _06831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  and (_06832_, _06026_, _05923_);
  and (_06833_, _06832_, _06807_);
  and (_06834_, _06833_, _06806_);
  and (_06835_, _06834_, _06805_);
  nand (_06836_, _06835_, _06803_);
  or (_06837_, _06835_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_06838_, _06837_, _06815_);
  and (_06839_, _06838_, _06836_);
  and (_06840_, _06820_, _05938_);
  and (_06841_, _06840_, _06372_);
  nand (_06842_, _06841_, _06359_);
  or (_06843_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_06844_, _06843_, _06012_);
  and (_06845_, _06844_, _06842_);
  and (_06846_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_06847_, _06846_, rst);
  or (_06848_, _06847_, _06845_);
  or (_05680_, _06848_, _06839_);
  or (_06849_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not (_06850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_06851_, _06530_, _06850_);
  and (_06852_, _06851_, _06071_);
  and (_05681_, _06852_, _06849_);
  nor (_06853_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_06854_, _06853_);
  and (_06855_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  not (_06856_, _06230_);
  not (_06857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_06858_, _06857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_06859_, _06858_);
  or (_06860_, _06859_, _06660_);
  not (_06861_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_06862_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _06861_);
  not (_06863_, _06862_);
  or (_06864_, _06863_, _06646_);
  and (_06865_, _06864_, _06860_);
  or (_06866_, _06862_, _06858_);
  or (_06867_, _06866_, _06690_);
  and (_06868_, _06867_, _06854_);
  nand (_06869_, _06868_, _06865_);
  or (_06870_, _06854_, _06623_);
  nand (_06871_, _06870_, _06869_);
  or (_06872_, _06871_, _06856_);
  or (_06873_, _06859_, _06655_);
  or (_06874_, _06863_, _06577_);
  and (_06875_, _06874_, _06873_);
  or (_06876_, _06866_, _06677_);
  and (_06877_, _06876_, _06854_);
  nand (_06878_, _06877_, _06875_);
  nand (_06879_, _06853_, _06138_);
  nand (_06880_, _06879_, _06878_);
  or (_06881_, _06880_, _06209_);
  nor (_06882_, _06881_, _06872_);
  and (_06883_, _06879_, _06878_);
  and (_06884_, _06883_, _06230_);
  and (_06885_, _06870_, _06869_);
  and (_06886_, _06885_, _06251_);
  nand (_06887_, _06886_, _06884_);
  or (_06888_, _06886_, _06884_);
  and (_06889_, _06888_, _06887_);
  and (_06890_, _06889_, _06882_);
  and (_06891_, _06885_, _06305_);
  and (_06892_, _06883_, _06251_);
  and (_06893_, _06892_, _06872_);
  nand (_06894_, _06893_, _06891_);
  or (_06895_, _06893_, _06891_);
  and (_06896_, _06895_, _06894_);
  and (_06897_, _06896_, _06890_);
  nand (_06898_, _06894_, _06887_);
  or (_06899_, _06880_, _06187_);
  or (_06900_, _06871_, _06166_);
  or (_06901_, _06900_, _06899_);
  nand (_06902_, _06900_, _06899_);
  and (_06903_, _06902_, _06901_);
  nand (_06904_, _06903_, _06898_);
  or (_06905_, _06903_, _06898_);
  and (_06906_, _06905_, _06904_);
  nand (_06907_, _06906_, _06897_);
  or (_06908_, _06906_, _06897_);
  and (_06910_, _06908_, _06907_);
  nand (_06911_, _06910_, _06855_);
  and (_06912_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nand (_06913_, _06896_, _06890_);
  or (_06914_, _06896_, _06890_);
  and (_06915_, _06914_, _06913_);
  nand (_06916_, _06915_, _06912_);
  and (_06917_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_06918_, _06889_, _06882_);
  nor (_06919_, _06918_, _06890_);
  nand (_06920_, _06919_, _06917_);
  or (_06921_, _06915_, _06912_);
  nand (_06922_, _06921_, _06916_);
  or (_06923_, _06922_, _06920_);
  and (_06924_, _06923_, _06916_);
  or (_06925_, _06910_, _06855_);
  nand (_06926_, _06925_, _06911_);
  or (_06927_, _06926_, _06924_);
  and (_06928_, _06927_, _06911_);
  and (_06929_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  and (_06930_, _06906_, _06897_);
  and (_06931_, _06903_, _06898_);
  and (_06932_, _06883_, _06304_);
  and (_06933_, _06932_, _06891_);
  or (_06934_, _06880_, _06298_);
  or (_06935_, _06934_, _06900_);
  and (_06936_, _06885_, _06297_);
  or (_06937_, _06936_, _06932_);
  and (_06938_, _06937_, _06935_);
  nand (_06939_, _06938_, _06933_);
  or (_06940_, _06938_, _06933_);
  and (_06941_, _06940_, _06939_);
  nand (_06942_, _06941_, _06931_);
  or (_06943_, _06941_, _06931_);
  and (_06944_, _06943_, _06942_);
  nand (_06945_, _06944_, _06930_);
  or (_06946_, _06944_, _06930_);
  and (_06947_, _06946_, _06945_);
  nand (_06948_, _06947_, _06929_);
  or (_06949_, _06947_, _06929_);
  nand (_06951_, _06949_, _06948_);
  or (_06952_, _06951_, _06928_);
  not (_06954_, _06952_);
  and (_06955_, _06951_, _06928_);
  nor (_06956_, _06955_, _06954_);
  and (_05682_, _06956_, _06071_);
  or (_06957_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not (_06958_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_06959_, _06530_, _06958_);
  and (_06960_, _06959_, _06071_);
  and (_05683_, _06960_, _06957_);
  or (_06961_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not (_06962_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_06963_, _06530_, _06962_);
  and (_06964_, _06963_, _06071_);
  and (_05684_, _06964_, _06961_);
  and (_06965_, _06384_, _06367_);
  and (_06966_, _06965_, _06011_);
  not (_06967_, _06966_);
  and (_06968_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_06969_, _06166_, _06302_);
  nor (_06970_, _06646_, _06120_);
  or (_06971_, _06970_, _06969_);
  and (_06972_, _06971_, _06127_);
  nor (_06973_, _06309_, _06302_);
  nor (_06974_, _06254_, _06120_);
  nor (_06975_, _06974_, _06973_);
  and (_06976_, _06975_, _06304_);
  nor (_06977_, _06975_, _06304_);
  nor (_06978_, _06977_, _06976_);
  and (_06979_, _06978_, _06145_);
  nor (_06980_, _06979_, _06972_);
  nor (_06981_, _06355_, _06166_);
  not (_06982_, _06981_);
  and (_06983_, _06649_, _06324_);
  not (_06984_, _06983_);
  nor (_06985_, _06648_, _06337_);
  not (_06986_, _06985_);
  and (_06987_, _06647_, _06332_);
  and (_06988_, _06339_, _06166_);
  nor (_06989_, _06988_, _06987_);
  and (_06990_, _06989_, _06986_);
  and (_06991_, _06990_, _06984_);
  and (_06992_, _06991_, _06982_);
  and (_06993_, _06992_, _06980_);
  nor (_06994_, _06993_, _06967_);
  or (_06995_, _06994_, _06968_);
  and (_05750_, _06995_, _06071_);
  not (_06996_, _06375_);
  nor (_06997_, _06434_, _06996_);
  and (_06998_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_06999_, _06998_, _06390_);
  or (_07000_, _06999_, _06997_);
  or (_07001_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_07002_, _07001_, _06071_);
  and (_05935_, _07002_, _07000_);
  and (_07003_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _06071_);
  not (_07004_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_07005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_07006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_07007_, _07006_, _07005_);
  or (_07008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_07009_, _07008_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_07010_, _07009_, _07007_);
  and (_07011_, _07010_, _07004_);
  and (_07012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _06071_);
  and (_07013_, _07012_, _07011_);
  or (_05942_, _07013_, _07003_);
  and (_07014_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_07015_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_07016_, _06939_);
  not (_07017_, _06934_);
  and (_07018_, _06885_, _06303_);
  not (_07019_, _07018_);
  nand (_07020_, _07019_, _06935_);
  or (_07021_, _06935_, _06276_);
  and (_07022_, _07021_, _07020_);
  nand (_07023_, _07022_, _07017_);
  or (_07024_, _07018_, _07017_);
  and (_07025_, _07024_, _07023_);
  and (_07026_, _07025_, _07016_);
  or (_07027_, _06871_, _06113_);
  or (_07028_, _06880_, _06276_);
  or (_07029_, _07028_, _07027_);
  nand (_07030_, _07028_, _07027_);
  and (_07031_, _07030_, _07029_);
  not (_07032_, _07031_);
  or (_07033_, _07032_, _07021_);
  or (_07034_, _07032_, _07023_);
  nand (_07035_, _07032_, _07023_);
  nand (_07036_, _07035_, _07034_);
  nand (_07037_, _07036_, _07021_);
  and (_07038_, _07037_, _07033_);
  nand (_07039_, _07038_, _07026_);
  or (_07040_, _07038_, _07026_);
  and (_07041_, _07040_, _07039_);
  nand (_07042_, _07024_, _07023_);
  or (_07043_, _07042_, _06942_);
  not (_07044_, _06945_);
  and (_07045_, _06942_, _06939_);
  nand (_07046_, _07045_, _07042_);
  or (_07047_, _07045_, _07042_);
  and (_07048_, _07047_, _07046_);
  nand (_07049_, _07048_, _07044_);
  nand (_07050_, _07049_, _07043_);
  nand (_07051_, _07050_, _07041_);
  nand (_07053_, _07051_, _07039_);
  and (_07054_, _06883_, _06776_);
  and (_07055_, _07054_, _07019_);
  and (_07056_, _07033_, _07034_);
  not (_07057_, _07056_);
  nand (_07058_, _07057_, _07055_);
  or (_07059_, _07057_, _07055_);
  and (_07060_, _07059_, _07058_);
  nand (_07061_, _07060_, _07053_);
  and (_07062_, _07058_, _07029_);
  nand (_07063_, _07062_, _07061_);
  nand (_07064_, _07063_, _07015_);
  or (_07065_, _07063_, _07015_);
  nand (_07067_, _07065_, _07064_);
  and (_07068_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_07070_, _07060_, _07053_);
  and (_07071_, _07070_, _07061_);
  nand (_07073_, _07071_, _07068_);
  and (_07075_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or (_07076_, _07050_, _07041_);
  and (_07078_, _07076_, _07051_);
  nand (_07079_, _07078_, _07075_);
  or (_07081_, _07078_, _07075_);
  nand (_07083_, _07081_, _07079_);
  and (_07084_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_07085_, _07048_, _07044_);
  and (_07086_, _07085_, _07049_);
  nand (_07087_, _07086_, _07084_);
  or (_07088_, _07086_, _07084_);
  nand (_07089_, _07088_, _07087_);
  and (_07090_, _06952_, _06948_);
  or (_07091_, _07090_, _07089_);
  and (_07092_, _07091_, _07087_);
  or (_07093_, _07092_, _07083_);
  and (_07094_, _07093_, _07079_);
  or (_07095_, _07071_, _07068_);
  nand (_07096_, _07095_, _07073_);
  or (_07097_, _07096_, _07094_);
  and (_07098_, _07097_, _07073_);
  or (_07099_, _07098_, _07067_);
  nand (_07100_, _07099_, _07064_);
  nand (_07101_, _07100_, _07014_);
  or (_07102_, _07100_, _07014_);
  and (_07103_, _07102_, _07101_);
  and (_05974_, _07103_, _06071_);
  and (_07104_, _06026_, _06012_);
  and (_07105_, _06804_, _05981_);
  and (_07106_, _06840_, _07105_);
  nand (_07107_, _07106_, _07104_);
  and (_07108_, _06331_, _06321_);
  and (_07109_, _06625_, _06138_);
  nor (_07110_, _07109_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_07112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07113_, _06634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_07114_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07115_, _06623_, _07114_);
  nand (_07116_, _07115_, _07113_);
  or (_07117_, _06593_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07118_, _06138_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07119_, _07118_, _07117_);
  and (_07120_, _07119_, _07116_);
  or (_07121_, _06701_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07122_, _06593_, _07114_);
  nand (_07123_, _07122_, _07121_);
  or (_07124_, _06408_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07126_, _06634_, _07114_);
  nand (_07127_, _07126_, _07124_);
  and (_07128_, _07127_, _07123_);
  nand (_07129_, _07128_, _07120_);
  and (_07130_, _07129_, _07112_);
  nor (_07132_, _07130_, _07110_);
  or (_07133_, _06666_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07134_, _06701_, _07114_);
  nand (_07135_, _07134_, _07133_);
  and (_07136_, _07135_, _07112_);
  and (_07137_, _07119_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07138_, _07137_, _07136_);
  nor (_07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07140_, _07139_, _06113_);
  nor (_07141_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_07142_, _07141_);
  and (_07143_, _07142_, _07140_);
  not (_07144_, _07143_);
  or (_07145_, _06674_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07146_, _06408_, _07114_);
  and (_07147_, _07146_, _07145_);
  or (_07148_, _07147_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07149_, _07116_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07150_, _07149_, _07148_);
  or (_07151_, _07150_, _07144_);
  nor (_07152_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_07153_, _07152_);
  nand (_07154_, _07139_, _06276_);
  and (_07155_, _07154_, _07153_);
  not (_07156_, _07155_);
  and (_07157_, _06666_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07158_, _07157_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07159_, _07123_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07160_, _07159_, _07158_);
  or (_07161_, _07160_, _07156_);
  nand (_07162_, _07149_, _07148_);
  or (_07163_, _07162_, _07143_);
  and (_07164_, _07163_, _07151_);
  not (_07165_, _07164_);
  or (_07166_, _07165_, _07161_);
  and (_07167_, _07166_, _07151_);
  nand (_07168_, _07159_, _07158_);
  or (_07169_, _07168_, _07155_);
  and (_07170_, _07169_, _07161_);
  and (_07171_, _07170_, _07164_);
  not (_07172_, _07139_);
  or (_07173_, _07172_, _06297_);
  nor (_07174_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_07175_, _07174_);
  nand (_07176_, _07175_, _07173_);
  and (_07177_, _06674_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07178_, _07177_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07179_, _07127_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07180_, _07179_, _07178_);
  or (_07181_, _07180_, _07176_);
  nor (_07182_, _07135_, _07112_);
  nor (_07183_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_07184_, _07183_);
  nand (_07185_, _07139_, _06166_);
  and (_07186_, _07185_, _07184_);
  not (_07187_, _07186_);
  or (_07188_, _07187_, _07182_);
  and (_07189_, _07175_, _07173_);
  nand (_07190_, _07179_, _07178_);
  or (_07191_, _07190_, _07189_);
  nand (_07192_, _07191_, _07181_);
  or (_07193_, _07192_, _07188_);
  nand (_07194_, _07193_, _07181_);
  nand (_07195_, _07194_, _07171_);
  and (_07196_, _07195_, _07167_);
  and (_07197_, _07147_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07198_, _07197_);
  nor (_07199_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_07200_, _07199_);
  nand (_07201_, _07139_, _06187_);
  and (_07202_, _07201_, _07200_);
  nand (_07203_, _07202_, _07198_);
  or (_07204_, _07202_, _07198_);
  nand (_07205_, _07204_, _07203_);
  nand (_07206_, _07157_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07207_, _07172_, _06251_);
  nor (_07208_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_07209_, _07208_);
  and (_07210_, _07209_, _07207_);
  nand (_07211_, _07210_, _07206_);
  and (_07212_, _07177_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07213_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_07214_, _07213_);
  or (_07215_, _07172_, _06230_);
  nand (_07216_, _07215_, _07214_);
  and (_07217_, _07216_, _07212_);
  or (_07218_, _07210_, _07206_);
  nand (_07219_, _07218_, _07211_);
  or (_07220_, _07219_, _07217_);
  and (_07221_, _07220_, _07211_);
  or (_07222_, _07221_, _07205_);
  nand (_07223_, _07222_, _07203_);
  not (_07224_, _07182_);
  or (_07225_, _07186_, _07224_);
  and (_07226_, _07225_, _07188_);
  and (_07227_, _07191_, _07181_);
  and (_07228_, _07227_, _07226_);
  and (_07229_, _07228_, _07171_);
  nand (_07230_, _07229_, _07223_);
  nand (_07231_, _07230_, _07196_);
  not (_07232_, _07138_);
  and (_07233_, _07232_, _07132_);
  nand (_07235_, _07233_, _07231_);
  and (_07236_, _07235_, _07143_);
  not (_07237_, _07236_);
  and (_07239_, _07233_, _07231_);
  and (_07240_, _07180_, _07176_);
  not (_07241_, _07188_);
  and (_07242_, _07226_, _07223_);
  nor (_07243_, _07242_, _07241_);
  or (_07244_, _07243_, _07240_);
  and (_07245_, _07244_, _07181_);
  not (_07246_, _07245_);
  nand (_07247_, _07246_, _07170_);
  and (_07248_, _07247_, _07161_);
  nand (_07249_, _07248_, _07164_);
  or (_07250_, _07248_, _07164_);
  nand (_07251_, _07250_, _07249_);
  nand (_07252_, _07251_, _07239_);
  and (_07253_, _07252_, _07237_);
  or (_07254_, _07253_, _07138_);
  or (_07255_, _07246_, _07170_);
  nand (_07256_, _07255_, _07247_);
  nand (_07257_, _07256_, _07239_);
  and (_07259_, _07235_, _07156_);
  not (_07261_, _07259_);
  and (_07262_, _07261_, _07257_);
  nand (_07263_, _07262_, _07162_);
  nand (_07264_, _07253_, _07138_);
  nand (_07265_, _07264_, _07254_);
  or (_07266_, _07265_, _07263_);
  and (_07267_, _07266_, _07254_);
  and (_07268_, _07264_, _07254_);
  or (_07269_, _07262_, _07162_);
  and (_07270_, _07269_, _07263_);
  and (_07271_, _07270_, _07268_);
  nand (_07272_, _07192_, _07243_);
  or (_07273_, _07192_, _07243_);
  nand (_07274_, _07273_, _07272_);
  nand (_07275_, _07274_, _07239_);
  and (_07276_, _07235_, _07176_);
  not (_07277_, _07276_);
  and (_07278_, _07277_, _07275_);
  and (_07279_, _07278_, _07168_);
  nor (_07280_, _07226_, _07223_);
  or (_07281_, _07280_, _07242_);
  and (_07282_, _07281_, _07239_);
  and (_07283_, _07235_, _07187_);
  nor (_07284_, _07283_, _07282_);
  and (_07285_, _07284_, _07190_);
  nor (_07286_, _07278_, _07168_);
  or (_07287_, _07286_, _07279_);
  not (_07288_, _07287_);
  and (_07289_, _07288_, _07285_);
  nor (_07290_, _07289_, _07279_);
  and (_07291_, _07221_, _07205_);
  not (_07292_, _07291_);
  and (_07293_, _07292_, _07222_);
  or (_07294_, _07293_, _07235_);
  or (_07295_, _07239_, _07202_);
  and (_07296_, _07295_, _07294_);
  nor (_07297_, _07296_, _07224_);
  not (_07298_, _07297_);
  not (_07299_, _07212_);
  or (_07300_, _07235_, _07299_);
  nand (_07301_, _07300_, _07216_);
  or (_07302_, _07300_, _07216_);
  and (_07303_, _07302_, _07301_);
  nand (_07304_, _07303_, _07206_);
  or (_07305_, _07303_, _07206_);
  and (_07306_, _07305_, _07304_);
  and (_07307_, _07139_, _06209_);
  nor (_07308_, _07139_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_07309_, _07308_, _07307_);
  nor (_07310_, _07309_, _07299_);
  not (_07311_, _07310_);
  nand (_07312_, _07311_, _07306_);
  nand (_07313_, _07312_, _07304_);
  and (_07314_, _07219_, _07217_);
  not (_07315_, _07314_);
  and (_07316_, _07315_, _07220_);
  or (_07317_, _07316_, _07235_);
  or (_07318_, _07239_, _07210_);
  and (_07319_, _07318_, _07317_);
  nand (_07320_, _07319_, _07198_);
  or (_07321_, _07319_, _07198_);
  and (_07322_, _07321_, _07320_);
  nand (_07323_, _07322_, _07313_);
  and (_07324_, _07296_, _07224_);
  not (_07325_, _07324_);
  and (_07326_, _07325_, _07320_);
  nand (_07327_, _07326_, _07323_);
  and (_07328_, _07327_, _07298_);
  nor (_07329_, _07284_, _07190_);
  nor (_07330_, _07329_, _07285_);
  and (_07331_, _07288_, _07330_);
  nand (_07332_, _07331_, _07328_);
  nand (_07333_, _07332_, _07290_);
  nand (_07334_, _07333_, _07271_);
  nand (_07335_, _07334_, _07267_);
  and (_07336_, _07335_, _07132_);
  nand (_07337_, _07333_, _07270_);
  or (_07338_, _07333_, _07270_);
  nand (_07339_, _07338_, _07337_);
  nand (_07340_, _07339_, _07336_);
  or (_07341_, _07336_, _07262_);
  and (_07342_, _07341_, _07340_);
  nand (_07343_, _07342_, _07108_);
  and (_07344_, _06344_, _06124_);
  and (_07345_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not (_07346_, _07345_);
  or (_07347_, _07073_, _07067_);
  nand (_07348_, _07347_, _07064_);
  and (_07349_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_07350_, _07349_, _07014_);
  and (_07351_, _07350_, _07348_);
  nor (_07352_, _07096_, _07067_);
  nand (_07353_, _07350_, _07352_);
  nor (_07354_, _07353_, _07094_);
  or (_07355_, _07354_, _07351_);
  and (_07356_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  not (_07357_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_07358_, _06853_, _07357_);
  and (_07360_, _07358_, _07356_);
  and (_07361_, _07360_, _07355_);
  and (_07362_, _07361_, _07346_);
  nand (_07363_, _07360_, _07355_);
  and (_07364_, _07363_, _07345_);
  or (_07365_, _07364_, _07362_);
  nand (_07366_, _07365_, _07344_);
  nor (_07367_, _06708_, _06642_);
  nor (_07368_, _07367_, _06709_);
  nor (_07369_, _07368_, _06616_);
  not (_07370_, _07369_);
  nor (_07371_, _06743_, _06737_);
  nor (_07372_, _07371_, _06716_);
  and (_07373_, _07372_, _06745_);
  not (_07374_, _06756_);
  nor (_07375_, _06623_, _06120_);
  nor (_07376_, _07375_, _06128_);
  and (_07377_, _07376_, _07374_);
  and (_07378_, _06311_, _06120_);
  nor (_07379_, _06297_, _06120_);
  and (_07380_, _07379_, _06255_);
  nor (_07381_, _07380_, _07378_);
  nor (_07383_, _07381_, _06276_);
  not (_07384_, _07383_);
  and (_07385_, _07381_, _06276_);
  nor (_07386_, _07385_, _06585_);
  and (_07387_, _07386_, _07384_);
  nor (_07388_, _07387_, _07377_);
  nor (_07389_, _06299_, _06113_);
  not (_07390_, _07389_);
  and (_07391_, _06767_, _07390_);
  not (_07392_, _07391_);
  and (_07393_, _06754_, _06297_);
  nor (_07394_, _07393_, _06303_);
  nor (_07395_, _07394_, _07392_);
  not (_07396_, _07395_);
  and (_07397_, _07392_, _06760_);
  nor (_07398_, _07391_, _06755_);
  and (_07399_, _07398_, _06303_);
  nor (_07400_, _07399_, _07397_);
  and (_07401_, _07400_, _07396_);
  nor (_07402_, _07401_, _06759_);
  and (_07403_, _06628_, _06324_);
  and (_07404_, _06626_, _06332_);
  nor (_07405_, _06627_, _06337_);
  and (_07406_, _06339_, _06276_);
  or (_07407_, _07406_, _07405_);
  or (_07409_, _07407_, _07404_);
  nor (_07410_, _07409_, _07403_);
  not (_07411_, _06350_);
  or (_07412_, _07411_, _06113_);
  and (_07413_, _06352_, _06297_);
  and (_07414_, _06349_, _06303_);
  nor (_07415_, _07414_, _07413_);
  and (_07416_, _07415_, _07412_);
  and (_07417_, _07416_, _07410_);
  not (_07418_, _07417_);
  nor (_07419_, _07418_, _07402_);
  and (_07420_, _07419_, _07388_);
  not (_07421_, _07420_);
  nor (_07422_, _07421_, _07373_);
  and (_07423_, _07422_, _07370_);
  and (_07424_, _07423_, _07366_);
  nand (_07425_, _07424_, _07343_);
  not (_07426_, _07425_);
  nor (_07427_, _07426_, _07107_);
  and (_07428_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05686_);
  and (_07429_, _07428_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_07430_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_07431_, _07430_, _07429_);
  or (_07432_, _07431_, _07427_);
  not (_07433_, _07429_);
  and (_07434_, _06623_, _06349_);
  and (_07435_, _06777_, _06251_);
  and (_07437_, _06646_, _06120_);
  not (_07438_, _07437_);
  nor (_07439_, _06690_, _06113_);
  and (_07440_, _07439_, _06312_);
  and (_07441_, _07440_, _06666_);
  and (_07442_, _07441_, _06408_);
  and (_07443_, _07442_, _06701_);
  or (_07444_, _07443_, _06302_);
  and (_07445_, _07444_, _07438_);
  and (_07446_, _06300_, _06113_);
  and (_07447_, _06690_, _06677_);
  and (_07448_, _06655_, _06660_);
  and (_07449_, _07448_, _07447_);
  and (_07450_, _07449_, _07446_);
  nor (_07451_, _07450_, _06120_);
  not (_07452_, _07451_);
  and (_07453_, _06577_, _06120_);
  and (_07454_, _06646_, _06577_);
  nor (_07455_, _07454_, _06120_);
  nor (_07456_, _07455_, _07453_);
  and (_07457_, _07456_, _07452_);
  and (_07458_, _07457_, _07445_);
  and (_07459_, _07458_, _06623_);
  nor (_07460_, _07458_, _06623_);
  nor (_07461_, _07460_, _07459_);
  and (_07462_, _07461_, _06145_);
  and (_07463_, _06623_, _06120_);
  nor (_07464_, _06276_, _06120_);
  or (_07465_, _07464_, _07463_);
  and (_07466_, _07465_, _06127_);
  or (_07467_, _07466_, _07462_);
  or (_07468_, _07467_, _07435_);
  and (_07469_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_07470_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07471_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06284_);
  nor (_07473_, _07471_, _07470_);
  not (_07474_, _07473_);
  nor (_07475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07477_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06172_);
  nor (_07478_, _07477_, _07475_);
  not (_07479_, _07478_);
  nor (_07480_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_07481_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06193_);
  nor (_07483_, _07481_, _07480_);
  not (_07484_, _07483_);
  nor (_07486_, _07484_, _06749_);
  nor (_07487_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_07488_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06210_);
  nor (_07489_, _07488_, _07487_);
  and (_07490_, _07489_, _07486_);
  nor (_07491_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07492_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06243_);
  nor (_07493_, _07492_, _07491_);
  nand (_07494_, _07493_, _07490_);
  or (_07495_, _07494_, _07479_);
  nor (_07496_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_07497_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06151_);
  nor (_07498_, _07497_, _07496_);
  not (_07499_, _07498_);
  or (_07500_, _07499_, _07495_);
  or (_07501_, _07500_, _07474_);
  nor (_07502_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_07503_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06261_);
  nor (_07504_, _07503_, _07502_);
  not (_07505_, _07504_);
  and (_07506_, _07505_, _07501_);
  not (_07507_, _07506_);
  nor (_07508_, _07505_, _07501_);
  nor (_07509_, _07508_, _06716_);
  and (_07511_, _07509_, _07507_);
  and (_07512_, _07090_, _07089_);
  not (_07514_, _07512_);
  and (_07515_, _07514_, _07091_);
  and (_07516_, _07515_, _07344_);
  or (_07517_, _07516_, _07511_);
  or (_07518_, _07517_, _07469_);
  or (_07519_, _07518_, _07468_);
  or (_07520_, _07519_, _07434_);
  or (_07521_, _07520_, _07433_);
  and (_07523_, _07521_, _06071_);
  and (_06034_, _07523_, _07432_);
  and (_07525_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_07526_, _06804_, _06371_);
  and (_07527_, _07526_, _06840_);
  and (_07528_, _07527_, _06814_);
  and (_07530_, _07528_, _06009_);
  nand (_07531_, _07335_, _07132_);
  or (_07532_, _07322_, _07313_);
  and (_07533_, _07532_, _07323_);
  or (_07534_, _07533_, _07531_);
  or (_07535_, _07336_, _07319_);
  and (_07536_, _07535_, _07534_);
  and (_07537_, _07536_, _07108_);
  and (_07538_, _07103_, _07344_);
  or (_07540_, _06729_, _06727_);
  nor (_07541_, _06730_, _06716_);
  and (_07542_, _07541_, _07540_);
  and (_07543_, _06697_, _06687_);
  or (_07544_, _07543_, _06698_);
  and (_07545_, _07544_, _06615_);
  and (_07546_, _06252_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07547_, _06752_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07548_, _07547_, _06230_);
  nor (_07549_, _07548_, _06429_);
  or (_07550_, _07549_, _07546_);
  and (_07551_, _07550_, _06751_);
  nor (_07552_, _07411_, _06187_);
  and (_07553_, _06349_, _06251_);
  and (_07554_, _06352_, _06230_);
  or (_07555_, _07554_, _07553_);
  nor (_07556_, _07555_, _07552_);
  and (_07557_, _07556_, _06428_);
  and (_07558_, _07557_, _06424_);
  nand (_07559_, _07558_, _06418_);
  or (_07560_, _07559_, _07551_);
  or (_07561_, _07560_, _07545_);
  or (_07562_, _07561_, _07542_);
  or (_07563_, _07562_, _07538_);
  or (_07564_, _07563_, _07537_);
  and (_07565_, _07564_, _07530_);
  or (_07566_, _07565_, _07525_);
  or (_07567_, _07566_, _07429_);
  or (_07569_, _07493_, _07490_);
  and (_07570_, _07494_, _06715_);
  and (_07571_, _07570_, _07569_);
  nor (_07572_, _07441_, _06302_);
  and (_07573_, _07447_, _07446_);
  nor (_07574_, _07573_, _06120_);
  nor (_07575_, _07574_, _07572_);
  nand (_07576_, _07575_, _06408_);
  or (_07577_, _07575_, _06408_);
  and (_07578_, _07577_, _06145_);
  and (_07579_, _07578_, _07576_);
  or (_07580_, _06919_, _06917_);
  and (_07581_, _07580_, _06920_);
  and (_07583_, _07581_, _07344_);
  and (_07584_, _06777_, _06303_);
  and (_07585_, _06251_, _06127_);
  and (_07586_, _06408_, _06349_);
  and (_07587_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_07588_, _07587_, _07586_);
  or (_07590_, _07588_, _07585_);
  or (_07591_, _07590_, _07584_);
  or (_07592_, _07591_, _07583_);
  or (_07593_, _07592_, _07579_);
  or (_07594_, _07593_, _07571_);
  or (_07595_, _07594_, _07433_);
  and (_07596_, _07595_, _06071_);
  and (_06049_, _07596_, _07567_);
  and (_07597_, _07330_, _07328_);
  nor (_07598_, _07597_, _07285_);
  nand (_07599_, _07287_, _07598_);
  or (_07600_, _07287_, _07598_);
  nand (_07601_, _07600_, _07599_);
  nand (_07602_, _07601_, _07336_);
  or (_07603_, _07336_, _07278_);
  and (_07604_, _07603_, _07602_);
  nand (_07605_, _07604_, _07108_);
  nand (_07606_, _07356_, _07355_);
  nor (_07607_, _07358_, _07606_);
  and (_07608_, _07358_, _07606_);
  or (_07609_, _07608_, _07607_);
  nand (_07610_, _07609_, _07344_);
  nor (_07611_, _06707_, _06645_);
  nor (_07612_, _07611_, _06708_);
  nor (_07613_, _07612_, _06616_);
  not (_07614_, _07613_);
  nor (_07615_, _06647_, _06596_);
  or (_07616_, _07615_, _06739_);
  not (_07617_, _07616_);
  nor (_07618_, _07617_, _06736_);
  or (_07619_, _07618_, _06716_);
  nor (_07621_, _07619_, _06737_);
  nor (_07622_, _07393_, _06755_);
  nor (_07623_, _07622_, _07392_);
  and (_07624_, _07622_, _07392_);
  or (_07625_, _07624_, _06759_);
  nor (_07626_, _07625_, _07623_);
  and (_07627_, _06349_, _06297_);
  not (_07628_, _07627_);
  nor (_07630_, _06353_, _06166_);
  nor (_07631_, _07411_, _06276_);
  nor (_07632_, _07631_, _07630_);
  and (_07633_, _07632_, _07628_);
  and (_07634_, _07633_, _06607_);
  not (_07635_, _07634_);
  nor (_07636_, _07635_, _07626_);
  and (_07637_, _07636_, _06590_);
  not (_07638_, _07637_);
  nor (_07639_, _07638_, _07621_);
  and (_07641_, _07639_, _07614_);
  and (_07642_, _07641_, _07610_);
  and (_07643_, _07642_, _07605_);
  nor (_07644_, _07643_, _07107_);
  and (_07645_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_07646_, _07645_, _07429_);
  or (_07647_, _07646_, _07644_);
  and (_07648_, _06593_, _06349_);
  and (_07650_, _06777_, _06230_);
  and (_07651_, _07450_, _06646_);
  nor (_07652_, _07651_, _06120_);
  not (_07653_, _07652_);
  and (_07654_, _07653_, _07445_);
  and (_07655_, _07654_, _06577_);
  nor (_07656_, _07654_, _06577_);
  nor (_07657_, _07656_, _07655_);
  nor (_07658_, _07657_, _06585_);
  not (_07659_, _07379_);
  nor (_07660_, _07453_, _06128_);
  and (_07661_, _07660_, _07659_);
  or (_07662_, _07661_, _07658_);
  or (_07663_, _07662_, _07650_);
  and (_07664_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  and (_07665_, _07500_, _07474_);
  not (_07666_, _07665_);
  and (_07667_, _07501_, _06715_);
  and (_07668_, _07667_, _07666_);
  and (_07669_, _06956_, _07344_);
  or (_07670_, _07669_, _07668_);
  or (_07671_, _07670_, _07664_);
  or (_07672_, _07671_, _07663_);
  nor (_07673_, _07672_, _07648_);
  nand (_07674_, _07673_, _07429_);
  and (_07675_, _07674_, _06071_);
  and (_06052_, _07675_, _07647_);
  and (_06060_, _07609_, _06071_);
  nor (_07676_, _07330_, _07328_);
  or (_07677_, _07676_, _07597_);
  nand (_07678_, _07677_, _07336_);
  or (_07679_, _07336_, _07284_);
  and (_07680_, _07679_, _07678_);
  nand (_07681_, _07680_, _07108_);
  or (_07682_, _07356_, _07355_);
  and (_07683_, _07682_, _07606_);
  nand (_07684_, _07683_, _07344_);
  nor (_07685_, _06706_, _06649_);
  and (_07686_, _06706_, _06649_);
  nor (_07687_, _07686_, _07685_);
  and (_07688_, _07687_, _06615_);
  not (_07689_, _07688_);
  nor (_07690_, _06735_, _06649_);
  not (_07691_, _07690_);
  nor (_07692_, _06736_, _06716_);
  and (_07693_, _07692_, _07691_);
  and (_07694_, _06753_, _06166_);
  not (_07695_, _07694_);
  nor (_07696_, _06752_, _06759_);
  and (_07697_, _07696_, _06304_);
  not (_07698_, _07697_);
  nor (_07699_, _06353_, _06187_);
  not (_07700_, _07699_);
  nand (_07701_, _06350_, _06297_);
  not (_07702_, _07701_);
  and (_07703_, _06349_, _06304_);
  nor (_07704_, _07703_, _07702_);
  and (_07705_, _07704_, _07700_);
  and (_07706_, _07705_, _07698_);
  and (_07707_, _07706_, _07695_);
  and (_07709_, _07707_, _06991_);
  and (_07710_, _07709_, _06980_);
  not (_07711_, _07710_);
  nor (_07712_, _07711_, _07693_);
  and (_07713_, _07712_, _07689_);
  and (_07714_, _07713_, _07684_);
  and (_07715_, _07714_, _07681_);
  nor (_07716_, _07715_, _07107_);
  and (_07717_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_07718_, _07717_, _07429_);
  or (_07719_, _07718_, _07716_);
  and (_07720_, _06634_, _06349_);
  and (_07721_, _06777_, _06306_);
  and (_07722_, _07452_, _07444_);
  nor (_07723_, _07722_, _06634_);
  and (_07724_, _07722_, _06634_);
  or (_07725_, _07724_, _06585_);
  nor (_07726_, _07725_, _07723_);
  and (_07727_, _06166_, _06302_);
  not (_07728_, _07727_);
  nor (_07729_, _07437_, _06128_);
  and (_07730_, _07729_, _07728_);
  or (_07731_, _07730_, _07726_);
  or (_07732_, _07731_, _07721_);
  and (_07733_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and (_07734_, _07499_, _07495_);
  not (_07735_, _07734_);
  and (_07737_, _07500_, _06715_);
  and (_07738_, _07737_, _07735_);
  and (_07739_, _06926_, _06924_);
  not (_07740_, _07739_);
  and (_07741_, _07740_, _06927_);
  and (_07742_, _07741_, _07344_);
  or (_07743_, _07742_, _07738_);
  or (_07744_, _07743_, _07733_);
  or (_07745_, _07744_, _07732_);
  nor (_07746_, _07745_, _07720_);
  nand (_07747_, _07746_, _07429_);
  and (_07748_, _07747_, _06071_);
  and (_06063_, _07748_, _07719_);
  and (_06074_, _07683_, _06071_);
  not (_07749_, _07349_);
  and (_07750_, _07749_, _07101_);
  or (_07751_, _07750_, _07355_);
  nor (_06092_, _07751_, rst);
  not (_07752_, _05993_);
  and (_07753_, _06004_, _05981_);
  and (_07754_, _07753_, _07752_);
  and (_07755_, _07104_, _07754_);
  and (_07756_, _07755_, _06840_);
  nor (_07757_, _07756_, _07429_);
  or (_07758_, _07757_, _07564_);
  not (_07759_, _07757_);
  or (_07760_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_07761_, _07760_, _06071_);
  and (_06096_, _07761_, _07758_);
  nand (_07762_, _07759_, _07643_);
  or (_07763_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_07764_, _07763_, _06071_);
  and (_06130_, _07764_, _07762_);
  not (_07765_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_07766_, _07428_, _07765_);
  not (_07767_, _05937_);
  and (_07768_, _07767_, _05923_);
  and (_07769_, _07768_, _05968_);
  and (_07770_, _07769_, _06372_);
  and (_07771_, _07770_, _06012_);
  nor (_07772_, _07771_, _07766_);
  not (_07773_, _07772_);
  or (_07774_, _07336_, _07253_);
  and (_07775_, _07337_, _07263_);
  nand (_07776_, _07775_, _07268_);
  or (_07777_, _07775_, _07268_);
  nand (_07778_, _07777_, _07776_);
  nand (_07779_, _07778_, _07336_);
  nand (_07781_, _07779_, _07774_);
  nand (_07782_, _07781_, _07108_);
  and (_07783_, _06854_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_07784_, _07363_, _07346_);
  nand (_07785_, _07784_, _07783_);
  or (_07786_, _07784_, _07783_);
  nand (_07787_, _07786_, _07785_);
  nand (_07788_, _07787_, _07344_);
  not (_07789_, _06327_);
  and (_07790_, _06710_, _07789_);
  nor (_07791_, _06710_, _07789_);
  nor (_07792_, _07791_, _07790_);
  and (_07793_, _07792_, _06615_);
  not (_07794_, _07793_);
  nor (_07795_, _06747_, _07789_);
  and (_07796_, _06747_, _07789_);
  or (_07797_, _07796_, _07795_);
  nor (_07798_, _07797_, _06716_);
  nor (_07799_, _07391_, _06760_);
  nor (_07800_, _07799_, _06113_);
  and (_07801_, _07799_, _06113_);
  nor (_07802_, _07801_, _07800_);
  nor (_07803_, _07802_, _06759_);
  nor (_07804_, _06353_, _06276_);
  and (_07805_, _06787_, _06302_);
  nor (_07806_, _07805_, _07804_);
  and (_07807_, _06349_, _06776_);
  and (_07808_, _06789_, _06306_);
  nor (_07809_, _07808_, _07807_);
  and (_07810_, _07809_, _07806_);
  and (_07811_, _07810_, _06343_);
  not (_07812_, _07811_);
  nor (_07813_, _07812_, _07803_);
  and (_07814_, _07813_, _06319_);
  not (_07815_, _07814_);
  nor (_07816_, _07815_, _07798_);
  and (_07817_, _07816_, _07794_);
  and (_07818_, _07817_, _07788_);
  nand (_07819_, _07818_, _07782_);
  nand (_07820_, _07819_, _07773_);
  not (_07821_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_07822_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05686_);
  and (_07823_, _07822_, _07821_);
  nor (_07824_, _05954_, _05937_);
  and (_07825_, _07824_, _06833_);
  and (_07826_, _07825_, _06815_);
  and (_07827_, _07826_, _06805_);
  and (_07828_, _07827_, _06803_);
  nor (_07829_, _07827_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_07830_, _07823_);
  and (_07831_, _07830_, _07772_);
  not (_07832_, _07831_);
  nor (_07833_, _07832_, _07829_);
  not (_07834_, _07833_);
  nor (_07835_, _07834_, _07828_);
  nor (_07836_, _07835_, _07823_);
  nand (_07837_, _07836_, _07820_);
  nor (_07838_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_07839_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _06086_);
  nor (_07840_, _07839_, _07838_);
  and (_07841_, _07840_, _07508_);
  nor (_07843_, _07840_, _07508_);
  or (_07844_, _07843_, _06716_);
  or (_07845_, _07844_, _07841_);
  and (_07846_, _07092_, _07083_);
  not (_07847_, _07846_);
  and (_07848_, _07847_, _07093_);
  and (_07849_, _07848_, _07344_);
  nor (_07850_, _07463_, _07375_);
  not (_07851_, _07850_);
  and (_07852_, _07851_, _07458_);
  nor (_07853_, _07852_, _06139_);
  and (_07854_, _07852_, _06139_);
  nor (_07855_, _07854_, _07853_);
  and (_07856_, _07855_, _06145_);
  and (_07857_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_07858_, _06127_, _06120_);
  or (_07859_, _07858_, _06349_);
  and (_07860_, _07859_, _06139_);
  or (_07861_, _07860_, _07857_);
  and (_07862_, _06777_, _06305_);
  and (_07863_, _06761_, _06127_);
  or (_07864_, _07863_, _07862_);
  nor (_07865_, _07864_, _07861_);
  not (_07866_, _07865_);
  nor (_07867_, _07866_, _07856_);
  not (_07868_, _07867_);
  nor (_07869_, _07868_, _07849_);
  nand (_07870_, _07869_, _07845_);
  or (_07871_, _07870_, _07830_);
  and (_07872_, _07871_, _07837_);
  and (_06199_, _07872_, _06071_);
  and (_07873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_07874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_07875_, _07874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_07876_, _07875_);
  nor (_07877_, _07876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not (_07878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_07879_, _07878_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_07880_, _07879_, _07877_);
  nor (_07881_, _07880_, _07873_);
  or (_07882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_07883_, _07882_, _06071_);
  nor (_06346_, _07883_, _07881_);
  and (_07884_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_07886_, _07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_07887_, _07886_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_07888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_07889_, _07885_, _07888_);
  and (_07890_, _07889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_07891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_07892_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _07891_);
  not (_07893_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_07894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _07893_);
  and (_07895_, _07894_, _07892_);
  and (_07896_, _07895_, _07890_);
  nor (_07897_, _07896_, _07887_);
  not (_07898_, _07897_);
  and (_07899_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  not (_07900_, _07890_);
  nor (_07901_, _07895_, _07900_);
  not (_07902_, _07885_);
  and (_07903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_07904_, _07903_, _07902_);
  not (_07905_, _07904_);
  and (_07906_, _07888_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not (_07907_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_07908_, _07885_, _07907_);
  and (_07909_, _07908_, _07906_);
  nor (_07910_, _07909_, _07890_);
  and (_07911_, _07910_, _07905_);
  nor (_07912_, _07911_, _07901_);
  not (_07913_, _07887_);
  nand (_07914_, _07913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_07915_, _07914_, _07912_);
  or (_07916_, _07915_, _07899_);
  and (_07917_, _07916_, _06560_);
  or (_06379_, _07917_, _07884_);
  and (_07918_, _06922_, _06920_);
  not (_07919_, _07918_);
  and (_07920_, _07919_, _06923_);
  and (_06589_, _07920_, _06071_);
  and (_06604_, _07581_, _06071_);
  and (_07922_, _06881_, _06872_);
  nor (_07923_, _07922_, _06882_);
  and (_06606_, _07923_, _06071_);
  and (_07924_, _06885_, _06306_);
  and (_06617_, _07924_, _06071_);
  and (_07925_, _06701_, _06127_);
  nor (_07926_, _06253_, _06120_);
  nor (_07927_, _06308_, _06302_);
  nor (_07928_, _07927_, _07926_);
  and (_07929_, _07928_, _06305_);
  not (_07930_, _07929_);
  nor (_07931_, _07928_, _06305_);
  nor (_07932_, _07931_, _06585_);
  and (_07933_, _07932_, _07930_);
  nor (_07934_, _07933_, _07925_);
  nor (_07935_, _06656_, _06337_);
  and (_07936_, _06659_, _06324_);
  nor (_07937_, _07936_, _07935_);
  and (_07938_, _06657_, _06332_);
  and (_07939_, _06339_, _06187_);
  nor (_07940_, _07939_, _07938_);
  nor (_07941_, _06355_, _06187_);
  not (_07942_, _07941_);
  and (_07943_, _07942_, _07940_);
  and (_07944_, _07943_, _07937_);
  and (_07945_, _07944_, _07934_);
  and (_07946_, _06374_, _06011_);
  nand (_07947_, _07946_, _07945_);
  or (_07948_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_07949_, _07948_, _06071_);
  and (_06658_, _07949_, _07947_);
  and (_07950_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  not (_07951_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_07952_, _07897_, _07951_);
  nand (_07953_, _07913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_07954_, _07953_, _07912_);
  or (_07955_, _07954_, _07952_);
  and (_07956_, _07955_, _06560_);
  or (_06679_, _07956_, _07950_);
  not (_07957_, _06374_);
  nand (_07958_, _06438_, _07957_);
  and (_07959_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_07960_, _06691_, _06332_);
  and (_07961_, _06339_, _06209_);
  nor (_07962_, _07961_, _07960_);
  and (_07963_, _06674_, _06127_);
  and (_07964_, _06145_, _06209_);
  nor (_07965_, _07964_, _07963_);
  nor (_07966_, _07808_, _06788_);
  and (_07967_, _07966_, _07965_);
  and (_07968_, _07967_, _07962_);
  nor (_07969_, _06691_, _06770_);
  nor (_07970_, _07969_, _06336_);
  or (_07971_, _07970_, _06692_);
  nor (_07972_, _06352_, _06349_);
  and (_07973_, _07972_, _06348_);
  nor (_07974_, _07973_, _06209_);
  not (_07975_, _07974_);
  and (_07976_, _07975_, _07971_);
  and (_07977_, _07976_, _07968_);
  not (_07978_, _07977_);
  and (_07979_, _06377_, _06011_);
  and (_07980_, _07979_, _07978_);
  or (_07981_, _06384_, _06362_);
  and (_07983_, _07981_, _06373_);
  and (_07984_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_07985_, _07984_, _07983_);
  or (_07986_, _07985_, _07980_);
  or (_07988_, _07986_, _07959_);
  and (_06778_, _07988_, _06071_);
  and (_07989_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_07990_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_07991_, _07901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_07992_, _07904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_07993_, _07992_, _07910_);
  or (_07994_, _07993_, _07991_);
  and (_07996_, _07994_, _07913_);
  or (_07997_, _07996_, _07990_);
  and (_07998_, _07997_, _06560_);
  or (_06783_, _07998_, _07989_);
  and (_07999_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_08000_, _06993_, _06611_);
  or (_08001_, _08000_, _07999_);
  and (_06811_, _08001_, _06071_);
  and (_08002_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_06909_, _08002_, _07884_);
  and (_06950_, _05768_, _06071_);
  not (_08003_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_08004_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08003_);
  and (_08005_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_08006_, _08005_, _08004_);
  and (_06953_, _08006_, _06071_);
  nor (_08007_, _07344_, _06857_);
  and (_08008_, _07344_, _06857_);
  or (_08009_, _08008_, _08007_);
  and (_07052_, _08009_, _06071_);
  and (_07066_, _05788_, _06071_);
  and (_07069_, _05810_, _06071_);
  and (_07072_, _05829_, _06071_);
  and (_07074_, _05847_, _06071_);
  and (_07077_, _05880_, _06071_);
  and (_07080_, _05726_, _06071_);
  and (_07082_, _05747_, _06071_);
  nor (_08010_, _06609_, _06996_);
  and (_08011_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_08012_, _08011_, _06390_);
  or (_08013_, _08012_, _08010_);
  or (_08014_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_08015_, _08014_, _06071_);
  and (_07111_, _08015_, _08013_);
  and (_08016_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_08018_, _08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_08019_, _08017_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_08020_, _08019_, _08018_);
  or (_08021_, _08020_, _08016_);
  and (_07125_, _08021_, _06071_);
  and (_08022_, _08003_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_08023_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_08024_, _08023_, _08022_);
  and (_07131_, _08024_, _06071_);
  nand (_08025_, _07336_, _07212_);
  and (_08026_, _08025_, _07309_);
  nor (_08027_, _08025_, _07309_);
  or (_08028_, _08027_, _08026_);
  nand (_08029_, _08028_, _07108_);
  not (_08030_, _07097_);
  and (_08031_, _07096_, _07094_);
  nor (_08032_, _08031_, _08030_);
  and (_08033_, _08032_, _07344_);
  and (_08034_, _06350_, _06230_);
  nor (_08035_, _06751_, _06349_);
  nor (_08036_, _08035_, _06209_);
  nor (_08037_, _08036_, _08034_);
  nor (_08038_, _06693_, _06302_);
  nor (_08039_, _08038_, _06726_);
  nor (_08040_, _06715_, _06615_);
  not (_08041_, _08040_);
  and (_08042_, _08041_, _08039_);
  and (_08043_, _06781_, _06776_);
  and (_08044_, _06777_, _06302_);
  nor (_08045_, _08044_, _08043_);
  and (_08046_, _08045_, _07965_);
  nand (_08047_, _08046_, _07962_);
  nor (_08048_, _08047_, _08042_);
  and (_08049_, _08048_, _08037_);
  and (_08050_, _08049_, _07971_);
  not (_08051_, _08050_);
  nor (_08052_, _08051_, _08033_);
  and (_08053_, _08052_, _08029_);
  nand (_08054_, _08053_, _07759_);
  or (_08056_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_08057_, _08056_, _06071_);
  and (_07234_, _08057_, _08054_);
  or (_08058_, _07311_, _07306_);
  and (_08059_, _08058_, _07312_);
  or (_08060_, _08059_, _07531_);
  or (_08061_, _07336_, _07303_);
  and (_08062_, _08061_, _08060_);
  nand (_08063_, _08062_, _07108_);
  nand (_08064_, _07098_, _07067_);
  and (_08065_, _08064_, _07099_);
  nand (_08066_, _08065_, _07344_);
  and (_08067_, _06695_, _06689_);
  nor (_08068_, _08067_, _06696_);
  nor (_08069_, _08068_, _06616_);
  not (_08070_, _08069_);
  and (_08071_, _06666_, _06127_);
  nor (_08072_, _06230_, _06209_);
  and (_08073_, _06230_, _06209_);
  nor (_08074_, _08073_, _08072_);
  nor (_08075_, _08074_, _06302_);
  and (_08076_, _08074_, _06302_);
  nor (_08077_, _08076_, _08075_);
  nor (_08078_, _08077_, _06585_);
  nor (_08079_, _08078_, _08071_);
  nand (_08080_, _06350_, _06251_);
  nor (_08081_, _06353_, _06209_);
  and (_08082_, _06349_, _06230_);
  nor (_08083_, _08082_, _08081_);
  and (_08084_, _08083_, _08080_);
  and (_08086_, _06669_, _06324_);
  nor (_08087_, _06668_, _06337_);
  not (_08088_, _08087_);
  and (_08090_, _06667_, _06332_);
  nor (_08091_, _06426_, _06230_);
  nor (_08092_, _08091_, _08090_);
  nand (_08093_, _08092_, _08088_);
  nor (_08094_, _08093_, _08086_);
  and (_08095_, _08094_, _08084_);
  and (_08096_, _08095_, _08079_);
  and (_08097_, _07547_, _06230_);
  nor (_08098_, _08097_, _07548_);
  nor (_08099_, _08098_, _06759_);
  nor (_08100_, _06691_, _06669_);
  or (_08101_, _08100_, _06719_);
  and (_08102_, _08101_, _06726_);
  nor (_08103_, _08101_, _06726_);
  or (_08104_, _08103_, _08102_);
  and (_08105_, _08104_, _06715_);
  nor (_08106_, _08105_, _08099_);
  and (_08107_, _08106_, _08096_);
  and (_08108_, _08107_, _08070_);
  and (_08109_, _08108_, _08066_);
  and (_08110_, _08109_, _08063_);
  nand (_08111_, _08110_, _07759_);
  or (_08112_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_08113_, _08112_, _06071_);
  and (_07238_, _08113_, _08111_);
  nor (_08114_, _08053_, _07107_);
  and (_08115_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_08116_, _08115_, _07429_);
  or (_08117_, _08116_, _08114_);
  and (_08118_, _07484_, _06749_);
  nor (_08119_, _08118_, _07486_);
  and (_08120_, _08119_, _06715_);
  nand (_08121_, _07336_, _07108_);
  nor (_08122_, _06761_, _06121_);
  not (_08123_, _08122_);
  nor (_08124_, _08123_, _06314_);
  and (_08125_, _08124_, _06674_);
  nor (_08126_, _08124_, _06674_);
  nor (_08127_, _08126_, _08125_);
  and (_08128_, _08127_, _06145_);
  and (_08129_, _06674_, _06349_);
  and (_08130_, _07924_, _07344_);
  and (_08131_, _06777_, _06304_);
  nor (_08132_, _06209_, _06128_);
  or (_08133_, _08132_, _08131_);
  or (_08134_, _08133_, _08130_);
  nor (_08135_, _08134_, _08129_);
  not (_08136_, _08135_);
  nor (_08137_, _08136_, _08128_);
  nand (_08138_, _08137_, _08121_);
  or (_08139_, _08138_, _08120_);
  or (_08140_, _08139_, _07433_);
  and (_08141_, _08140_, _06071_);
  and (_07258_, _08141_, _08117_);
  nor (_08142_, _08110_, _07107_);
  and (_08143_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_08144_, _08143_, _07429_);
  or (_08145_, _08144_, _08142_);
  and (_08146_, _06666_, _06349_);
  and (_08147_, _06777_, _06297_);
  nor (_08148_, _07440_, _06302_);
  and (_08150_, _06690_, _07446_);
  nor (_08151_, _08150_, _06120_);
  or (_08152_, _08151_, _08148_);
  nor (_08153_, _08152_, _06666_);
  and (_08154_, _08152_, _06666_);
  nor (_08155_, _08154_, _08153_);
  nor (_08156_, _08155_, _06585_);
  and (_08158_, _06230_, _06127_);
  or (_08159_, _08158_, _08156_);
  or (_08160_, _08159_, _08147_);
  and (_08161_, _07239_, _07108_);
  nor (_08162_, _07489_, _07486_);
  nor (_08163_, _08162_, _07490_);
  and (_08164_, _08163_, _06715_);
  and (_08165_, _07923_, _07344_);
  or (_08166_, _08165_, _08164_);
  or (_08167_, _08166_, _08161_);
  or (_08168_, _08167_, _08160_);
  nor (_08169_, _08168_, _08146_);
  nand (_08170_, _08169_, _07429_);
  and (_08171_, _08170_, _06071_);
  and (_07260_, _08171_, _08145_);
  nor (_08172_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_08173_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_08174_, _08173_, _08172_);
  not (_08175_, _08174_);
  not (_08176_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_08177_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_08178_, _06530_, _08177_);
  nor (_08179_, _08178_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_08180_, _08178_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08181_, _08180_, _08179_);
  nor (_08182_, _08181_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08183_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_08184_, _08183_, _08182_);
  nor (_08185_, _08184_, _08176_);
  and (_08186_, _08184_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_08187_, _08186_, _08185_);
  nor (_08188_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_08189_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_08190_, _08189_, _08188_);
  and (_08191_, _06530_, _08177_);
  nor (_08192_, _08191_, _08178_);
  nor (_08193_, _08192_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08194_, _08003_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_08195_, _08194_, _08193_);
  nor (_08196_, _08195_, _08190_);
  not (_08197_, _08196_);
  nor (_08198_, _08197_, _08187_);
  or (_08199_, _08198_, _08175_);
  and (_08200_, _08195_, _08190_);
  not (_08201_, _08200_);
  nor (_08202_, _08184_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_08203_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_08204_, _08184_, _08203_);
  or (_08205_, _08204_, _08202_);
  nor (_08206_, _08205_, _08201_);
  not (_08207_, _08190_);
  nor (_08208_, _08195_, _08207_);
  not (_08209_, _08208_);
  not (_08210_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08211_, _08184_, _08210_);
  and (_08212_, _08184_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08213_, _08212_, _08211_);
  nor (_08214_, _08213_, _08209_);
  not (_08215_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_08217_, _08184_, _08215_);
  nor (_08218_, _08184_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08219_, _08218_, _08217_);
  not (_08220_, _08219_);
  and (_08221_, _08195_, _08207_);
  and (_08222_, _08221_, _08220_);
  or (_08223_, _08222_, _08214_);
  or (_08224_, _08223_, _08206_);
  nor (_08225_, _08224_, _08199_);
  nor (_08227_, _08184_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_08228_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08229_, _08184_, _08228_);
  or (_08230_, _08229_, _08227_);
  nor (_08231_, _08230_, _08201_);
  nor (_08232_, _08231_, _08174_);
  not (_08233_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08234_, _08184_, _08233_);
  nor (_08235_, _08184_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08236_, _08235_, _08234_);
  not (_08237_, _08236_);
  nand (_08238_, _08237_, _08221_);
  and (_08239_, _08184_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_08240_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_08241_, _08184_, _08240_);
  nor (_08242_, _08241_, _08239_);
  nor (_08243_, _08242_, _08209_);
  nor (_08244_, _08184_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_08245_, _08244_);
  not (_08246_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08247_, _08184_, _08246_);
  nor (_08248_, _08247_, _08197_);
  and (_08249_, _08248_, _08245_);
  nor (_08250_, _08249_, _08243_);
  and (_08251_, _08250_, _08238_);
  and (_08252_, _08251_, _08232_);
  nor (_08253_, _08252_, _08225_);
  not (_08254_, _08253_);
  and (_08255_, _08254_, word_in[7]);
  not (_08256_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_08257_, _08174_, _08256_);
  or (_08258_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_08259_, _08258_, _08257_);
  and (_08260_, _08259_, _08196_);
  or (_08261_, _08260_, _08184_);
  not (_08262_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08263_, _08174_, _08262_);
  or (_08264_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_08266_, _08264_, _08263_);
  and (_08267_, _08266_, _08221_);
  not (_08268_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08269_, _08174_, _08268_);
  or (_08270_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_08271_, _08270_, _08269_);
  and (_08272_, _08271_, _08200_);
  or (_08273_, _08272_, _08267_);
  not (_08274_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_08275_, _08174_, _08274_);
  or (_08276_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_08277_, _08276_, _08275_);
  and (_08278_, _08277_, _08208_);
  or (_08279_, _08278_, _08273_);
  or (_08280_, _08279_, _08261_);
  not (_08281_, _08184_);
  not (_08282_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_08283_, _08174_, _08282_);
  or (_08284_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_08285_, _08284_, _08283_);
  and (_08286_, _08285_, _08196_);
  or (_08287_, _08286_, _08281_);
  not (_08288_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_08289_, _08174_, _08288_);
  or (_08290_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_08291_, _08290_, _08289_);
  and (_08292_, _08291_, _08221_);
  not (_08293_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_08294_, _08174_, _08293_);
  or (_08295_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_08296_, _08295_, _08294_);
  and (_08297_, _08296_, _08200_);
  or (_08298_, _08297_, _08292_);
  not (_08299_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08300_, _08174_, _08299_);
  or (_08301_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_08302_, _08301_, _08300_);
  and (_08303_, _08302_, _08208_);
  or (_08304_, _08303_, _08298_);
  or (_08305_, _08304_, _08287_);
  and (_08306_, _08305_, _08280_);
  and (_08307_, _08306_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08307_, _08255_);
  and (_08308_, _08207_, _08174_);
  not (_08309_, _08308_);
  and (_08310_, _08190_, _08174_);
  and (_08311_, _08310_, _08195_);
  nor (_08312_, _08310_, _08195_);
  nor (_08313_, _08312_, _08311_);
  not (_08314_, _08313_);
  nor (_08315_, _08314_, _08230_);
  nor (_08316_, _08311_, _08281_);
  not (_08317_, _08195_);
  nor (_08318_, _08317_, _08184_);
  and (_08319_, _08310_, _08318_);
  nor (_08320_, _08319_, _08316_);
  and (_08321_, _08320_, _08314_);
  and (_08322_, _08321_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_08323_, _08320_, _08313_);
  and (_08324_, _08323_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08325_, _08324_, _08322_);
  nor (_08326_, _08325_, _08315_);
  nor (_08327_, _08326_, _08309_);
  nor (_08328_, _08190_, _08174_);
  not (_08329_, _08328_);
  nor (_08330_, _08314_, _08219_);
  and (_08331_, _08321_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08332_, _08323_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08333_, _08332_, _08331_);
  nor (_08334_, _08333_, _08330_);
  nor (_08335_, _08334_, _08329_);
  nor (_08336_, _08335_, _08327_);
  not (_08337_, _08310_);
  nor (_08338_, _08314_, _08236_);
  and (_08339_, _08321_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_08340_, _08323_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08341_, _08340_, _08339_);
  nor (_08342_, _08341_, _08338_);
  nor (_08343_, _08342_, _08337_);
  and (_08344_, _08190_, _08175_);
  not (_08345_, _08344_);
  and (_08346_, _08313_, _08281_);
  and (_08347_, _08346_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08348_, _08323_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08349_, _08321_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_08350_, _08313_, _08184_);
  and (_08351_, _08350_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_08352_, _08351_, _08349_);
  or (_08353_, _08352_, _08348_);
  nor (_08354_, _08353_, _08347_);
  nor (_08355_, _08354_, _08345_);
  nor (_08356_, _08355_, _08343_);
  and (_08357_, _08356_, _08336_);
  or (_08358_, _08328_, _08310_);
  not (_08359_, _08358_);
  not (_08360_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_08361_, _08174_, _08360_);
  or (_08362_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_08363_, _08362_, _08361_);
  and (_08364_, _08363_, _08359_);
  not (_08365_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_08366_, _08174_, _08365_);
  or (_08367_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_08368_, _08367_, _08366_);
  and (_08369_, _08368_, _08358_);
  or (_08370_, _08369_, _08364_);
  and (_08371_, _08370_, _08323_);
  not (_08372_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_08373_, _08174_, _08372_);
  or (_08374_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_08375_, _08374_, _08373_);
  and (_08376_, _08375_, _08359_);
  not (_08377_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_08378_, _08174_, _08377_);
  or (_08379_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_08380_, _08379_, _08378_);
  and (_08381_, _08380_, _08358_);
  or (_08382_, _08381_, _08376_);
  and (_08383_, _08382_, _08321_);
  not (_08384_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08386_, _08174_, _08384_);
  or (_08387_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_08388_, _08387_, _08386_);
  and (_08389_, _08388_, _08359_);
  not (_08390_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_08391_, _08174_, _08390_);
  or (_08392_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_08393_, _08392_, _08391_);
  and (_08394_, _08393_, _08358_);
  or (_08395_, _08394_, _08389_);
  and (_08396_, _08395_, _08346_);
  not (_08397_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_08398_, _08174_, _08397_);
  or (_08399_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_08400_, _08399_, _08398_);
  and (_08401_, _08400_, _08359_);
  not (_08402_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08403_, _08174_, _08402_);
  or (_08404_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_08405_, _08404_, _08403_);
  and (_08406_, _08405_, _08358_);
  or (_08407_, _08406_, _08401_);
  and (_08408_, _08407_, _08350_);
  or (_08409_, _08408_, _08396_);
  or (_08410_, _08409_, _08383_);
  nor (_08411_, _08410_, _08371_);
  nor (_08412_, _08411_, _08357_);
  and (_08413_, _08357_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08413_, _08412_);
  nor (_08414_, _08200_, _08196_);
  not (_08415_, _08414_);
  nor (_08416_, _08415_, _08205_);
  and (_08417_, _08200_, _08184_);
  nor (_08418_, _08200_, _08184_);
  nor (_08419_, _08418_, _08417_);
  and (_08420_, _08415_, _08419_);
  and (_08421_, _08420_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08422_, _08414_, _08419_);
  and (_08423_, _08422_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08424_, _08423_, _08421_);
  nor (_08425_, _08424_, _08416_);
  nor (_08426_, _08425_, _08309_);
  not (_08427_, _08426_);
  and (_08428_, _08344_, _08318_);
  nand (_08429_, _08428_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08430_, _08415_, _08236_);
  and (_08431_, _08422_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08432_, _08431_, _08430_);
  or (_08433_, _08432_, _08345_);
  and (_08434_, _08433_, _08429_);
  and (_08435_, _08434_, _08427_);
  nor (_08436_, _08415_, _08230_);
  and (_08437_, _08420_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08438_, _08422_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08439_, _08438_, _08437_);
  nor (_08440_, _08439_, _08436_);
  nor (_08441_, _08440_, _08329_);
  nor (_08442_, _08415_, _08219_);
  and (_08443_, _08420_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08444_, _08422_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08445_, _08444_, _08443_);
  nor (_08446_, _08445_, _08442_);
  nor (_08448_, _08446_, _08337_);
  nor (_08449_, _08448_, _08441_);
  and (_08450_, _08449_, _08435_);
  and (_08451_, _08450_, word_in[23]);
  and (_08452_, _08266_, _08208_);
  and (_08453_, _08277_, _08196_);
  or (_08454_, _08453_, _08452_);
  and (_08455_, _08271_, _08221_);
  and (_08456_, _08259_, _08200_);
  or (_08457_, _08456_, _08455_);
  or (_08458_, _08457_, _08454_);
  or (_08459_, _08458_, _08419_);
  not (_08460_, _08419_);
  and (_08461_, _08291_, _08208_);
  and (_08462_, _08302_, _08196_);
  or (_08463_, _08462_, _08461_);
  and (_08464_, _08296_, _08221_);
  and (_08465_, _08285_, _08200_);
  or (_08466_, _08465_, _08464_);
  or (_08467_, _08466_, _08463_);
  or (_08468_, _08467_, _08460_);
  nand (_08469_, _08468_, _08459_);
  nor (_08470_, _08469_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08470_, _08451_);
  nor (_08471_, _08329_, _08195_);
  nand (_08472_, _08329_, _08195_);
  not (_08473_, _08472_);
  nor (_08474_, _08473_, _08471_);
  not (_08475_, _08474_);
  nor (_08476_, _08475_, _08236_);
  nor (_08477_, _08472_, _08184_);
  and (_08478_, _08472_, _08184_);
  nor (_08479_, _08478_, _08477_);
  and (_08480_, _08479_, _08475_);
  and (_08481_, _08480_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08482_, _08479_, _08474_);
  and (_08483_, _08482_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08484_, _08483_, _08481_);
  nor (_08485_, _08484_, _08476_);
  nor (_08486_, _08485_, _08309_);
  and (_08487_, _08471_, _08211_);
  nor (_08488_, _08475_, _08205_);
  and (_08489_, _08482_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08490_, _08489_, _08488_);
  and (_08491_, _08490_, _08328_);
  nor (_08492_, _08491_, _08487_);
  not (_08493_, _08492_);
  nor (_08494_, _08493_, _08486_);
  nor (_08495_, _08475_, _08230_);
  and (_08496_, _08480_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_08497_, _08482_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08498_, _08497_, _08496_);
  nor (_08499_, _08498_, _08495_);
  nor (_08500_, _08499_, _08337_);
  nor (_08501_, _08475_, _08219_);
  and (_08502_, _08480_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08503_, _08482_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08504_, _08503_, _08502_);
  nor (_08505_, _08504_, _08501_);
  nor (_08506_, _08505_, _08345_);
  nor (_08507_, _08506_, _08500_);
  and (_08508_, _08507_, _08494_);
  and (_08509_, _08368_, _08359_);
  and (_08510_, _08363_, _08358_);
  or (_08511_, _08510_, _08509_);
  and (_08512_, _08511_, _08482_);
  and (_08513_, _08380_, _08359_);
  and (_08514_, _08375_, _08358_);
  or (_08515_, _08514_, _08513_);
  and (_08516_, _08515_, _08480_);
  and (_08517_, _08474_, _08281_);
  and (_08518_, _08393_, _08359_);
  and (_08519_, _08388_, _08358_);
  or (_08520_, _08519_, _08518_);
  and (_08521_, _08520_, _08517_);
  and (_08522_, _08474_, _08184_);
  and (_08523_, _08405_, _08359_);
  and (_08524_, _08400_, _08358_);
  or (_08525_, _08524_, _08523_);
  and (_08526_, _08525_, _08522_);
  or (_08527_, _08526_, _08521_);
  or (_08528_, _08527_, _08516_);
  nor (_08529_, _08528_, _08512_);
  nor (_08530_, _08529_, _08508_);
  and (_08531_, _08508_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08531_, _08530_);
  and (_08532_, _08195_, _08184_);
  nor (_08533_, _08417_, _08203_);
  or (_08534_, _08533_, _08532_);
  and (_07359_, _08534_, _06071_);
  not (_08535_, _06526_);
  or (_08536_, _08535_, _05810_);
  or (_08537_, _06526_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_08538_, _08537_, _06071_);
  and (_07382_, _08538_, _08536_);
  and (_08539_, _08508_, _06071_);
  and (_08540_, _08539_, word_in[31]);
  and (_08541_, _08532_, _08328_);
  and (_08542_, _08539_, _08541_);
  and (_08543_, _08542_, _08540_);
  not (_08544_, _08542_);
  and (_08545_, _08450_, _06071_);
  and (_08546_, _08545_, _08414_);
  and (_08547_, _08546_, _08419_);
  and (_08548_, _08547_, _08308_);
  not (_08549_, _08548_);
  and (_08550_, _08357_, _06071_);
  and (_08551_, _08550_, _08344_);
  and (_08552_, _08551_, _08350_);
  and (_08553_, _08225_, _06071_);
  and (_08554_, _08553_, _08190_);
  nor (_08555_, _08253_, rst);
  and (_08556_, _08555_, _08532_);
  and (_08557_, _08556_, _08554_);
  and (_08558_, _08555_, word_in[7]);
  and (_08559_, _08558_, _08557_);
  nor (_08560_, _08557_, _08293_);
  nor (_08561_, _08560_, _08559_);
  nor (_08562_, _08561_, _08552_);
  and (_08563_, _08552_, word_in[15]);
  or (_08564_, _08563_, _08562_);
  and (_08565_, _08564_, _08549_);
  and (_08566_, _08545_, word_in[23]);
  and (_08567_, _08566_, _08548_);
  or (_08568_, _08567_, _08565_);
  and (_08569_, _08568_, _08544_);
  or (_14025_, _08569_, _08543_);
  or (_08570_, _08480_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07408_, _08570_, _06071_);
  or (_08571_, _08197_, _08184_);
  nor (_08572_, _08417_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_08573_, _08572_, _08571_);
  and (_07436_, _08573_, _06071_);
  and (_08574_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_08575_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_08576_, _08575_, _07912_);
  or (_08577_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_08578_, _08577_, _06560_);
  and (_08579_, _08578_, _08576_);
  or (_07472_, _08579_, _08574_);
  and (_08580_, _08311_, _08184_);
  not (_08581_, _08571_);
  nor (_08582_, _08581_, _08580_);
  not (_08583_, _08312_);
  or (_08584_, _08583_, _08184_);
  nor (_08585_, _08584_, _08207_);
  nor (_08586_, _08585_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_08587_, _08586_, _08582_);
  and (_07476_, _08587_, _06071_);
  and (_08588_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_08589_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_08590_, _08589_, _07912_);
  or (_08591_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_08592_, _08591_, _06560_);
  and (_08593_, _08592_, _08590_);
  or (_07482_, _08593_, _08588_);
  or (_08594_, _08535_, _05880_);
  or (_08595_, _06526_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_08596_, _08595_, _06071_);
  and (_07485_, _08596_, _08594_);
  and (_08597_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_08598_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_08599_, _08598_, _07912_);
  or (_08600_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_08601_, _08600_, _06560_);
  and (_08602_, _08601_, _08599_);
  or (_07510_, _08602_, _08597_);
  and (_08603_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_08604_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_08605_, _08604_, _07912_);
  or (_08606_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_08607_, _08606_, _06560_);
  and (_08608_, _08607_, _08605_);
  or (_07513_, _08608_, _08603_);
  or (_08609_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_08611_, _08609_, _07912_);
  or (_08612_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_08613_, _08612_, _06560_);
  and (_08614_, _08613_, _08611_);
  or (_07522_, _08614_, _06559_);
  not (_08615_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor (_08616_, _08016_, _08615_);
  nor (_08617_, _08616_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_08618_, _08616_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_08619_, _08618_, _08617_);
  nor (_07524_, _08619_, rst);
  not (_08620_, _08321_);
  and (_08621_, _08517_, _08310_);
  or (_08622_, _08195_, _08184_);
  or (_08623_, _08622_, _08344_);
  and (_08624_, _08623_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08625_, _08624_, _08621_);
  and (_08626_, _08625_, _08620_);
  and (_08627_, _08211_, _08196_);
  or (_08628_, _08627_, _08585_);
  or (_08629_, _08628_, _08626_);
  and (_08630_, _08629_, _08582_);
  or (_08631_, _08627_, _08625_);
  and (_08632_, _08631_, _08580_);
  or (_08633_, _08632_, _08581_);
  or (_08634_, _08633_, _08630_);
  and (_07529_, _08634_, _06071_);
  or (_08635_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_08636_, _08635_, _07912_);
  and (_08637_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_08638_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_08639_, _08638_, _06560_);
  or (_08640_, _08639_, _08637_);
  and (_07539_, _08640_, _08636_);
  or (_08641_, _08535_, _05788_);
  or (_08642_, _06526_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_08643_, _08642_, _06071_);
  and (_07568_, _08643_, _08641_);
  and (_08644_, _08328_, _08318_);
  or (_08645_, _08644_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08646_, _08645_, _08622_);
  or (_08647_, _08646_, _08621_);
  and (_08648_, _08647_, _08620_);
  and (_08649_, _08645_, _08580_);
  nand (_08650_, _08195_, _08174_);
  nand (_08651_, _08418_, _08650_);
  nor (_08652_, _08651_, _08309_);
  and (_08653_, _08471_, _08281_);
  and (_08654_, _08653_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08655_, _08654_, _08652_);
  or (_08656_, _08655_, _08649_);
  or (_08657_, _08656_, _08585_);
  or (_08658_, _08657_, _08648_);
  and (_07582_, _08658_, _06071_);
  and (_08659_, _08016_, _08615_);
  nor (_08660_, _08659_, _08616_);
  and (_07589_, _08660_, _06071_);
  or (_08661_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_08662_, _08661_, _07912_);
  and (_08663_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_08664_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and (_08665_, _08664_, _06560_);
  or (_08666_, _08665_, _08663_);
  and (_07620_, _08666_, _08662_);
  or (_08667_, _07887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_08668_, _08667_, _07912_);
  and (_08669_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_08670_, _07897_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and (_08671_, _08670_, _06560_);
  or (_08672_, _08671_, _08669_);
  and (_07629_, _08672_, _08668_);
  not (_08673_, _08417_);
  and (_08674_, _08584_, _08673_);
  and (_08675_, _08201_, _08184_);
  or (_08676_, _08675_, _08318_);
  not (_08677_, _08418_);
  or (_08678_, _08644_, _08621_);
  or (_08679_, _08678_, _08677_);
  and (_08680_, _08679_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08681_, _08585_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08682_, _08308_, _08318_);
  and (_08683_, _08581_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08684_, _08683_, _08682_);
  or (_08685_, _08684_, _08681_);
  or (_08686_, _08685_, _08680_);
  or (_08687_, _08316_, _08477_);
  and (_08688_, _08687_, _08686_);
  and (_08689_, _08517_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08690_, _08689_, _08644_);
  or (_08691_, _08690_, _08688_);
  and (_08692_, _08691_, _08676_);
  and (_08693_, _08686_, _08580_);
  or (_08694_, _08683_, _08621_);
  or (_08695_, _08694_, _08681_);
  or (_08696_, _08695_, _08693_);
  or (_08697_, _08696_, _08692_);
  and (_08698_, _08697_, _08674_);
  and (_08699_, _08532_, _08344_);
  and (_08700_, _08691_, _08699_);
  or (_08701_, _08683_, _08585_);
  or (_08702_, _08701_, _08693_);
  or (_08703_, _08702_, _08700_);
  or (_08704_, _08703_, _08698_);
  and (_07640_, _08704_, _06071_);
  and (_08705_, _06527_, _05689_);
  not (_08706_, _08705_);
  or (_08707_, _08706_, _05829_);
  not (_08708_, _05689_);
  nor (_08709_, _06527_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_08710_, _08709_, _08708_);
  nand (_08711_, _08710_, _08707_);
  or (_08712_, _08706_, _05847_);
  nor (_08713_, _06527_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_08714_, _08713_, _08708_);
  nand (_08715_, _08714_, _08712_);
  and (_08717_, _08715_, _08711_);
  or (_08718_, _08706_, _05788_);
  nor (_08719_, _06527_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_08720_, _08719_, _08708_);
  nand (_08721_, _08720_, _08718_);
  or (_08722_, _08706_, _05810_);
  nor (_08723_, _06527_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_08724_, _08723_, _08708_);
  and (_08725_, _08724_, _08722_);
  not (_08726_, _08725_);
  and (_08727_, _08726_, _08721_);
  and (_08728_, _08727_, _08717_);
  or (_08729_, _08706_, _05880_);
  nor (_08730_, _06527_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_08731_, _08730_, _08708_);
  and (_08732_, _08731_, _08729_);
  or (_08733_, _08706_, _05768_);
  nor (_08734_, _06527_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_08735_, _08734_, _08708_);
  and (_08736_, _08735_, _08733_);
  or (_08737_, _08706_, _05747_);
  nor (_08739_, _06527_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_08740_, _08739_, _08708_);
  nand (_08741_, _08740_, _08737_);
  or (_08742_, _08706_, _05726_);
  nor (_08744_, _06527_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_08745_, _08744_, _08708_);
  nand (_08746_, _08745_, _08742_);
  nor (_08748_, _08746_, _08741_);
  and (_08749_, _08748_, _08736_);
  and (_08750_, _08749_, _08732_);
  nand (_08752_, _08750_, _08728_);
  and (_08753_, _08720_, _08718_);
  and (_08754_, _08725_, _08711_);
  and (_08756_, _08754_, _08715_);
  and (_08757_, _08756_, _08753_);
  and (_08758_, _08746_, _08741_);
  and (_08760_, _08758_, _08736_);
  and (_08761_, _08760_, _08757_);
  not (_08762_, _08761_);
  not (_08764_, _08732_);
  and (_08765_, _08749_, _08764_);
  and (_08767_, _08765_, _08728_);
  and (_08768_, _08765_, _08756_);
  nor (_08769_, _08768_, _08767_);
  and (_08770_, _08769_, _08762_);
  and (_08771_, _08770_, _08752_);
  and (_08772_, _08732_, _08715_);
  and (_08773_, _08772_, _08749_);
  and (_08774_, _08773_, _08754_);
  and (_08775_, _06527_, _06071_);
  not (_08776_, _08775_);
  or (_08777_, _08776_, _08768_);
  or (_08778_, _08777_, _08774_);
  or (_07649_, _08778_, _08771_);
  or (_08779_, _08428_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08780_, _08779_, _08651_);
  and (_08781_, _08780_, _08677_);
  and (_08782_, _08678_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08783_, _08782_, _08682_);
  or (_08784_, _08783_, _08781_);
  and (_08785_, _08784_, _08687_);
  and (_08786_, _08779_, _08580_);
  and (_08787_, _08585_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08788_, _08581_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08789_, _08788_, _08621_);
  or (_08790_, _08789_, _08787_);
  or (_08791_, _08790_, _08644_);
  or (_08792_, _08791_, _08786_);
  or (_08793_, _08792_, _08785_);
  and (_07708_, _08793_, _06071_);
  nand (_08794_, _07823_, _07520_);
  or (_08795_, _07772_, _07425_);
  nor (_08796_, _07826_, _06271_);
  nor (_08797_, _08796_, _07773_);
  not (_08798_, _08797_);
  not (_08799_, _06803_);
  and (_08800_, _06004_, _07752_);
  and (_08801_, _08800_, _05982_);
  and (_08802_, _08801_, _08799_);
  nor (_08803_, _08801_, _06271_);
  nor (_08804_, _08803_, _08802_);
  and (_08805_, _07831_, _07826_);
  not (_08806_, _08805_);
  nor (_08807_, _08806_, _08804_);
  nor (_08808_, _08807_, _08798_);
  nor (_08809_, _08808_, _07823_);
  nand (_08810_, _08809_, _08795_);
  nand (_08811_, _08810_, _08794_);
  and (_07736_, _08811_, _06071_);
  not (_08812_, _08320_);
  and (_08813_, _08653_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08814_, _08517_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_08815_, _08814_, _08329_);
  or (_08816_, _08815_, _08813_);
  or (_08817_, _08428_, _08184_);
  and (_08818_, _08817_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_08819_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_08820_, _08190_, _08819_);
  and (_08821_, _08820_, _08318_);
  or (_08822_, _08821_, _08319_);
  or (_08823_, _08822_, _08818_);
  or (_08824_, _08823_, _08816_);
  and (_08825_, _08824_, _08812_);
  or (_08826_, _08821_, _08428_);
  or (_08827_, _08826_, _08815_);
  or (_08828_, _08827_, _08825_);
  and (_08829_, _08828_, _08677_);
  and (_08830_, _08824_, _08580_);
  or (_08831_, _08813_, _08644_);
  or (_08832_, _08831_, _08814_);
  or (_08833_, _08832_, _08682_);
  or (_08834_, _08833_, _08830_);
  or (_08835_, _08834_, _08829_);
  and (_07780_, _08835_, _06071_);
  nor (_08836_, _08482_, _08281_);
  and (_08837_, _08836_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08838_, _08471_, _08184_);
  nor (_08839_, _08195_, _08246_);
  or (_08840_, _08839_, _08311_);
  and (_08841_, _08840_, _08281_);
  and (_08842_, _08644_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08843_, _08842_, _08682_);
  or (_08844_, _08843_, _08841_);
  or (_08845_, _08844_, _08428_);
  or (_08847_, _08845_, _08838_);
  or (_08848_, _08847_, _08837_);
  and (_07842_, _08848_, _06071_);
  and (_08849_, _08478_, _08308_);
  nor (_08851_, _08675_, _08311_);
  nor (_08852_, _08851_, _08849_);
  or (_08854_, _08682_, _08653_);
  or (_08856_, _08854_, _08852_);
  or (_08857_, _08856_, _08699_);
  or (_08859_, _08857_, _08517_);
  and (_08861_, _08859_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08862_, _08861_, _08420_);
  and (_07921_, _08862_, _06071_);
  and (_08864_, _06381_, _06011_);
  not (_08865_, _08864_);
  and (_08867_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_08869_, _08865_, _07945_);
  or (_08871_, _08869_, _08867_);
  and (_07982_, _08871_, _06071_);
  or (_08873_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_08874_, _06530_, _05815_);
  and (_08876_, _08874_, _06071_);
  and (_07987_, _08876_, _08873_);
  and (_08877_, _08532_, _08308_);
  or (_08878_, _08877_, _08522_);
  or (_08879_, _08878_, _08699_);
  and (_08880_, _08316_, _08197_);
  and (_08881_, _08428_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08882_, _08678_, _08682_);
  and (_08883_, _08882_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08884_, _08883_, _08881_);
  and (_08885_, _08849_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_08886_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08887_, _08358_, _08886_);
  and (_08888_, _08887_, _08517_);
  and (_08889_, _08653_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08891_, _08522_, _08344_);
  and (_08892_, _08583_, _08239_);
  or (_08893_, _08892_, _08891_);
  or (_08895_, _08893_, _08889_);
  or (_08896_, _08895_, _08888_);
  or (_08897_, _08896_, _08885_);
  or (_08898_, _08897_, _08884_);
  and (_08899_, _08898_, _08880_);
  or (_08900_, _08319_, _08838_);
  and (_08901_, _08900_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08902_, _08901_, _08849_);
  or (_08903_, _08902_, _08899_);
  and (_08904_, _08903_, _08879_);
  or (_08905_, _08901_, _08898_);
  and (_08906_, _08905_, _08580_);
  and (_08907_, _08414_, _08281_);
  and (_08908_, _08907_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08909_, _08571_, _08886_);
  or (_08910_, _08909_, _08319_);
  or (_08911_, _08910_, _08881_);
  or (_08912_, _08911_, _08908_);
  or (_08913_, _08912_, _08838_);
  or (_08914_, _08913_, _08906_);
  or (_08915_, _08914_, _08904_);
  and (_07995_, _08915_, _06071_);
  and (_08916_, _08532_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08917_, _08208_, _08184_);
  or (_08918_, _08174_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08919_, _08918_, _08917_);
  and (_08920_, _08208_, _08281_);
  and (_08921_, _08920_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08922_, _08921_, _08919_);
  or (_08923_, _08922_, _08916_);
  and (_08924_, _08212_, _08196_);
  not (_08925_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08926_, _08184_, _08925_);
  and (_08927_, _08926_, _08209_);
  or (_08928_, _08927_, _08924_);
  or (_08929_, _08928_, _08923_);
  and (_08930_, _08929_, _08350_);
  or (_08931_, _08924_, _08891_);
  or (_08932_, _08931_, _08930_);
  and (_08933_, _08932_, _08197_);
  and (_08934_, _08929_, _08580_);
  or (_08935_, _08934_, _08838_);
  or (_08936_, _08935_, _08849_);
  or (_08937_, _08936_, _08926_);
  or (_08938_, _08937_, _08933_);
  and (_08055_, _08938_, _06071_);
  or (_08939_, _07772_, _07643_);
  not (_08940_, _07826_);
  and (_08941_, _07831_, _08940_);
  and (_08942_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_08943_, _08799_, _06032_);
  nor (_08944_, _06032_, _06292_);
  nor (_08945_, _08944_, _08943_);
  nor (_08946_, _08945_, _08806_);
  nor (_08947_, _08946_, _08942_);
  and (_08948_, _08947_, _07830_);
  nand (_08949_, _08948_, _08939_);
  and (_08950_, _07823_, _07673_);
  not (_08951_, _08950_);
  and (_08952_, _08951_, _08949_);
  and (_08085_, _08952_, _06071_);
  or (_08953_, _08053_, _07772_);
  and (_08954_, _07826_, _06383_);
  and (_08955_, _08954_, _06803_);
  nor (_08956_, _08954_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_08957_, _08956_, _07832_);
  not (_08958_, _08957_);
  nor (_08959_, _08958_, _08955_);
  nor (_08961_, _08959_, _07823_);
  nand (_08962_, _08961_, _08953_);
  or (_08963_, _08139_, _07830_);
  and (_08964_, _08963_, _08962_);
  and (_08089_, _08964_, _06071_);
  and (_08966_, _08532_, _08329_);
  and (_08967_, _08966_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08968_, _08190_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08970_, _08968_, _08517_);
  and (_08971_, _08838_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_08973_, _08571_, _08233_);
  and (_08974_, _08318_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_08975_, _08974_, _08973_);
  or (_08977_, _08975_, _08971_);
  or (_08978_, _08977_, _08522_);
  or (_08979_, _08978_, _08970_);
  or (_08980_, _08979_, _08967_);
  and (_08149_, _08980_, _06071_);
  and (_08982_, _07104_, _06383_);
  and (_08984_, _08982_, _05968_);
  nand (_08985_, _08984_, _06365_);
  and (_08986_, _08985_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_08987_, _06365_, _05968_);
  and (_08988_, _08987_, _08982_);
  not (_08989_, _08988_);
  nor (_08990_, _08989_, _06993_);
  nor (_08991_, _08990_, _08986_);
  nor (_08157_, _08991_, rst);
  not (_08992_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_08993_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_08994_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08993_);
  not (_08995_, _08994_);
  and (_08996_, _07902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_08997_, _08996_, _08995_);
  and (_08998_, _08997_, _07900_);
  nor (_08999_, _08998_, _08992_);
  and (_09000_, _08998_, rxd_i);
  or (_09001_, _09000_, rst);
  or (_08216_, _09001_, _08999_);
  not (_09002_, rxd_i);
  nor (_09003_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_09004_, _09003_, _07892_);
  and (_09005_, _07890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09006_, _09005_, _09004_);
  nand (_09007_, _09006_, _09002_);
  or (_09008_, _09006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_09009_, _09008_, _06071_);
  and (_08226_, _09009_, _09007_);
  and (_09010_, _08190_, _08184_);
  or (_09011_, _08346_, _09010_);
  and (_09012_, _09011_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_09013_, _09012_, _08207_);
  and (_09014_, _09013_, _08966_);
  or (_09015_, _08541_, _08917_);
  nor (_09016_, _09010_, _08532_);
  and (_09017_, _09016_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_09018_, _09017_, _09015_);
  or (_09019_, _09018_, _09014_);
  and (_08265_, _09019_, _06071_);
  or (_09020_, _08350_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08385_, _09020_, _06071_);
  or (_09021_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not (_09022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_09023_, _06530_, _09022_);
  and (_09024_, _09023_, _06071_);
  and (_08447_, _09024_, _09021_);
  not (_09025_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nor (_09026_, _05954_, _07767_);
  and (_09027_, _09026_, _06809_);
  and (_09028_, _09027_, _06815_);
  nand (_09029_, _09028_, _06362_);
  nand (_09030_, _09029_, _09025_);
  and (_09031_, _09030_, _08989_);
  or (_09032_, _09029_, _08799_);
  and (_09033_, _09032_, _09031_);
  nor (_09034_, _06355_, _06856_);
  not (_09035_, _09034_);
  and (_09036_, _09035_, _08094_);
  and (_09037_, _09036_, _08079_);
  nor (_09038_, _09037_, _08989_);
  or (_09039_, _09038_, _09033_);
  and (_08610_, _09039_, _06071_);
  nand (_09040_, _07946_, _06434_);
  or (_09041_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_09042_, _09041_, _06071_);
  and (_08716_, _09042_, _09040_);
  and (_09043_, _08539_, word_in[24]);
  and (_09044_, _08539_, _08877_);
  and (_09045_, _09044_, _09043_);
  and (_09046_, _08545_, _08699_);
  not (_09047_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_09048_, _08555_, _08190_);
  nor (_09049_, _09048_, _08553_);
  and (_09050_, _08555_, _08622_);
  not (_09051_, _09050_);
  and (_09052_, _09051_, _09049_);
  and (_09053_, _09052_, _08555_);
  nor (_09054_, _09053_, _09047_);
  and (_09056_, _08555_, word_in[0]);
  and (_09057_, _09056_, _09052_);
  or (_09059_, _09057_, _09054_);
  and (_09061_, _08550_, _08580_);
  not (_09062_, _09061_);
  and (_09063_, _09062_, _09059_);
  and (_09064_, _09061_, word_in[8]);
  or (_09066_, _09064_, _09063_);
  or (_09067_, _09066_, _09046_);
  not (_09068_, _09044_);
  not (_09070_, _09046_);
  or (_09071_, _09070_, word_in[16]);
  and (_09072_, _09071_, _09068_);
  and (_09073_, _09072_, _09067_);
  or (_08738_, _09073_, _09045_);
  and (_09075_, _08539_, word_in[25]);
  and (_09076_, _09075_, _09044_);
  not (_09078_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_09079_, _09053_, _09078_);
  and (_09080_, _08555_, word_in[1]);
  and (_09081_, _09080_, _09052_);
  or (_09082_, _09081_, _09079_);
  or (_09083_, _09082_, _09061_);
  or (_09084_, _09062_, word_in[9]);
  and (_09085_, _09084_, _09070_);
  and (_09086_, _09085_, _09083_);
  and (_09088_, _09046_, word_in[17]);
  or (_09089_, _09088_, _09086_);
  and (_09090_, _09089_, _09068_);
  or (_08743_, _09090_, _09076_);
  or (_09091_, _09062_, word_in[10]);
  and (_09092_, _09091_, _09070_);
  not (_09093_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_09094_, _09053_, _09093_);
  and (_09095_, _09053_, word_in[2]);
  or (_09096_, _09095_, _09094_);
  or (_09097_, _09096_, _09061_);
  and (_09098_, _09097_, _09092_);
  and (_09099_, _09046_, word_in[18]);
  or (_09100_, _09099_, _09044_);
  or (_09101_, _09100_, _09098_);
  or (_09102_, _09068_, word_in[26]);
  and (_08747_, _09102_, _09101_);
  and (_09103_, _08539_, word_in[27]);
  and (_09104_, _09103_, _09044_);
  not (_09105_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_09106_, _09053_, _09105_);
  and (_09107_, _09053_, word_in[3]);
  or (_09108_, _09107_, _09106_);
  and (_09109_, _09108_, _09062_);
  and (_09110_, _09061_, word_in[11]);
  or (_09111_, _09110_, _09109_);
  and (_09112_, _09111_, _09070_);
  and (_09113_, _08545_, word_in[19]);
  and (_09114_, _09113_, _08699_);
  or (_09115_, _09114_, _09112_);
  and (_09116_, _09115_, _09068_);
  or (_08751_, _09116_, _09104_);
  or (_09117_, _09062_, word_in[12]);
  and (_09118_, _09117_, _09070_);
  and (_09119_, _09053_, word_in[4]);
  not (_09120_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_09121_, _09053_, _09120_);
  or (_09122_, _09121_, _09119_);
  or (_09123_, _09122_, _09061_);
  and (_09124_, _09123_, _09118_);
  and (_09125_, _09046_, word_in[20]);
  or (_09126_, _09125_, _09044_);
  or (_09127_, _09126_, _09124_);
  or (_09128_, _09068_, word_in[28]);
  and (_08755_, _09128_, _09127_);
  or (_09129_, _09062_, word_in[13]);
  and (_09130_, _09129_, _09070_);
  not (_09131_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_09132_, _09053_, _09131_);
  and (_09133_, _09053_, word_in[5]);
  or (_09134_, _09133_, _09132_);
  or (_09135_, _09134_, _09061_);
  and (_09136_, _09135_, _09130_);
  and (_09137_, _09046_, word_in[21]);
  or (_09138_, _09137_, _09136_);
  and (_09139_, _09138_, _09068_);
  and (_09140_, _08539_, word_in[29]);
  and (_09141_, _09140_, _09044_);
  or (_08759_, _09141_, _09139_);
  or (_09142_, _09062_, word_in[14]);
  and (_09143_, _09142_, _09070_);
  not (_09144_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_09145_, _09053_, _09144_);
  and (_09146_, _09053_, word_in[6]);
  or (_09147_, _09146_, _09145_);
  or (_09149_, _09147_, _09061_);
  and (_09150_, _09149_, _09143_);
  and (_09151_, _09046_, word_in[22]);
  or (_09152_, _09151_, _09044_);
  or (_09153_, _09152_, _09150_);
  or (_09154_, _09068_, word_in[30]);
  and (_08763_, _09154_, _09153_);
  or (_09155_, _09068_, word_in[31]);
  nor (_09156_, _09053_, _08377_);
  and (_09157_, _09053_, _08558_);
  or (_09158_, _09157_, _09156_);
  or (_09159_, _09158_, _09061_);
  or (_09160_, _09062_, word_in[15]);
  and (_09162_, _09160_, _09070_);
  and (_09163_, _09162_, _09159_);
  and (_09165_, _08566_, _08699_);
  or (_09166_, _09165_, _09044_);
  or (_09167_, _09166_, _09163_);
  and (_08766_, _09167_, _09155_);
  and (_09168_, _08545_, word_in[16]);
  and (_09169_, _08545_, _08310_);
  and (_09170_, _09169_, _08422_);
  and (_09171_, _09170_, _09168_);
  not (_09172_, _09170_);
  and (_09173_, _08550_, _08328_);
  and (_09174_, _09173_, _08321_);
  not (_09175_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_09177_, _08553_, _08207_);
  and (_09178_, _09177_, _09051_);
  nor (_09180_, _09178_, _09175_);
  and (_09181_, _09178_, _09056_);
  nor (_09182_, _09181_, _09180_);
  nor (_09183_, _09182_, _09174_);
  and (_09184_, _09174_, word_in[8]);
  or (_09185_, _09184_, _09183_);
  and (_09187_, _09185_, _09172_);
  or (_09188_, _09187_, _09171_);
  and (_09189_, _08539_, _08699_);
  not (_09190_, _09189_);
  and (_09191_, _09190_, _09188_);
  and (_09192_, _09189_, word_in[24]);
  or (_08846_, _09192_, _09191_);
  and (_09194_, _08545_, word_in[17]);
  and (_09195_, _09170_, _09194_);
  and (_09196_, _09178_, _09080_);
  not (_09197_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09198_, _09178_, _09197_);
  nor (_09199_, _09198_, _09196_);
  nor (_09200_, _09199_, _09174_);
  and (_09201_, _09174_, word_in[9]);
  or (_09202_, _09201_, _09200_);
  and (_09203_, _09202_, _09172_);
  or (_09204_, _09203_, _09195_);
  and (_09205_, _09204_, _09190_);
  and (_09206_, _09189_, word_in[25]);
  or (_08850_, _09206_, _09205_);
  nor (_09207_, t2_i, rst);
  and (_08853_, _09207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not (_09208_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09209_, _09178_, _09208_);
  and (_09210_, _08555_, word_in[2]);
  and (_09211_, _09178_, _09210_);
  nor (_09212_, _09211_, _09209_);
  nor (_09213_, _09212_, _09174_);
  and (_09214_, _09174_, word_in[10]);
  or (_09215_, _09214_, _09213_);
  and (_09216_, _09215_, _09172_);
  and (_09217_, _08545_, word_in[18]);
  and (_09218_, _09170_, _09217_);
  or (_09219_, _09218_, _09216_);
  and (_09220_, _09219_, _09190_);
  and (_09221_, _09189_, word_in[26]);
  or (_08855_, _09221_, _09220_);
  not (_09222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_09223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _09222_);
  not (_09224_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_09225_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_09226_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _06445_);
  nor (_09227_, _09226_, _09225_);
  nor (_09228_, _09227_, _06444_);
  nor (_09229_, _09228_, _09224_);
  and (_09230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_09231_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _06445_);
  nor (_09232_, _09231_, _09230_);
  nor (_09233_, _09232_, _06444_);
  not (_09234_, _09233_);
  and (_09236_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_09237_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _06445_);
  nor (_09238_, _09237_, _09236_);
  nor (_09239_, _09238_, _06444_);
  and (_09240_, _09239_, _09234_);
  nand (_09241_, _09240_, _09229_);
  and (_09242_, _09241_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_09243_, _09242_, _09223_);
  and (_09244_, _06032_, _06378_);
  and (_09245_, _06840_, _09244_);
  and (_09246_, _09245_, _06815_);
  or (_09247_, _09246_, _09243_);
  and (_09248_, _06383_, _06027_);
  and (_09249_, _09248_, _06840_);
  not (_09250_, _09249_);
  and (_09251_, _09250_, _09247_);
  nand (_09252_, _09246_, _06803_);
  and (_09254_, _09252_, _09251_);
  nor (_09255_, _09250_, _06609_);
  or (_09256_, _09255_, _09254_);
  and (_08858_, _09256_, _06071_);
  not (_09258_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09259_, _09178_, _09258_);
  and (_09260_, _08555_, word_in[3]);
  and (_09262_, _09178_, _09260_);
  nor (_09263_, _09262_, _09259_);
  nor (_09264_, _09263_, _09174_);
  and (_09265_, _09174_, word_in[11]);
  or (_09267_, _09265_, _09264_);
  and (_09268_, _09267_, _09172_);
  and (_09269_, _09170_, _09113_);
  or (_09271_, _09269_, _09268_);
  and (_09272_, _09271_, _09190_);
  and (_09273_, _09189_, word_in[27]);
  or (_08860_, _09273_, _09272_);
  not (_09275_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09276_, _09178_, _09275_);
  and (_09277_, _08555_, word_in[4]);
  and (_09279_, _09178_, _09277_);
  or (_09280_, _09279_, _09276_);
  or (_09282_, _09280_, _09174_);
  not (_09283_, _09174_);
  or (_09284_, _09283_, word_in[12]);
  and (_09285_, _09284_, _09282_);
  and (_09286_, _09285_, _09172_);
  and (_09287_, _08545_, word_in[20]);
  and (_09288_, _09170_, _09287_);
  or (_09289_, _09288_, _09286_);
  or (_09290_, _09289_, _09189_);
  or (_09291_, _09190_, word_in[28]);
  and (_08863_, _09291_, _09290_);
  and (_09292_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_09293_, _06967_, _06609_);
  or (_09294_, _09293_, _09292_);
  and (_08866_, _09294_, _06071_);
  not (_09295_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09296_, _09178_, _09295_);
  and (_09297_, _08555_, word_in[5]);
  and (_09298_, _09178_, _09297_);
  or (_09299_, _09298_, _09296_);
  or (_09301_, _09299_, _09174_);
  or (_09302_, _09283_, word_in[13]);
  and (_09303_, _09302_, _09301_);
  or (_09304_, _09303_, _09170_);
  and (_09305_, _08545_, word_in[21]);
  or (_09306_, _09172_, _09305_);
  and (_09307_, _09306_, _09304_);
  or (_09308_, _09307_, _09189_);
  or (_09309_, _09190_, word_in[29]);
  and (_08868_, _09309_, _09308_);
  nor (_09310_, _06434_, _06400_);
  and (_09311_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_09312_, _09311_, _09310_);
  and (_08870_, _09312_, _06071_);
  not (_09313_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09314_, _09178_, _09313_);
  and (_09315_, _08555_, word_in[6]);
  and (_09316_, _09178_, _09315_);
  nor (_09317_, _09316_, _09314_);
  nor (_09318_, _09317_, _09174_);
  and (_09319_, _09174_, word_in[14]);
  or (_09320_, _09319_, _09318_);
  and (_09321_, _09320_, _09172_);
  and (_09322_, _08545_, word_in[22]);
  and (_09323_, _09170_, _09322_);
  or (_09324_, _09323_, _09321_);
  and (_09325_, _09324_, _09190_);
  and (_09326_, _09189_, word_in[30]);
  or (_08872_, _09326_, _09325_);
  and (_09327_, _09170_, _08566_);
  and (_09328_, _09178_, _08558_);
  nor (_09329_, _09178_, _08256_);
  nor (_09330_, _09329_, _09328_);
  nor (_09331_, _09330_, _09174_);
  and (_09332_, _09174_, word_in[15]);
  or (_09333_, _09332_, _09331_);
  and (_09334_, _09333_, _09172_);
  or (_09335_, _09334_, _09327_);
  and (_09336_, _09335_, _09190_);
  and (_09337_, _09189_, word_in[31]);
  or (_08875_, _09337_, _09336_);
  nor (_09338_, _06355_, _06276_);
  not (_09339_, _09338_);
  and (_09340_, _09339_, _07410_);
  and (_09341_, _09340_, _07388_);
  nor (_09342_, _09341_, _06967_);
  and (_09343_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_09344_, _09343_, _09342_);
  and (_08890_, _09344_, _06071_);
  or (_09345_, _06965_, _06391_);
  nor (_09346_, _09345_, _06392_);
  or (_09347_, _09346_, _06390_);
  and (_09348_, _09347_, _06400_);
  or (_09349_, _09348_, _06392_);
  and (_09350_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_09351_, _07945_, _06400_);
  and (_09352_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_09353_, _09352_, _09345_);
  or (_09354_, _09353_, _09351_);
  or (_09355_, _09354_, _09350_);
  and (_08894_, _09355_, _06071_);
  and (_09357_, _08545_, _08328_);
  and (_09358_, _09357_, _08422_);
  not (_09359_, _09358_);
  and (_09361_, _08550_, _08308_);
  and (_09362_, _09361_, _08321_);
  not (_09364_, _08553_);
  and (_09365_, _09048_, _09364_);
  and (_09367_, _09365_, _09051_);
  and (_09368_, _09367_, _09056_);
  not (_09369_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_09370_, _09367_, _09369_);
  nor (_09372_, _09370_, _09368_);
  nor (_09374_, _09372_, _09362_);
  and (_09375_, _09362_, word_in[8]);
  or (_09377_, _09375_, _09374_);
  and (_09378_, _09377_, _09359_);
  and (_09380_, _08539_, _08580_);
  and (_09381_, _09358_, _09168_);
  or (_09382_, _09381_, _09380_);
  or (_09383_, _09382_, _09378_);
  not (_09384_, _09380_);
  or (_09385_, _09384_, word_in[24]);
  and (_08960_, _09385_, _09383_);
  not (_09386_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09387_, _09367_, _09386_);
  and (_09388_, _09367_, _09080_);
  or (_09389_, _09388_, _09387_);
  or (_09390_, _09389_, _09362_);
  not (_09391_, _09362_);
  or (_09392_, _09391_, word_in[9]);
  and (_09393_, _09392_, _09390_);
  or (_09394_, _09393_, _09358_);
  or (_09395_, _09359_, _09194_);
  and (_09396_, _09395_, _09384_);
  and (_09397_, _09396_, _09394_);
  and (_09398_, _09380_, word_in[25]);
  or (_08965_, _09398_, _09397_);
  and (_09399_, _09367_, _09210_);
  not (_09400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09401_, _09367_, _09400_);
  nor (_09402_, _09401_, _09399_);
  nor (_09403_, _09402_, _09362_);
  and (_09404_, _09362_, word_in[10]);
  or (_09405_, _09404_, _09403_);
  and (_09406_, _09405_, _09359_);
  and (_09407_, _09358_, _09217_);
  or (_09408_, _09407_, _09380_);
  or (_09409_, _09408_, _09406_);
  or (_09410_, _09384_, word_in[26]);
  and (_08969_, _09410_, _09409_);
  and (_09411_, _09358_, _09113_);
  and (_09412_, _09367_, _09260_);
  not (_09413_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09414_, _09367_, _09413_);
  nor (_09415_, _09414_, _09412_);
  nor (_09416_, _09415_, _09362_);
  and (_09417_, _09362_, word_in[11]);
  or (_09418_, _09417_, _09416_);
  and (_09419_, _09418_, _09359_);
  or (_09420_, _09419_, _09411_);
  and (_09421_, _09420_, _09384_);
  and (_09422_, _09380_, word_in[27]);
  or (_08972_, _09422_, _09421_);
  and (_09423_, _09367_, _09277_);
  not (_09424_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09425_, _09367_, _09424_);
  nor (_09426_, _09425_, _09423_);
  nor (_09427_, _09426_, _09362_);
  and (_09428_, _09362_, word_in[12]);
  or (_09429_, _09428_, _09427_);
  and (_09430_, _09429_, _09359_);
  and (_09431_, _09358_, _09287_);
  or (_09432_, _09431_, _09380_);
  or (_09433_, _09432_, _09430_);
  or (_09434_, _09384_, word_in[28]);
  and (_08976_, _09434_, _09433_);
  not (_09435_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_09436_, _09367_, _09435_);
  and (_09437_, _09367_, _09297_);
  or (_09438_, _09437_, _09436_);
  or (_09439_, _09438_, _09362_);
  or (_09440_, _09391_, word_in[13]);
  and (_09441_, _09440_, _09439_);
  or (_09442_, _09441_, _09358_);
  or (_09443_, _09359_, _09305_);
  and (_09444_, _09443_, _09384_);
  and (_09445_, _09444_, _09442_);
  and (_09446_, _09380_, word_in[29]);
  or (_14026_, _09446_, _09445_);
  and (_09447_, _09367_, _09315_);
  not (_09448_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09449_, _09367_, _09448_);
  nor (_09450_, _09449_, _09447_);
  nor (_09451_, _09450_, _09362_);
  and (_09452_, _09362_, word_in[14]);
  or (_09453_, _09452_, _09451_);
  and (_09454_, _09453_, _09359_);
  and (_09455_, _09358_, _09322_);
  or (_09456_, _09455_, _09380_);
  or (_09457_, _09456_, _09454_);
  or (_09458_, _09384_, word_in[30]);
  and (_08981_, _09458_, _09457_);
  and (_09459_, _09358_, _08566_);
  and (_09460_, _09367_, _08558_);
  nor (_09461_, _09367_, _08372_);
  nor (_09462_, _09461_, _09460_);
  nor (_09463_, _09462_, _09362_);
  and (_09464_, _09362_, word_in[15]);
  or (_09465_, _09464_, _09463_);
  and (_09466_, _09465_, _09359_);
  or (_09467_, _09466_, _09459_);
  and (_09468_, _09467_, _09384_);
  and (_09469_, _09380_, word_in[31]);
  or (_08983_, _09469_, _09468_);
  and (_09470_, _08539_, _08653_);
  not (_09471_, _09470_);
  and (_09472_, _08545_, _08308_);
  and (_09473_, _09472_, _08422_);
  not (_09474_, _09473_);
  and (_09475_, _08551_, _08321_);
  not (_09476_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_09477_, _09051_, _08554_);
  nor (_09478_, _09477_, _09476_);
  and (_09479_, _09477_, _09056_);
  nor (_09480_, _09479_, _09478_);
  nor (_09481_, _09480_, _09475_);
  and (_09482_, _09475_, word_in[8]);
  or (_09483_, _09482_, _09481_);
  and (_09484_, _09483_, _09474_);
  and (_09485_, _09473_, _09168_);
  or (_09486_, _09485_, _09484_);
  and (_09487_, _09486_, _09471_);
  and (_09488_, _09470_, word_in[24]);
  or (_14027_, _09488_, _09487_);
  and (_09489_, _09477_, _09080_);
  not (_09490_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09491_, _09477_, _09490_);
  nor (_09492_, _09491_, _09489_);
  nor (_09493_, _09492_, _09475_);
  and (_09494_, _09475_, word_in[9]);
  or (_09495_, _09494_, _09493_);
  and (_09496_, _09495_, _09474_);
  and (_09497_, _09473_, _09194_);
  or (_09498_, _09497_, _09496_);
  and (_09499_, _09498_, _09471_);
  and (_09500_, _09470_, word_in[25]);
  or (_09055_, _09500_, _09499_);
  and (_09501_, _09477_, _09210_);
  not (_09502_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09503_, _09477_, _09502_);
  nor (_09504_, _09503_, _09501_);
  nor (_09505_, _09504_, _09475_);
  and (_09506_, _09475_, word_in[10]);
  or (_09507_, _09506_, _09505_);
  and (_09508_, _09507_, _09474_);
  and (_09509_, _09473_, _09217_);
  or (_09510_, _09509_, _09508_);
  and (_09511_, _09510_, _09471_);
  and (_09512_, _09470_, word_in[26]);
  or (_09058_, _09512_, _09511_);
  not (_09513_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09514_, _09477_, _09513_);
  and (_09515_, _09477_, _09260_);
  nor (_09516_, _09515_, _09514_);
  nor (_09517_, _09516_, _09475_);
  and (_09518_, _09475_, word_in[11]);
  or (_09519_, _09518_, _09517_);
  and (_09520_, _09519_, _09474_);
  and (_09521_, _09473_, _09113_);
  or (_09522_, _09521_, _09520_);
  and (_09523_, _09522_, _09471_);
  and (_09524_, _09470_, word_in[27]);
  or (_09060_, _09524_, _09523_);
  not (_09525_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_09526_, _09477_, _09525_);
  and (_09527_, _09477_, _09277_);
  nor (_09528_, _09527_, _09526_);
  nor (_09529_, _09528_, _09475_);
  and (_09530_, _09475_, word_in[12]);
  or (_09531_, _09530_, _09529_);
  and (_09532_, _09531_, _09474_);
  and (_09533_, _09473_, _09287_);
  or (_09534_, _09533_, _09532_);
  and (_09535_, _09534_, _09471_);
  and (_09536_, _09470_, word_in[28]);
  or (_09065_, _09536_, _09535_);
  and (_09537_, _09477_, _09297_);
  not (_09538_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_09539_, _09477_, _09538_);
  nor (_09540_, _09539_, _09537_);
  nor (_09541_, _09540_, _09475_);
  and (_09542_, _09475_, word_in[13]);
  or (_09543_, _09542_, _09541_);
  and (_09544_, _09543_, _09474_);
  and (_09545_, _09473_, _09305_);
  or (_09546_, _09545_, _09544_);
  and (_09548_, _09546_, _09471_);
  and (_09549_, _09470_, word_in[29]);
  or (_09069_, _09549_, _09548_);
  not (_09550_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_09552_, _09477_, _09550_);
  and (_09553_, _09477_, _09315_);
  or (_09554_, _09553_, _09552_);
  or (_09555_, _09554_, _09475_);
  not (_09556_, word_in[14]);
  nand (_09557_, _09475_, _09556_);
  and (_09558_, _09557_, _09555_);
  or (_09559_, _09558_, _09473_);
  or (_09560_, _09474_, _09322_);
  and (_09561_, _09560_, _09471_);
  and (_09562_, _09561_, _09559_);
  and (_09563_, _09470_, word_in[30]);
  or (_09074_, _09563_, _09562_);
  nor (_09564_, _09477_, _08274_);
  and (_09565_, _09477_, _08558_);
  nor (_09566_, _09565_, _09564_);
  nor (_09567_, _09566_, _09475_);
  and (_09568_, _09475_, word_in[15]);
  or (_09569_, _09568_, _09567_);
  and (_09570_, _09569_, _09474_);
  and (_09571_, _09473_, _08566_);
  or (_09572_, _09571_, _09570_);
  and (_09573_, _09572_, _09471_);
  and (_09574_, _09470_, word_in[31]);
  or (_09077_, _09574_, _09573_);
  and (_09575_, _06400_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_09576_, _07977_, _06390_);
  and (_09577_, _09576_, _06398_);
  or (_09578_, _09577_, _09575_);
  and (_09087_, _09578_, _06071_);
  and (_09579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_09580_, _09579_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_09581_, _09580_, _07900_);
  and (_09582_, _07904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_09583_, _09582_, _09005_);
  or (_09584_, _09583_, _09581_);
  and (_09585_, _09005_, _09579_);
  or (_09586_, _09585_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_09587_, _09586_, _06071_);
  and (_09148_, _09587_, _09584_);
  and (_09588_, _08546_, _08460_);
  and (_09589_, _09588_, _08344_);
  not (_09590_, _09589_);
  and (_09591_, _08550_, _08621_);
  not (_09592_, _09591_);
  not (_09593_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_09594_, _08555_, _08318_);
  and (_09595_, _09594_, _09049_);
  nor (_09596_, _09595_, _09593_);
  and (_09597_, _09595_, word_in[0]);
  or (_09598_, _09597_, _09596_);
  and (_09599_, _09598_, _09592_);
  and (_09600_, _09591_, word_in[8]);
  or (_09601_, _09600_, _09599_);
  and (_09602_, _09601_, _09590_);
  and (_09603_, _08539_, _08474_);
  and (_09604_, _09603_, _08479_);
  and (_09605_, _09604_, _08308_);
  and (_09606_, _09589_, _09168_);
  or (_09607_, _09606_, _09605_);
  or (_09608_, _09607_, _09602_);
  not (_09609_, _09605_);
  or (_09610_, _09609_, _09043_);
  and (_09161_, _09610_, _09608_);
  not (_09611_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_09612_, _09595_, _09611_);
  and (_09613_, _09595_, word_in[1]);
  or (_09614_, _09613_, _09612_);
  and (_09615_, _09614_, _09592_);
  and (_09616_, _09591_, word_in[9]);
  or (_09617_, _09616_, _09615_);
  and (_09618_, _09617_, _09590_);
  and (_09619_, _09589_, _09194_);
  or (_09620_, _09619_, _09605_);
  or (_09621_, _09620_, _09618_);
  or (_09622_, _09609_, _09075_);
  and (_09164_, _09622_, _09621_);
  not (_09623_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_09624_, _09595_, _09623_);
  and (_09625_, _09595_, word_in[2]);
  or (_09626_, _09625_, _09624_);
  and (_09627_, _09626_, _09592_);
  and (_09628_, _09591_, word_in[10]);
  or (_09629_, _09628_, _09627_);
  and (_09630_, _09629_, _09590_);
  and (_09631_, _09589_, _09217_);
  or (_09632_, _09631_, _09605_);
  or (_09633_, _09632_, _09630_);
  and (_09634_, _08539_, word_in[26]);
  or (_09635_, _09609_, _09634_);
  and (_14028_, _09635_, _09633_);
  not (_09636_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_09637_, _09595_, _09636_);
  and (_09638_, _09595_, word_in[3]);
  or (_09639_, _09638_, _09637_);
  and (_09640_, _09639_, _09592_);
  and (_09641_, _09591_, word_in[11]);
  or (_09642_, _09641_, _09640_);
  and (_09643_, _09642_, _09590_);
  and (_09644_, _09589_, _09113_);
  or (_09645_, _09644_, _09605_);
  or (_09646_, _09645_, _09643_);
  or (_09647_, _09609_, _09103_);
  and (_14029_, _09647_, _09646_);
  not (_09648_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_09649_, _09595_, _09648_);
  and (_09650_, _09595_, word_in[4]);
  or (_09651_, _09650_, _09649_);
  or (_09652_, _09651_, _09591_);
  or (_09653_, _09592_, word_in[12]);
  and (_09654_, _09653_, _09652_);
  and (_09655_, _09654_, _09590_);
  and (_09656_, _09589_, _09287_);
  or (_09657_, _09656_, _09605_);
  or (_09658_, _09657_, _09655_);
  and (_09659_, _08539_, word_in[28]);
  or (_09660_, _09609_, _09659_);
  and (_14030_, _09660_, _09658_);
  not (_09661_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09662_, _09595_, _09661_);
  and (_09663_, _09595_, word_in[5]);
  or (_09664_, _09663_, _09662_);
  and (_09665_, _09664_, _09592_);
  and (_09666_, _09591_, word_in[13]);
  or (_09667_, _09666_, _09665_);
  and (_09668_, _09667_, _09590_);
  and (_09669_, _09589_, _09305_);
  or (_09670_, _09669_, _09605_);
  or (_09671_, _09670_, _09668_);
  or (_09672_, _09609_, _09140_);
  and (_14031_, _09672_, _09671_);
  not (_09673_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09674_, _09595_, _09673_);
  and (_09675_, _09595_, word_in[6]);
  or (_09676_, _09675_, _09674_);
  and (_09677_, _09676_, _09592_);
  and (_09678_, _09591_, word_in[14]);
  or (_09679_, _09678_, _09677_);
  and (_09680_, _09679_, _09590_);
  and (_09681_, _09589_, _09322_);
  or (_09682_, _09681_, _09605_);
  or (_09683_, _09682_, _09680_);
  and (_09684_, _08539_, word_in[30]);
  or (_09685_, _09609_, _09684_);
  and (_09176_, _09685_, _09683_);
  nor (_09686_, _09595_, _08390_);
  and (_09687_, _09595_, word_in[7]);
  or (_09688_, _09687_, _09686_);
  and (_09689_, _09688_, _09592_);
  and (_09690_, _09591_, word_in[15]);
  or (_09691_, _09690_, _09689_);
  and (_09692_, _09691_, _09590_);
  and (_09693_, _09589_, _08566_);
  or (_09694_, _09693_, _09605_);
  or (_09695_, _09694_, _09692_);
  or (_09696_, _09609_, _08540_);
  and (_09179_, _09696_, _09695_);
  nor (_09697_, _06527_, _06146_);
  nor (_09698_, _05705_, _05865_);
  and (_09699_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_09700_, _09699_, _09698_);
  not (_09701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_09702_, _05696_, _09701_);
  and (_09703_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_09704_, _09703_, _09702_);
  and (_09705_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_09706_, _05718_, _05862_);
  nor (_09707_, _09706_, _09705_);
  and (_09708_, _09707_, _09704_);
  and (_09709_, _09708_, _09700_);
  and (_09710_, _06527_, _05811_);
  not (_09711_, _09710_);
  nor (_09712_, _09711_, _09709_);
  nor (_09713_, _09712_, _09697_);
  nor (_09186_, _09713_, rst);
  and (_09714_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_09715_, _06993_, _06400_);
  and (_09716_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_09717_, _09716_, _09345_);
  or (_09718_, _09717_, _09715_);
  or (_09719_, _09718_, _09714_);
  and (_09193_, _09719_, _06071_);
  and (_09235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06071_);
  and (_09720_, _09604_, _08344_);
  not (_09721_, _09720_);
  and (_09722_, _09588_, _08310_);
  not (_09723_, _09722_);
  or (_09724_, _09723_, _09168_);
  and (_09725_, _09173_, _08346_);
  not (_09726_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_09727_, _09594_, _09177_);
  nor (_09728_, _09727_, _09726_);
  and (_09729_, _09727_, _09056_);
  or (_09730_, _09729_, _09728_);
  or (_09731_, _09730_, _09725_);
  not (_09732_, _09725_);
  or (_09733_, _09732_, word_in[8]);
  and (_09734_, _09733_, _09731_);
  or (_09735_, _09734_, _09722_);
  and (_09736_, _09735_, _09724_);
  and (_09737_, _09736_, _09721_);
  and (_09738_, _09720_, word_in[24]);
  or (_09253_, _09738_, _09737_);
  or (_09739_, _09723_, _09194_);
  not (_09740_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09741_, _09727_, _09740_);
  and (_09742_, _09727_, _09080_);
  or (_09743_, _09742_, _09741_);
  or (_09744_, _09743_, _09725_);
  or (_09745_, _09732_, word_in[9]);
  and (_09746_, _09745_, _09744_);
  or (_09747_, _09746_, _09722_);
  and (_09748_, _09747_, _09739_);
  or (_09749_, _09748_, _09720_);
  or (_09750_, _09721_, word_in[25]);
  and (_09257_, _09750_, _09749_);
  and (_09751_, _09727_, _09210_);
  not (_09752_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09753_, _09727_, _09752_);
  nor (_09754_, _09753_, _09751_);
  nor (_09755_, _09754_, _09725_);
  and (_09756_, _09725_, word_in[10]);
  or (_09757_, _09756_, _09755_);
  and (_09758_, _09757_, _09723_);
  and (_09759_, _09722_, _09217_);
  or (_09760_, _09759_, _09720_);
  or (_09761_, _09760_, _09758_);
  or (_09762_, _09721_, word_in[26]);
  and (_09261_, _09762_, _09761_);
  or (_09763_, _09723_, _09113_);
  not (_09764_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09765_, _09727_, _09764_);
  and (_09766_, _09727_, _09260_);
  or (_09767_, _09766_, _09765_);
  or (_09768_, _09767_, _09725_);
  or (_09769_, _09732_, word_in[11]);
  and (_09770_, _09769_, _09768_);
  or (_09771_, _09770_, _09722_);
  and (_09772_, _09771_, _09763_);
  or (_09773_, _09772_, _09720_);
  or (_09774_, _09721_, word_in[27]);
  and (_09266_, _09774_, _09773_);
  and (_09775_, _09727_, _09277_);
  not (_09776_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09777_, _09727_, _09776_);
  nor (_09778_, _09777_, _09775_);
  nor (_09779_, _09778_, _09725_);
  and (_09780_, _09725_, word_in[12]);
  or (_09781_, _09780_, _09779_);
  and (_09782_, _09781_, _09723_);
  and (_09783_, _09722_, _09287_);
  or (_09784_, _09783_, _09782_);
  and (_09785_, _09784_, _09721_);
  and (_09786_, _09720_, word_in[28]);
  or (_09270_, _09786_, _09785_);
  not (_09787_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09788_, _09727_, _09787_);
  and (_09789_, _09727_, _09297_);
  or (_09790_, _09789_, _09788_);
  or (_09791_, _09790_, _09725_);
  or (_09792_, _09732_, word_in[13]);
  and (_09793_, _09792_, _09791_);
  or (_09794_, _09793_, _09722_);
  or (_09795_, _09723_, _09305_);
  and (_09796_, _09795_, _09794_);
  or (_09797_, _09796_, _09720_);
  or (_09798_, _09721_, word_in[29]);
  and (_09274_, _09798_, _09797_);
  or (_09799_, _09723_, _09322_);
  not (_09800_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09801_, _09727_, _09800_);
  and (_09802_, _09727_, _09315_);
  or (_09803_, _09802_, _09801_);
  or (_09804_, _09803_, _09725_);
  nand (_09805_, _09725_, _09556_);
  and (_09806_, _09805_, _09804_);
  or (_09807_, _09806_, _09722_);
  and (_09808_, _09807_, _09799_);
  or (_09809_, _09808_, _09720_);
  or (_09810_, _09721_, word_in[30]);
  and (_09278_, _09810_, _09809_);
  or (_09811_, _09723_, _08566_);
  nor (_09812_, _09727_, _08262_);
  and (_09813_, _09727_, _08558_);
  or (_09814_, _09813_, _09812_);
  or (_09815_, _09814_, _09725_);
  or (_09816_, _09732_, word_in[15]);
  and (_09817_, _09816_, _09815_);
  or (_09818_, _09817_, _09722_);
  and (_09819_, _09818_, _09811_);
  or (_09820_, _09819_, _09720_);
  or (_09821_, _09721_, word_in[31]);
  and (_09281_, _09821_, _09820_);
  and (_09822_, _09588_, _08328_);
  not (_09823_, _09822_);
  and (_09824_, _09361_, _08346_);
  not (_09825_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_09826_, _09365_, _08318_);
  nor (_09827_, _09826_, _09825_);
  and (_09828_, _09826_, _09056_);
  nor (_09829_, _09828_, _09827_);
  nor (_09830_, _09829_, _09824_);
  and (_09831_, _09824_, word_in[8]);
  or (_09832_, _09831_, _09830_);
  and (_09833_, _09832_, _09823_);
  and (_09834_, _09604_, _08310_);
  and (_09835_, _09822_, _09168_);
  or (_09836_, _09835_, _09834_);
  or (_09837_, _09836_, _09833_);
  not (_09838_, _09834_);
  or (_09839_, _09838_, word_in[24]);
  and (_09356_, _09839_, _09837_);
  or (_09840_, _09823_, _09194_);
  not (_09841_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_09842_, _09826_, _09841_);
  and (_09843_, _09826_, _09080_);
  or (_09844_, _09843_, _09842_);
  or (_09845_, _09844_, _09824_);
  not (_09846_, _09824_);
  or (_09847_, _09846_, word_in[9]);
  and (_09848_, _09847_, _09845_);
  or (_09849_, _09848_, _09822_);
  and (_09850_, _09849_, _09840_);
  or (_09851_, _09850_, _09834_);
  or (_09852_, _09838_, word_in[25]);
  and (_09360_, _09852_, _09851_);
  not (_09853_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_09854_, _09826_, _09853_);
  and (_09855_, _09826_, _09210_);
  or (_09856_, _09855_, _09854_);
  or (_09857_, _09856_, _09824_);
  or (_09858_, _09846_, word_in[10]);
  and (_09859_, _09858_, _09857_);
  or (_09860_, _09859_, _09822_);
  or (_09861_, _09823_, _09217_);
  and (_09862_, _09861_, _09860_);
  or (_09863_, _09862_, _09834_);
  or (_09864_, _09838_, word_in[26]);
  and (_09363_, _09864_, _09863_);
  not (_09865_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_09866_, _09826_, _09865_);
  and (_09867_, _09826_, _09260_);
  or (_09868_, _09867_, _09866_);
  or (_09869_, _09868_, _09824_);
  or (_09870_, _09846_, word_in[11]);
  and (_09871_, _09870_, _09869_);
  or (_09872_, _09871_, _09822_);
  or (_09873_, _09823_, _09113_);
  and (_09874_, _09873_, _09872_);
  or (_09875_, _09874_, _09834_);
  or (_09876_, _09838_, word_in[27]);
  and (_09366_, _09876_, _09875_);
  and (_09877_, _09826_, _09277_);
  not (_09878_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_09879_, _09826_, _09878_);
  nor (_09880_, _09879_, _09877_);
  nor (_09881_, _09880_, _09824_);
  and (_09882_, _09824_, word_in[12]);
  or (_09883_, _09882_, _09881_);
  and (_09884_, _09883_, _09823_);
  and (_09886_, _09822_, _09287_);
  or (_09887_, _09886_, _09834_);
  or (_09888_, _09887_, _09884_);
  or (_09890_, _09838_, word_in[28]);
  and (_09371_, _09890_, _09888_);
  not (_09891_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09893_, _09826_, _09891_);
  and (_09894_, _09826_, _09297_);
  or (_09896_, _09894_, _09893_);
  or (_09897_, _09896_, _09824_);
  or (_09899_, _09846_, word_in[13]);
  and (_09900_, _09899_, _09897_);
  or (_09901_, _09900_, _09822_);
  or (_09903_, _09823_, _09305_);
  and (_09904_, _09903_, _09901_);
  or (_09906_, _09904_, _09834_);
  or (_09908_, _09838_, word_in[29]);
  and (_09373_, _09908_, _09906_);
  and (_09909_, _09826_, _09315_);
  not (_09910_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09911_, _09826_, _09910_);
  nor (_09912_, _09911_, _09909_);
  nor (_09913_, _09912_, _09824_);
  and (_09914_, _09824_, word_in[14]);
  or (_09915_, _09914_, _09913_);
  and (_09916_, _09915_, _09823_);
  and (_09917_, _09822_, _09322_);
  or (_09918_, _09917_, _09834_);
  or (_09919_, _09918_, _09916_);
  or (_09920_, _09838_, word_in[30]);
  and (_09376_, _09920_, _09919_);
  nor (_09921_, _09826_, _08384_);
  and (_09922_, _09826_, _08558_);
  nor (_09923_, _09922_, _09921_);
  nor (_09924_, _09923_, _09824_);
  and (_09925_, _09824_, word_in[15]);
  or (_09926_, _09925_, _09924_);
  and (_09927_, _09926_, _09823_);
  and (_09928_, _09822_, _08566_);
  or (_09929_, _09928_, _09834_);
  or (_09930_, _09929_, _09927_);
  or (_09931_, _09838_, word_in[31]);
  and (_09379_, _09931_, _09930_);
  and (_09932_, _09588_, _08308_);
  and (_09933_, _08551_, _08346_);
  and (_09934_, _09594_, _08554_);
  and (_09935_, _09934_, _09056_);
  not (_09936_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_09937_, _09934_, _09936_);
  nor (_09938_, _09937_, _09935_);
  nor (_09939_, _09938_, _09933_);
  and (_09940_, _09933_, word_in[8]);
  or (_09941_, _09940_, _09939_);
  or (_09942_, _09941_, _09932_);
  and (_09943_, _08539_, _08644_);
  not (_09944_, _09943_);
  not (_09945_, _09932_);
  or (_09946_, _09945_, _09168_);
  and (_09947_, _09946_, _09944_);
  and (_09948_, _09947_, _09942_);
  and (_09949_, _09043_, _08644_);
  or (_14032_, _09949_, _09948_);
  not (_09950_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_09951_, _09934_, _09950_);
  and (_09952_, _09934_, _09080_);
  or (_09953_, _09952_, _09951_);
  or (_09954_, _09953_, _09933_);
  not (_09955_, _09933_);
  or (_09956_, _09955_, word_in[9]);
  and (_09957_, _09956_, _09954_);
  or (_09958_, _09957_, _09932_);
  or (_09959_, _09945_, _09194_);
  and (_09960_, _09959_, _09958_);
  or (_09961_, _09960_, _09943_);
  or (_09962_, _09944_, word_in[25]);
  and (_14033_, _09962_, _09961_);
  and (_09963_, _09634_, _08644_);
  and (_09964_, _09934_, _09210_);
  not (_09965_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_09966_, _09934_, _09965_);
  nor (_09967_, _09966_, _09964_);
  nor (_09968_, _09967_, _09933_);
  and (_09969_, _09933_, word_in[10]);
  or (_09970_, _09969_, _09968_);
  and (_09971_, _09970_, _09945_);
  and (_09972_, _09932_, _09217_);
  or (_09973_, _09972_, _09971_);
  and (_09974_, _09973_, _09944_);
  or (_14034_, _09974_, _09963_);
  and (_09975_, _09103_, _08644_);
  not (_09976_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_09977_, _09934_, _09976_);
  and (_09978_, _09934_, _09260_);
  or (_09979_, _09978_, _09977_);
  or (_09980_, _09979_, _09933_);
  or (_09981_, _09955_, word_in[11]);
  and (_09982_, _09981_, _09980_);
  or (_09984_, _09982_, _09932_);
  or (_09986_, _09945_, _09113_);
  and (_09987_, _09986_, _09944_);
  and (_09988_, _09987_, _09984_);
  or (_14035_, _09988_, _09975_);
  and (_09990_, _09943_, word_in[28]);
  not (_09991_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_09992_, _09934_, _09991_);
  and (_09993_, _09934_, _09277_);
  or (_09995_, _09993_, _09992_);
  or (_09997_, _09995_, _09933_);
  or (_09998_, _09955_, word_in[12]);
  and (_09999_, _09998_, _09997_);
  or (_10000_, _09999_, _09932_);
  or (_10002_, _09945_, _09287_);
  and (_10003_, _10002_, _09944_);
  and (_10004_, _10003_, _10000_);
  or (_14036_, _10004_, _09990_);
  and (_10006_, _09140_, _08644_);
  and (_10007_, _09934_, _09297_);
  not (_10008_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_10010_, _09934_, _10008_);
  nor (_10011_, _10010_, _10007_);
  nor (_10012_, _10011_, _09933_);
  and (_10013_, _09933_, word_in[13]);
  or (_10014_, _10013_, _10012_);
  and (_10015_, _10014_, _09945_);
  and (_10016_, _09932_, _09305_);
  or (_10017_, _10016_, _10015_);
  and (_10018_, _10017_, _09944_);
  or (_14037_, _10018_, _10006_);
  not (_10019_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_10020_, _09934_, _10019_);
  and (_10021_, _09934_, _09315_);
  or (_10022_, _10021_, _10020_);
  or (_10023_, _10022_, _09933_);
  nand (_10024_, _09933_, _09556_);
  and (_10025_, _10024_, _10023_);
  or (_10026_, _10025_, _09932_);
  or (_10027_, _09945_, _09322_);
  and (_10028_, _10027_, _09944_);
  and (_10029_, _10028_, _10026_);
  and (_10030_, _09943_, word_in[30]);
  or (_14038_, _10030_, _10029_);
  and (_10031_, _09934_, _08558_);
  nor (_10033_, _09934_, _08268_);
  nor (_10034_, _10033_, _10031_);
  nor (_10035_, _10034_, _09933_);
  and (_10036_, _09933_, word_in[15]);
  or (_10037_, _10036_, _10035_);
  and (_10038_, _10037_, _09945_);
  and (_10039_, _09932_, _08566_);
  or (_10040_, _10039_, _10038_);
  and (_10041_, _10040_, _09944_);
  and (_10042_, _09943_, word_in[31]);
  or (_14039_, _10042_, _10041_);
  and (_10043_, _08539_, _08482_);
  and (_10044_, _10043_, _08308_);
  not (_10045_, _10044_);
  and (_10046_, _08545_, _08428_);
  not (_10047_, _10046_);
  or (_10048_, _10047_, word_in[16]);
  and (_10049_, _08550_, _08319_);
  not (_10050_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10051_, _08317_, _08184_);
  and (_10052_, _08555_, _10051_);
  and (_10053_, _10052_, _09049_);
  nor (_10054_, _10053_, _10050_);
  and (_10055_, _10053_, _09056_);
  or (_10056_, _10055_, _10054_);
  or (_10057_, _10056_, _10049_);
  not (_10058_, _10049_);
  or (_10059_, _10058_, word_in[8]);
  and (_10060_, _10059_, _10057_);
  or (_10061_, _10060_, _10046_);
  and (_10062_, _10061_, _10048_);
  and (_10063_, _10062_, _10045_);
  and (_10064_, _10044_, word_in[24]);
  or (_09547_, _10064_, _10063_);
  and (_10065_, _10046_, word_in[17]);
  not (_10066_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_10067_, _10053_, _10066_);
  and (_10068_, _10053_, word_in[1]);
  or (_10069_, _10068_, _10067_);
  and (_10070_, _10069_, _10058_);
  and (_10071_, _10049_, word_in[9]);
  or (_10072_, _10071_, _10070_);
  and (_10073_, _10072_, _10047_);
  or (_10074_, _10073_, _10065_);
  and (_10075_, _10074_, _10045_);
  and (_10076_, _10044_, word_in[25]);
  or (_09551_, _10076_, _10075_);
  and (_10078_, _10046_, word_in[18]);
  not (_10079_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_10080_, _10053_, _10079_);
  and (_10082_, _10053_, word_in[2]);
  or (_10083_, _10082_, _10080_);
  and (_10084_, _10083_, _10058_);
  and (_10085_, _10049_, word_in[10]);
  or (_10087_, _10085_, _10084_);
  and (_10088_, _10087_, _10047_);
  or (_10089_, _10088_, _10078_);
  and (_10090_, _10089_, _10045_);
  and (_10092_, _10044_, word_in[26]);
  or (_14040_, _10092_, _10090_);
  and (_10093_, _10046_, word_in[19]);
  not (_10095_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_10096_, _10053_, _10095_);
  and (_10097_, _10053_, word_in[3]);
  or (_10098_, _10097_, _10096_);
  and (_10100_, _10098_, _10058_);
  and (_10101_, _10049_, word_in[11]);
  or (_10102_, _10101_, _10100_);
  and (_10103_, _10102_, _10047_);
  or (_10105_, _10103_, _10093_);
  and (_10107_, _10105_, _10045_);
  and (_10108_, _10044_, word_in[27]);
  or (_14041_, _10108_, _10107_);
  and (_10109_, _10046_, word_in[20]);
  not (_10110_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_10111_, _10053_, _10110_);
  and (_10112_, _10053_, word_in[4]);
  or (_10113_, _10112_, _10111_);
  and (_10114_, _10113_, _10058_);
  and (_10115_, _10049_, word_in[12]);
  or (_10116_, _10115_, _10114_);
  and (_10117_, _10116_, _10047_);
  or (_10118_, _10117_, _10109_);
  and (_10119_, _10118_, _10045_);
  and (_10120_, _10044_, word_in[28]);
  or (_14042_, _10120_, _10119_);
  not (_10121_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_10122_, _10053_, _10121_);
  and (_10123_, _10053_, word_in[5]);
  or (_10124_, _10123_, _10122_);
  and (_10125_, _10124_, _10058_);
  and (_10126_, _10049_, word_in[13]);
  or (_10127_, _10126_, _10125_);
  and (_10128_, _10127_, _10047_);
  and (_10129_, _10046_, word_in[21]);
  or (_10130_, _10129_, _10128_);
  and (_10131_, _10130_, _10045_);
  and (_10132_, _10044_, word_in[29]);
  or (_14043_, _10132_, _10131_);
  and (_10133_, _10046_, word_in[22]);
  not (_10134_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_10135_, _10053_, _10134_);
  and (_10136_, _10053_, word_in[6]);
  or (_10137_, _10136_, _10135_);
  and (_10138_, _10137_, _10058_);
  and (_10139_, _10049_, word_in[14]);
  or (_10140_, _10139_, _10138_);
  and (_10141_, _10140_, _10047_);
  or (_10142_, _10141_, _10133_);
  and (_10143_, _10142_, _10045_);
  and (_10144_, _10044_, word_in[30]);
  or (_14044_, _10144_, _10143_);
  and (_10145_, _10046_, word_in[23]);
  nor (_10146_, _10053_, _08365_);
  and (_10147_, _10053_, word_in[7]);
  or (_10148_, _10147_, _10146_);
  and (_10149_, _10148_, _10058_);
  and (_10150_, _10049_, word_in[15]);
  or (_10151_, _10150_, _10149_);
  and (_10152_, _10151_, _10047_);
  or (_10153_, _10152_, _10145_);
  and (_10154_, _10153_, _10045_);
  and (_10155_, _10044_, word_in[31]);
  or (_14045_, _10155_, _10154_);
  and (_10156_, _09169_, _08420_);
  not (_10157_, _10156_);
  and (_10158_, _09173_, _08323_);
  and (_10159_, _10052_, _09177_);
  and (_10160_, _10159_, _09056_);
  not (_10161_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_10162_, _10159_, _10161_);
  nor (_10163_, _10162_, _10160_);
  nor (_10164_, _10163_, _10158_);
  and (_10165_, _10158_, word_in[8]);
  or (_10166_, _10165_, _10164_);
  and (_10167_, _10166_, _10157_);
  and (_10168_, _10043_, _08344_);
  and (_10169_, _10156_, _09168_);
  or (_10171_, _10169_, _10168_);
  or (_10172_, _10171_, _10167_);
  not (_10173_, _10168_);
  or (_10175_, _10173_, _09043_);
  and (_14046_, _10175_, _10172_);
  not (_10177_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_10179_, _10159_, _10177_);
  and (_10181_, _10159_, _09080_);
  or (_10182_, _10181_, _10179_);
  or (_10183_, _10182_, _10158_);
  not (_10185_, _10158_);
  or (_10186_, _10185_, word_in[9]);
  and (_10188_, _10186_, _10183_);
  or (_10189_, _10188_, _10156_);
  or (_10191_, _10157_, _09194_);
  and (_10192_, _10191_, _10173_);
  and (_10193_, _10192_, _10189_);
  and (_10194_, _10168_, _09075_);
  or (_14047_, _10194_, _10193_);
  not (_10195_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_10196_, _10159_, _10195_);
  and (_10197_, _10159_, _09210_);
  or (_10198_, _10197_, _10196_);
  or (_10199_, _10198_, _10158_);
  or (_10200_, _10185_, word_in[10]);
  and (_10201_, _10200_, _10199_);
  or (_10202_, _10201_, _10156_);
  or (_10203_, _10157_, _09217_);
  and (_10204_, _10203_, _10173_);
  and (_10205_, _10204_, _10202_);
  and (_10206_, _10168_, _09634_);
  or (_14048_, _10206_, _10205_);
  and (_10207_, _10159_, _09260_);
  not (_10208_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_10209_, _10159_, _10208_);
  nor (_10210_, _10209_, _10207_);
  nor (_10211_, _10210_, _10158_);
  and (_10212_, _10158_, word_in[11]);
  or (_10213_, _10212_, _10211_);
  and (_10214_, _10213_, _10157_);
  and (_10215_, _10156_, _09113_);
  or (_10216_, _10215_, _10168_);
  or (_10217_, _10216_, _10214_);
  or (_10218_, _10173_, _09103_);
  and (_14049_, _10218_, _10217_);
  and (_10219_, _10159_, _09277_);
  not (_10220_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_10221_, _10159_, _10220_);
  nor (_10222_, _10221_, _10219_);
  nor (_10223_, _10222_, _10158_);
  and (_10224_, _10158_, word_in[12]);
  or (_10225_, _10224_, _10223_);
  and (_10226_, _10225_, _10157_);
  and (_10227_, _10156_, _09287_);
  or (_10228_, _10227_, _10168_);
  or (_10229_, _10228_, _10226_);
  or (_10230_, _10173_, _09659_);
  and (_14050_, _10230_, _10229_);
  and (_10231_, _10159_, _09297_);
  not (_10232_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_10233_, _10159_, _10232_);
  nor (_10234_, _10233_, _10231_);
  nor (_10235_, _10234_, _10158_);
  and (_10236_, _10158_, word_in[13]);
  or (_10237_, _10236_, _10235_);
  and (_10238_, _10237_, _10157_);
  and (_10239_, _10156_, _09305_);
  or (_10240_, _10239_, _10168_);
  or (_10241_, _10240_, _10238_);
  or (_10242_, _10173_, _09140_);
  and (_14051_, _10242_, _10241_);
  and (_10243_, _10159_, _09315_);
  not (_10244_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_10245_, _10159_, _10244_);
  nor (_10246_, _10245_, _10243_);
  nor (_10247_, _10246_, _10158_);
  and (_10248_, _10158_, word_in[14]);
  or (_10249_, _10248_, _10247_);
  and (_10250_, _10249_, _10157_);
  and (_10251_, _10156_, _09322_);
  or (_10252_, _10251_, _10168_);
  or (_10253_, _10252_, _10250_);
  or (_10254_, _10173_, _09684_);
  and (_14052_, _10254_, _10253_);
  and (_10255_, _10159_, _08558_);
  nor (_10256_, _10159_, _08282_);
  nor (_10257_, _10256_, _10255_);
  nor (_10258_, _10257_, _10158_);
  and (_10259_, _10158_, word_in[15]);
  or (_10260_, _10259_, _10258_);
  and (_10261_, _10260_, _10157_);
  and (_10262_, _10156_, _08566_);
  or (_10263_, _10262_, _10168_);
  or (_10264_, _10263_, _10261_);
  or (_10265_, _10173_, _08540_);
  and (_14053_, _10265_, _10264_);
  and (_10266_, _10043_, _08310_);
  and (_10267_, _09357_, _08420_);
  and (_10268_, _09361_, _08323_);
  not (_10269_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10270_, _10052_, _09365_);
  nor (_10271_, _10270_, _10269_);
  and (_10272_, _10270_, _09056_);
  or (_10273_, _10272_, _10271_);
  or (_10274_, _10273_, _10268_);
  not (_10275_, _10268_);
  or (_10276_, _10275_, word_in[8]);
  and (_10277_, _10276_, _10274_);
  or (_10278_, _10277_, _10267_);
  not (_10279_, _10267_);
  or (_10280_, _10279_, _09168_);
  and (_10281_, _10280_, _10278_);
  or (_10282_, _10281_, _10266_);
  not (_10283_, _10266_);
  or (_10284_, _10283_, word_in[24]);
  and (_14008_, _10284_, _10282_);
  not (_10285_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_10286_, _10270_, _10285_);
  and (_10287_, _10270_, _09080_);
  or (_10288_, _10287_, _10286_);
  or (_10289_, _10288_, _10268_);
  or (_10290_, _10275_, word_in[9]);
  and (_10291_, _10290_, _10289_);
  or (_10292_, _10291_, _10267_);
  or (_10293_, _10279_, _09194_);
  and (_10294_, _10293_, _10283_);
  and (_10295_, _10294_, _10292_);
  and (_10296_, _10266_, word_in[25]);
  or (_14009_, _10296_, _10295_);
  and (_10297_, _10270_, _09210_);
  not (_10298_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_10299_, _10270_, _10298_);
  nor (_10300_, _10299_, _10297_);
  nor (_10301_, _10300_, _10268_);
  and (_10302_, _10268_, word_in[10]);
  or (_10303_, _10302_, _10301_);
  and (_10304_, _10303_, _10279_);
  and (_10305_, _10267_, _09217_);
  or (_10306_, _10305_, _10266_);
  or (_10307_, _10306_, _10304_);
  or (_10308_, _10283_, word_in[26]);
  and (_14010_, _10308_, _10307_);
  and (_10309_, _10270_, _09260_);
  not (_10310_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_10311_, _10270_, _10310_);
  nor (_10312_, _10311_, _10309_);
  nor (_10313_, _10312_, _10268_);
  and (_10314_, _10268_, word_in[11]);
  or (_10315_, _10314_, _10313_);
  and (_10316_, _10315_, _10279_);
  and (_10317_, _10267_, _09113_);
  or (_10318_, _10317_, _10266_);
  or (_10319_, _10318_, _10316_);
  or (_10320_, _10283_, word_in[27]);
  and (_14011_, _10320_, _10319_);
  and (_10321_, _10267_, _09287_);
  and (_10322_, _10270_, _09277_);
  not (_10323_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_10324_, _10270_, _10323_);
  nor (_10325_, _10324_, _10322_);
  nor (_10326_, _10325_, _10268_);
  and (_10327_, _10268_, word_in[12]);
  or (_10328_, _10327_, _10326_);
  and (_10329_, _10328_, _10279_);
  or (_10330_, _10329_, _10321_);
  and (_10331_, _10330_, _10283_);
  and (_10332_, _10266_, word_in[28]);
  or (_14012_, _10332_, _10331_);
  and (_10333_, _10270_, _09297_);
  not (_10334_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_10335_, _10270_, _10334_);
  nor (_10336_, _10335_, _10333_);
  nor (_10337_, _10336_, _10268_);
  and (_10338_, _10268_, word_in[13]);
  or (_10339_, _10338_, _10337_);
  and (_10340_, _10339_, _10279_);
  and (_10341_, _10267_, _09305_);
  or (_10342_, _10341_, _10266_);
  or (_10343_, _10342_, _10340_);
  or (_10344_, _10283_, word_in[29]);
  and (_14013_, _10344_, _10343_);
  and (_10345_, _10270_, _09315_);
  not (_10346_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_10347_, _10270_, _10346_);
  nor (_10348_, _10347_, _10345_);
  nor (_10349_, _10348_, _10268_);
  and (_10350_, _10268_, word_in[14]);
  or (_10351_, _10350_, _10349_);
  and (_10352_, _10351_, _10279_);
  and (_10353_, _10267_, _09322_);
  or (_10354_, _10353_, _10266_);
  or (_10355_, _10354_, _10352_);
  or (_10356_, _10283_, word_in[30]);
  and (_14014_, _10356_, _10355_);
  nor (_10357_, _10270_, _08360_);
  and (_10358_, _10270_, _08558_);
  or (_10359_, _10358_, _10357_);
  or (_10360_, _10359_, _10268_);
  or (_10361_, _10275_, word_in[15]);
  and (_10362_, _10361_, _10360_);
  or (_10363_, _10362_, _10267_);
  or (_10364_, _10279_, _08566_);
  and (_10365_, _10364_, _10363_);
  and (_10366_, _10365_, _10283_);
  and (_10367_, _10266_, word_in[31]);
  or (_14015_, _10367_, _10366_);
  and (_10368_, _09472_, _08420_);
  not (_10369_, _10368_);
  and (_10370_, _08551_, _08323_);
  not (_10371_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_10372_, _10052_, _08554_);
  nor (_10373_, _10372_, _10371_);
  and (_10374_, _10372_, _09056_);
  or (_10375_, _10374_, _10373_);
  or (_10376_, _10375_, _10370_);
  not (_10377_, _10370_);
  or (_10378_, _10377_, word_in[8]);
  and (_10379_, _10378_, _10376_);
  and (_10380_, _10379_, _10369_);
  and (_10381_, _10043_, _08328_);
  and (_10382_, _10368_, _09168_);
  or (_10383_, _10382_, _10381_);
  or (_10384_, _10383_, _10380_);
  not (_10385_, _10381_);
  or (_10386_, _10385_, word_in[24]);
  and (_14016_, _10386_, _10384_);
  not (_10387_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_10388_, _10372_, _10387_);
  and (_10389_, _10372_, _09080_);
  or (_10390_, _10389_, _10388_);
  or (_10391_, _10390_, _10370_);
  or (_10392_, _10377_, word_in[9]);
  and (_10393_, _10392_, _10391_);
  or (_10394_, _10393_, _10368_);
  or (_10395_, _10369_, _09194_);
  and (_10396_, _10395_, _10394_);
  or (_10397_, _10396_, _10381_);
  or (_10398_, _10385_, word_in[25]);
  and (_14017_, _10398_, _10397_);
  not (_10399_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_10400_, _10372_, _10399_);
  and (_10401_, _10372_, _09210_);
  or (_10402_, _10401_, _10400_);
  or (_10403_, _10402_, _10370_);
  or (_10404_, _10377_, word_in[10]);
  and (_10405_, _10404_, _10403_);
  or (_10406_, _10405_, _10368_);
  or (_10407_, _10369_, _09217_);
  and (_10408_, _10407_, _10385_);
  and (_10409_, _10408_, _10406_);
  and (_10410_, _10381_, _09634_);
  or (_14018_, _10410_, _10409_);
  and (_10411_, _10372_, _09260_);
  not (_10412_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_10413_, _10372_, _10412_);
  nor (_10414_, _10413_, _10411_);
  nor (_10415_, _10414_, _10370_);
  and (_10416_, _10370_, word_in[11]);
  or (_10417_, _10416_, _10415_);
  and (_10418_, _10417_, _10369_);
  and (_10420_, _10368_, _09113_);
  or (_10421_, _10420_, _10381_);
  or (_10422_, _10421_, _10418_);
  or (_10423_, _10385_, _09103_);
  and (_14019_, _10423_, _10422_);
  not (_10425_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_10426_, _10372_, _10425_);
  and (_10428_, _10372_, _09277_);
  or (_10429_, _10428_, _10426_);
  or (_10431_, _10429_, _10370_);
  or (_10432_, _10377_, word_in[12]);
  and (_10434_, _10432_, _10431_);
  or (_10435_, _10434_, _10368_);
  or (_10436_, _10369_, _09287_);
  and (_10437_, _10436_, _10385_);
  and (_10438_, _10437_, _10435_);
  and (_10439_, _10381_, _09659_);
  or (_14020_, _10439_, _10438_);
  and (_10440_, _10372_, _09297_);
  not (_10441_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_10442_, _10372_, _10441_);
  nor (_10443_, _10442_, _10440_);
  nor (_10444_, _10443_, _10370_);
  and (_10445_, _10370_, word_in[13]);
  or (_10446_, _10445_, _10444_);
  and (_10447_, _10446_, _10369_);
  and (_10448_, _10368_, _09305_);
  or (_10450_, _10448_, _10381_);
  or (_10451_, _10450_, _10447_);
  or (_10452_, _10385_, _09140_);
  and (_14021_, _10452_, _10451_);
  and (_10453_, _10372_, _09315_);
  not (_10454_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_10455_, _10372_, _10454_);
  nor (_10456_, _10455_, _10453_);
  nor (_10457_, _10456_, _10370_);
  and (_10458_, _10370_, word_in[14]);
  or (_10460_, _10458_, _10457_);
  and (_10461_, _10460_, _10369_);
  and (_10462_, _10368_, _09322_);
  or (_10463_, _10462_, _10381_);
  or (_10464_, _10463_, _10461_);
  or (_10465_, _10385_, _09684_);
  and (_14022_, _10465_, _10464_);
  nor (_10466_, _10372_, _08299_);
  and (_10467_, _10372_, _08558_);
  or (_10468_, _10467_, _10466_);
  or (_10469_, _10468_, _10370_);
  or (_10470_, _10377_, word_in[15]);
  and (_10471_, _10470_, _10469_);
  or (_10472_, _10471_, _10368_);
  or (_10473_, _10369_, _08566_);
  and (_10474_, _10473_, _10385_);
  and (_10475_, _10474_, _10472_);
  and (_10476_, _10381_, _08540_);
  or (_14023_, _10476_, _10475_);
  and (_10477_, _08547_, _08344_);
  not (_10478_, _10477_);
  and (_10479_, _08522_, _08310_);
  and (_10481_, _08550_, _10479_);
  not (_10483_, _10481_);
  not (_10484_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_10485_, _09049_, _08556_);
  nor (_10486_, _10485_, _10484_);
  and (_10487_, _10485_, word_in[0]);
  or (_10488_, _10487_, _10486_);
  and (_10489_, _10488_, _10483_);
  and (_10490_, _10481_, word_in[8]);
  or (_10491_, _10490_, _10489_);
  and (_10492_, _10491_, _10478_);
  not (_10493_, _08479_);
  and (_10494_, _09603_, _10493_);
  and (_10495_, _10494_, _08308_);
  and (_10496_, _10477_, _09168_);
  or (_10497_, _10496_, _10495_);
  or (_10498_, _10497_, _10492_);
  not (_10499_, _10495_);
  or (_10500_, _10499_, _09043_);
  and (_09885_, _10500_, _10498_);
  not (_10501_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_10502_, _10485_, _10501_);
  and (_10503_, _10485_, word_in[1]);
  or (_10504_, _10503_, _10502_);
  and (_10505_, _10504_, _10483_);
  and (_10506_, _10481_, word_in[9]);
  or (_10507_, _10506_, _10505_);
  and (_10508_, _10507_, _10478_);
  and (_10509_, _10477_, _09194_);
  or (_10510_, _10509_, _10495_);
  or (_10511_, _10510_, _10508_);
  or (_10512_, _10499_, _09075_);
  and (_09889_, _10512_, _10511_);
  not (_10513_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_10514_, _10485_, _10513_);
  and (_10515_, _10485_, word_in[2]);
  or (_10516_, _10515_, _10514_);
  and (_10517_, _10516_, _10483_);
  and (_10518_, _10481_, word_in[10]);
  or (_10519_, _10518_, _10517_);
  and (_10520_, _10519_, _10478_);
  and (_10521_, _10477_, _09217_);
  or (_10522_, _10521_, _10495_);
  or (_10523_, _10522_, _10520_);
  or (_10524_, _10499_, _09634_);
  and (_09892_, _10524_, _10523_);
  not (_10525_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_10526_, _10485_, _10525_);
  and (_10527_, _10485_, word_in[3]);
  or (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _10483_);
  and (_10530_, _10481_, word_in[11]);
  or (_10531_, _10530_, _10529_);
  and (_10532_, _10531_, _10478_);
  and (_10533_, _10477_, _09113_);
  or (_10534_, _10533_, _10495_);
  or (_10535_, _10534_, _10532_);
  or (_10536_, _10499_, _09103_);
  and (_09895_, _10536_, _10535_);
  not (_10537_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_10538_, _10485_, _10537_);
  and (_10539_, _10485_, word_in[4]);
  or (_10540_, _10539_, _10538_);
  and (_10541_, _10540_, _10483_);
  and (_10542_, _10481_, word_in[12]);
  or (_10543_, _10542_, _10541_);
  and (_10544_, _10543_, _10478_);
  and (_10545_, _10477_, _09287_);
  or (_10546_, _10545_, _10495_);
  or (_10547_, _10546_, _10544_);
  or (_10548_, _10499_, _09659_);
  and (_09898_, _10548_, _10547_);
  not (_10549_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_10550_, _10485_, _10549_);
  and (_10551_, _10485_, word_in[5]);
  or (_10552_, _10551_, _10550_);
  and (_10553_, _10552_, _10483_);
  and (_10554_, _10481_, word_in[13]);
  or (_10555_, _10554_, _10553_);
  and (_10556_, _10555_, _10478_);
  and (_10557_, _10477_, _09305_);
  or (_10558_, _10557_, _10495_);
  or (_10559_, _10558_, _10556_);
  or (_10560_, _10499_, _09140_);
  and (_09902_, _10560_, _10559_);
  not (_10561_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_10562_, _10485_, _10561_);
  and (_10563_, _10485_, word_in[6]);
  or (_10564_, _10563_, _10562_);
  and (_10565_, _10564_, _10483_);
  and (_10566_, _10481_, word_in[14]);
  or (_10567_, _10566_, _10565_);
  and (_10568_, _10567_, _10478_);
  and (_10569_, _10477_, _09322_);
  or (_10570_, _10569_, _10495_);
  or (_10571_, _10570_, _10568_);
  or (_10572_, _10499_, _09684_);
  and (_09905_, _10572_, _10571_);
  nor (_10573_, _10485_, _08402_);
  and (_10574_, _10485_, word_in[7]);
  or (_10575_, _10574_, _10573_);
  and (_10576_, _10575_, _10483_);
  and (_10577_, _10481_, word_in[15]);
  or (_10578_, _10577_, _10576_);
  and (_10579_, _10578_, _10478_);
  and (_10580_, _10477_, _08566_);
  or (_10581_, _10580_, _10495_);
  or (_10582_, _10581_, _10579_);
  or (_10583_, _10499_, _08540_);
  and (_09907_, _10583_, _10582_);
  and (_10584_, _08547_, _08310_);
  not (_10585_, _10584_);
  and (_10586_, _09173_, _08350_);
  and (_10587_, _09177_, _08556_);
  and (_10588_, _10587_, _09056_);
  not (_10589_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_10590_, _10587_, _10589_);
  nor (_10591_, _10590_, _10588_);
  nor (_10592_, _10591_, _10586_);
  and (_10593_, _10586_, word_in[8]);
  or (_10594_, _10593_, _10592_);
  and (_10595_, _10594_, _10585_);
  and (_10596_, _10494_, _08344_);
  and (_10597_, _10584_, _09168_);
  or (_10598_, _10597_, _10596_);
  or (_10599_, _10598_, _10595_);
  not (_10600_, _10596_);
  or (_10601_, _10600_, word_in[24]);
  and (_14024_, _10601_, _10599_);
  nor (_10602_, _09341_, _08865_);
  and (_10603_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_10604_, _10603_, _10602_);
  and (_09983_, _10604_, _06071_);
  or (_10605_, _10585_, _09194_);
  not (_10606_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_10607_, _10587_, _10606_);
  and (_10608_, _10587_, _09080_);
  or (_10609_, _10608_, _10607_);
  or (_10610_, _10609_, _10586_);
  not (_10611_, _10586_);
  or (_10612_, _10611_, word_in[9]);
  and (_10613_, _10612_, _10610_);
  or (_10614_, _10613_, _10584_);
  and (_10615_, _10614_, _10605_);
  and (_10616_, _10615_, _10600_);
  and (_10617_, _10596_, word_in[25]);
  or (_09985_, _10617_, _10616_);
  or (_10618_, _10611_, word_in[10]);
  not (_10619_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_10620_, _10587_, _10619_);
  and (_10621_, _10587_, _09210_);
  or (_10622_, _10621_, _10620_);
  or (_10623_, _10622_, _10586_);
  and (_10624_, _10623_, _10585_);
  and (_10625_, _10624_, _10618_);
  and (_10626_, _10584_, _09217_);
  or (_10627_, _10626_, _10596_);
  or (_10628_, _10627_, _10625_);
  or (_10629_, _10600_, word_in[26]);
  and (_09989_, _10629_, _10628_);
  and (_10630_, _10587_, _09260_);
  not (_10631_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_10632_, _10587_, _10631_);
  nor (_10633_, _10632_, _10630_);
  nor (_10634_, _10633_, _10586_);
  and (_10635_, _10586_, word_in[11]);
  or (_10636_, _10635_, _10634_);
  and (_10637_, _10636_, _10585_);
  and (_10638_, _10584_, _09113_);
  or (_10639_, _10638_, _10596_);
  or (_10640_, _10639_, _10637_);
  or (_10641_, _10600_, word_in[27]);
  and (_09994_, _10641_, _10640_);
  and (_10642_, _10587_, _09277_);
  not (_10643_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_10644_, _10587_, _10643_);
  nor (_10645_, _10644_, _10642_);
  nor (_10646_, _10645_, _10586_);
  and (_10647_, _10586_, word_in[12]);
  or (_10648_, _10647_, _10646_);
  and (_10649_, _10648_, _10585_);
  and (_10650_, _10584_, _09287_);
  or (_10651_, _10650_, _10596_);
  or (_10652_, _10651_, _10649_);
  or (_10653_, _10600_, word_in[28]);
  and (_09996_, _10653_, _10652_);
  not (_10654_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_10655_, _10587_, _10654_);
  and (_10656_, _10587_, _09297_);
  or (_10657_, _10656_, _10655_);
  or (_10658_, _10657_, _10586_);
  or (_10659_, _10611_, word_in[13]);
  and (_10660_, _10659_, _10658_);
  or (_10661_, _10660_, _10584_);
  or (_10662_, _10585_, _09305_);
  and (_10663_, _10662_, _10661_);
  or (_10664_, _10663_, _10596_);
  or (_10665_, _10600_, word_in[29]);
  and (_10001_, _10665_, _10664_);
  or (_10666_, _10585_, _09322_);
  not (_10667_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_10668_, _10587_, _10667_);
  and (_10669_, _10587_, _09315_);
  or (_10670_, _10669_, _10668_);
  or (_10671_, _10670_, _10586_);
  nand (_10672_, _10586_, _09556_);
  and (_10673_, _10672_, _10671_);
  or (_10674_, _10673_, _10584_);
  and (_10675_, _10674_, _10666_);
  or (_10676_, _10675_, _10596_);
  or (_10677_, _10600_, word_in[30]);
  and (_10005_, _10677_, _10676_);
  and (_10678_, _10587_, _08558_);
  nor (_10679_, _10587_, _08288_);
  nor (_10680_, _10679_, _10678_);
  nor (_10681_, _10680_, _10586_);
  and (_10682_, _10586_, word_in[15]);
  or (_10683_, _10682_, _10681_);
  and (_10684_, _10683_, _10585_);
  and (_10685_, _10584_, _08566_);
  or (_10686_, _10685_, _10596_);
  or (_10687_, _10686_, _10684_);
  or (_10688_, _10600_, word_in[31]);
  and (_10009_, _10688_, _10687_);
  or (_10689_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_10690_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_10691_, _06530_, _10690_);
  and (_10692_, _10691_, _06071_);
  and (_10032_, _10692_, _10689_);
  and (_10693_, _10494_, _08310_);
  not (_10694_, _10693_);
  and (_10695_, _08547_, _08328_);
  not (_10696_, _10695_);
  and (_10697_, _09361_, _08350_);
  and (_10698_, _09365_, _08532_);
  and (_10699_, _10698_, _09056_);
  not (_10700_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_10701_, _10698_, _10700_);
  nor (_10702_, _10701_, _10699_);
  nor (_10703_, _10702_, _10697_);
  and (_10704_, _10697_, word_in[8]);
  or (_10705_, _10704_, _10703_);
  and (_10706_, _10705_, _10696_);
  and (_10707_, _10695_, _09168_);
  or (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _10694_);
  and (_10710_, _10693_, word_in[24]);
  or (_10077_, _10710_, _10709_);
  and (_10711_, _10698_, _09080_);
  not (_10712_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_10713_, _10698_, _10712_);
  nor (_10714_, _10713_, _10711_);
  nor (_10715_, _10714_, _10697_);
  and (_10716_, _10697_, word_in[9]);
  or (_10717_, _10716_, _10715_);
  and (_10718_, _10717_, _10696_);
  and (_10719_, _10695_, _09194_);
  or (_10720_, _10719_, _10693_);
  or (_10721_, _10720_, _10718_);
  or (_10722_, _10694_, word_in[25]);
  and (_10081_, _10722_, _10721_);
  and (_10723_, _10698_, _09210_);
  not (_10724_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_10725_, _10698_, _10724_);
  nor (_10726_, _10725_, _10723_);
  nor (_10727_, _10726_, _10697_);
  and (_10728_, _10697_, word_in[10]);
  or (_10729_, _10728_, _10727_);
  and (_10730_, _10729_, _10696_);
  and (_10731_, _10695_, _09217_);
  or (_10732_, _10731_, _10693_);
  or (_10733_, _10732_, _10730_);
  or (_10734_, _10694_, word_in[26]);
  and (_10086_, _10734_, _10733_);
  and (_10735_, _10698_, _09260_);
  not (_10736_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_10737_, _10698_, _10736_);
  nor (_10738_, _10737_, _10735_);
  nor (_10739_, _10738_, _10697_);
  and (_10740_, _10697_, word_in[11]);
  or (_10741_, _10740_, _10739_);
  and (_10742_, _10741_, _10696_);
  and (_10743_, _10695_, _09113_);
  or (_10744_, _10743_, _10693_);
  or (_10745_, _10744_, _10742_);
  or (_10746_, _10694_, word_in[27]);
  and (_10091_, _10746_, _10745_);
  not (_10747_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_10748_, _10698_, _10747_);
  and (_10749_, _10698_, _09277_);
  or (_10750_, _10749_, _10748_);
  or (_10751_, _10750_, _10697_);
  not (_10752_, _10697_);
  or (_10753_, _10752_, word_in[12]);
  and (_10754_, _10753_, _10751_);
  or (_10755_, _10754_, _10695_);
  or (_10756_, _10696_, _09287_);
  and (_10757_, _10756_, _10755_);
  or (_10758_, _10757_, _10693_);
  or (_10759_, _10694_, word_in[28]);
  and (_10094_, _10759_, _10758_);
  and (_10760_, _10698_, _09297_);
  not (_10761_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_10762_, _10698_, _10761_);
  nor (_10763_, _10762_, _10760_);
  nor (_10764_, _10763_, _10697_);
  and (_10765_, _10697_, word_in[13]);
  or (_10766_, _10765_, _10764_);
  and (_10767_, _10766_, _10696_);
  and (_10768_, _10695_, _09305_);
  or (_10769_, _10768_, _10693_);
  or (_10770_, _10769_, _10767_);
  or (_10771_, _10694_, word_in[29]);
  and (_10099_, _10771_, _10770_);
  and (_10772_, _10698_, _09315_);
  not (_10773_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_10774_, _10698_, _10773_);
  nor (_10775_, _10774_, _10772_);
  nor (_10776_, _10775_, _10697_);
  and (_10777_, _10697_, word_in[14]);
  or (_10778_, _10777_, _10776_);
  and (_10779_, _10778_, _10696_);
  and (_10780_, _10695_, _09322_);
  or (_10781_, _10780_, _10693_);
  or (_10782_, _10781_, _10779_);
  or (_10783_, _10694_, word_in[30]);
  and (_10104_, _10783_, _10782_);
  and (_10784_, _10698_, _08558_);
  nor (_10785_, _10698_, _08397_);
  nor (_10786_, _10785_, _10784_);
  nor (_10787_, _10786_, _10697_);
  and (_10788_, _10697_, word_in[15]);
  or (_10789_, _10788_, _10787_);
  and (_10790_, _10789_, _10696_);
  and (_10791_, _10695_, _08566_);
  or (_10792_, _10791_, _10693_);
  or (_10793_, _10792_, _10790_);
  or (_10794_, _10694_, word_in[31]);
  and (_10106_, _10794_, _10793_);
  not (_10795_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_10796_, _08557_, _10795_);
  and (_10797_, _09056_, _08557_);
  or (_10798_, _10797_, _10796_);
  or (_10799_, _10798_, _08552_);
  not (_10800_, _08552_);
  or (_10801_, _10800_, word_in[8]);
  and (_10802_, _10801_, _10799_);
  or (_10803_, _10802_, _08548_);
  or (_10804_, _09168_, _08549_);
  and (_10805_, _10804_, _08544_);
  and (_10806_, _10805_, _10803_);
  and (_10807_, _08542_, word_in[24]);
  or (_10170_, _10807_, _10806_);
  and (_10808_, _08542_, word_in[25]);
  not (_10809_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_10810_, _08557_, _10809_);
  and (_10811_, _09080_, _08557_);
  or (_10812_, _10811_, _10810_);
  or (_10813_, _10812_, _08552_);
  or (_10814_, _10800_, word_in[9]);
  and (_10815_, _10814_, _10813_);
  or (_10816_, _10815_, _08548_);
  or (_10817_, _09194_, _08549_);
  and (_10818_, _10817_, _08544_);
  and (_10819_, _10818_, _10816_);
  or (_10174_, _10819_, _10808_);
  not (_10820_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_10821_, _08557_, _10820_);
  and (_10822_, _09210_, _08557_);
  or (_10823_, _10822_, _10821_);
  or (_10824_, _10823_, _08552_);
  or (_10825_, _10800_, word_in[10]);
  and (_10826_, _10825_, _10824_);
  or (_10827_, _10826_, _08548_);
  or (_10828_, _09217_, _08549_);
  and (_10829_, _10828_, _08544_);
  and (_10830_, _10829_, _10827_);
  and (_10831_, _08542_, word_in[26]);
  or (_10176_, _10831_, _10830_);
  and (_10832_, _07979_, _06360_);
  and (_10833_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_10834_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_10835_, _10834_, _07983_);
  or (_10836_, _10835_, _10833_);
  or (_10837_, _10836_, _10832_);
  and (_10178_, _10837_, _06071_);
  not (_10838_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_10839_, _08557_, _10838_);
  and (_10840_, _09260_, _08557_);
  or (_10841_, _10840_, _10839_);
  or (_10842_, _10841_, _08552_);
  or (_10843_, _10800_, word_in[11]);
  and (_10844_, _10843_, _10842_);
  or (_10845_, _10844_, _08548_);
  or (_10846_, _09113_, _08549_);
  and (_10847_, _10846_, _08544_);
  and (_10848_, _10847_, _10845_);
  and (_10849_, _08542_, word_in[27]);
  or (_10180_, _10849_, _10848_);
  not (_10850_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_10851_, _08557_, _10850_);
  and (_10852_, _09277_, _08557_);
  or (_10853_, _10852_, _10851_);
  or (_10854_, _10853_, _08552_);
  or (_10855_, _10800_, word_in[12]);
  and (_10856_, _10855_, _10854_);
  or (_10857_, _10856_, _08548_);
  or (_10858_, _09287_, _08549_);
  and (_10859_, _10858_, _08544_);
  and (_10860_, _10859_, _10857_);
  and (_10861_, _08542_, word_in[28]);
  or (_10184_, _10861_, _10860_);
  not (_10862_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_10863_, _08557_, _10862_);
  and (_10864_, _09297_, _08557_);
  or (_10865_, _10864_, _10863_);
  or (_10866_, _10865_, _08552_);
  or (_10867_, _10800_, word_in[13]);
  and (_10868_, _10867_, _10866_);
  or (_10869_, _10868_, _08548_);
  or (_10870_, _09305_, _08549_);
  and (_10871_, _10870_, _08544_);
  and (_10872_, _10871_, _10869_);
  and (_10873_, _08542_, word_in[29]);
  or (_10187_, _10873_, _10872_);
  not (_10874_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_10875_, _08557_, _10874_);
  and (_10876_, _09315_, _08557_);
  or (_10878_, _10876_, _10875_);
  or (_10879_, _10878_, _08552_);
  nand (_10880_, _08552_, _09556_);
  and (_10881_, _10880_, _10879_);
  or (_10882_, _10881_, _08548_);
  or (_10883_, _09322_, _08549_);
  and (_10884_, _10883_, _08544_);
  and (_10885_, _10884_, _10882_);
  and (_10886_, _08542_, word_in[30]);
  or (_10190_, _10886_, _10885_);
  not (_10887_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_10888_, _09028_, _07105_);
  nand (_10889_, _10888_, _10887_);
  and (_10890_, _10889_, _08989_);
  or (_10891_, _10888_, _08799_);
  and (_10892_, _10891_, _10890_);
  nor (_10893_, _08989_, _07945_);
  or (_10894_, _10893_, _10892_);
  and (_10419_, _10894_, _06071_);
  and (_10895_, _09026_, _06815_);
  and (_10896_, _10895_, _06809_);
  not (_10897_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_10898_, _08801_, _10897_);
  nand (_10899_, _10898_, _10896_);
  or (_10900_, _10899_, _08802_);
  nand (_10902_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_10903_, _06735_, _06715_);
  and (_10904_, _06706_, _06615_);
  nor (_10905_, _10904_, _10903_);
  nor (_10906_, _10905_, _10902_);
  or (_10907_, _10902_, _06349_);
  and (_10908_, _10907_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_10910_, _10908_, _10896_);
  or (_10911_, _10910_, _10906_);
  and (_10912_, _10911_, _08985_);
  nor (_10913_, _09341_, _08985_);
  or (_10914_, _10913_, _10912_);
  and (_10915_, _10914_, _06071_);
  and (_10424_, _10915_, _10900_);
  not (_10916_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_10917_, _09028_, _06032_);
  nand (_10918_, _10917_, _10916_);
  and (_10919_, _10918_, _08989_);
  or (_10920_, _10917_, _08799_);
  and (_10921_, _10920_, _10919_);
  nor (_10922_, _08989_, _06609_);
  or (_10923_, _10922_, _10921_);
  and (_10427_, _10923_, _06071_);
  and (_10924_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_10925_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06071_);
  and (_10926_, _10925_, _07011_);
  or (_10430_, _10926_, _10924_);
  not (_10927_, _06006_);
  nor (_10928_, _06803_, _10927_);
  not (_10929_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_10930_, _06005_, _05982_);
  nor (_10931_, _10930_, _10929_);
  or (_10932_, _10931_, _10928_);
  and (_10933_, _10896_, _06071_);
  and (_10934_, _10933_, _10932_);
  not (_10935_, _10896_);
  and (_10936_, _10930_, _10927_);
  or (_10937_, _10936_, _10935_);
  and (_10938_, _10937_, _08157_);
  or (_10433_, _10938_, _10934_);
  and (_10939_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_10940_, _10939_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_10449_, _10940_, _06071_);
  and (_10941_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_10942_, _10941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_10459_, _10942_, _06071_);
  and (_10943_, _05954_, _07767_);
  and (_10944_, _06378_, _05923_);
  not (_10945_, _06815_);
  nor (_10946_, _10945_, _05967_);
  and (_10947_, _10946_, _10944_);
  and (_10948_, _10947_, _10943_);
  and (_10949_, _10948_, _06805_);
  or (_10950_, _10949_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_10951_, _07768_, _06820_);
  and (_10952_, _10951_, _09248_);
  not (_10953_, _10952_);
  and (_10954_, _10953_, _10950_);
  nand (_10955_, _10949_, _06803_);
  and (_10956_, _10955_, _10954_);
  nor (_10957_, _10953_, _06359_);
  or (_10958_, _10957_, _10956_);
  and (_10480_, _10958_, _06071_);
  and (_10959_, _10947_, _06806_);
  nand (_10960_, _10959_, _06004_);
  and (_10961_, _10960_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_10962_, _10961_, _09249_);
  or (_10963_, _07753_, _06005_);
  and (_10964_, _10963_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_10965_, _10964_, _08802_);
  and (_10966_, _10965_, _10959_);
  or (_10967_, _10966_, _10962_);
  nand (_10968_, _09341_, _09249_);
  and (_10969_, _10968_, _06071_);
  and (_10482_, _10969_, _10967_);
  and (_10970_, _09584_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and (_10971_, _09580_, _07891_);
  and (_10972_, _09005_, _10971_);
  or (_10973_, _10972_, _10970_);
  and (_10877_, _10973_, _06071_);
  and (_10974_, _07010_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_10976_, _10974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_10901_, _10976_, _06071_);
  nor (_10977_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_10978_, _10977_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_10979_, _10978_, _08110_);
  or (_10980_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_10981_, _10980_, _06071_);
  and (_10909_, _10981_, _10979_);
  not (_10982_, _08660_);
  and (_10984_, _10982_, _08619_);
  or (_10985_, _08018_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03483_, _10985_, _06071_);
  and (_10987_, _03483_, _08021_);
  and (_10975_, _10987_, _10984_);
  and (_10988_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  not (_10989_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor (_10990_, _06530_, _10989_);
  or (_10992_, _10990_, _10988_);
  and (_10983_, _10992_, _06071_);
  and (_10994_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  not (_10995_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_10997_, _06530_, _10995_);
  or (_10998_, _10997_, _10994_);
  and (_10986_, _10998_, _06071_);
  and (_11000_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11001_, _06530_, _09022_);
  or (_11002_, _11001_, _11000_);
  and (_10991_, _11002_, _06071_);
  and (_11003_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not (_11005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_11006_, _06530_, _11005_);
  or (_11007_, _11006_, _11003_);
  and (_10993_, _11007_, _06071_);
  and (_11008_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_11009_, _06530_, _05815_);
  or (_11010_, _11009_, _11008_);
  and (_10996_, _11010_, _06071_);
  and (_11011_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_11012_, _06530_, _05760_);
  or (_11013_, _11012_, _11011_);
  and (_10999_, _11013_, _06071_);
  and (_11014_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_11015_, _06530_, _05865_);
  or (_11016_, _11015_, _11014_);
  and (_11004_, _11016_, _06071_);
  and (_11017_, _06071_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_11018_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _06071_);
  and (_11019_, _11018_, _07011_);
  or (_11033_, _11019_, _11017_);
  and (_11020_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_11021_, _11020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_11034_, _11021_, _06071_);
  and (_11022_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  not (_11023_, _09037_);
  and (_11024_, _11023_, _06399_);
  and (_11025_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_11026_, _11025_, _09345_);
  or (_11027_, _11026_, _11024_);
  or (_11028_, _11027_, _11022_);
  and (_11072_, _11028_, _06071_);
  not (_11029_, _10978_);
  or (_11030_, _11029_, _07564_);
  or (_11031_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_11032_, _11031_, _06071_);
  and (_11159_, _11032_, _11030_);
  and (_11175_, _07239_, _06071_);
  not (_11035_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_11036_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_11037_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_11038_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_11039_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_11040_, _11039_, _11037_);
  and (_11041_, _11040_, _11038_);
  nor (_11042_, _11041_, _11037_);
  nor (_11043_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_11044_, _11043_, _11036_);
  not (_11045_, _11044_);
  nor (_11046_, _11045_, _11042_);
  nor (_11047_, _11046_, _11036_);
  not (_11048_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_11049_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_11050_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_11051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_11052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_11053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_11054_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_11055_, _11054_, _11053_);
  and (_11056_, _11055_, _11052_);
  and (_11057_, _11056_, _11051_);
  and (_11058_, _11057_, _11050_);
  and (_11059_, _11058_, _11049_);
  and (_11060_, _11059_, _11048_);
  and (_11061_, _11060_, _11047_);
  nor (_11062_, _11061_, _11035_);
  and (_11063_, _11061_, _11035_);
  nor (_11064_, _11063_, _11062_);
  not (_11065_, _11064_);
  and (_11066_, _11059_, _11047_);
  nor (_11067_, _11066_, _11048_);
  nor (_11068_, _11067_, _11061_);
  not (_11069_, _11068_);
  and (_11070_, _11047_, _11058_);
  nor (_11071_, _11070_, _11049_);
  or (_11073_, _11071_, _11066_);
  not (_11074_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_11075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_11076_, _11047_, _11057_);
  and (_11077_, _11076_, _11075_);
  nor (_11078_, _11077_, _11074_);
  or (_11079_, _11078_, _11070_);
  and (_11080_, _11047_, _11055_);
  and (_11081_, _11080_, _11052_);
  nor (_11082_, _11081_, _11051_);
  nor (_11083_, _11082_, _11076_);
  not (_11084_, _11083_);
  nor (_11085_, _11080_, _11052_);
  nor (_11086_, _11085_, _11081_);
  not (_11087_, _11086_);
  and (_11088_, _11047_, _11054_);
  nor (_11089_, _11088_, _11053_);
  nor (_11090_, _11089_, _11080_);
  not (_11091_, _11090_);
  nor (_11092_, _11047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11093_, _11047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_11094_, _11093_, _11092_);
  not (_11095_, _11094_);
  and (_11096_, _05769_, _05726_);
  and (_11097_, _11096_, _05880_);
  and (_11098_, _11097_, _05861_);
  not (_11099_, _11098_);
  nor (_11100_, _05810_, _05788_);
  and (_11101_, _11100_, _05848_);
  and (_11102_, _11101_, _05854_);
  nor (_11103_, _05880_, _05726_);
  and (_11104_, _05880_, _05726_);
  nor (_11105_, _11104_, _11103_);
  and (_11106_, _11105_, _11102_);
  and (_11107_, _05860_, _05788_);
  and (_11108_, _05768_, _05747_);
  and (_11109_, _11108_, _05727_);
  and (_11110_, _11109_, _05880_);
  and (_11111_, _11110_, _11107_);
  nor (_11112_, _11111_, _11106_);
  and (_11113_, _11112_, _11099_);
  nor (_11114_, _05860_, _05853_);
  nor (_11115_, _05768_, _05748_);
  and (_11116_, _11115_, _11103_);
  and (_11117_, _11108_, _05726_);
  and (_11118_, _11117_, _05880_);
  and (_11119_, _11107_, _11118_);
  nor (_11120_, _11119_, _11116_);
  nor (_11121_, _11120_, _11114_);
  and (_11122_, _11103_, _05769_);
  and (_11123_, _11101_, _11122_);
  and (_11124_, _11110_, _05847_);
  or (_11125_, _11124_, _11123_);
  nor (_11126_, _05880_, _05727_);
  and (_11127_, _11108_, _11126_);
  and (_11128_, _11107_, _11127_);
  and (_11129_, _05853_, _11122_);
  or (_11130_, _11129_, _11128_);
  or (_11131_, _11130_, _11125_);
  nor (_11132_, _11131_, _11121_);
  nand (_11133_, _11132_, _11113_);
  and (_11134_, _11102_, _11104_);
  and (_11135_, _11116_, _11101_);
  nor (_11136_, _11135_, _11134_);
  and (_11137_, _11126_, _05769_);
  and (_11138_, _11115_, _05726_);
  and (_11139_, _11138_, _05880_);
  nor (_11140_, _11139_, _11137_);
  nor (_11141_, _11140_, _05857_);
  and (_11142_, _05880_, _05727_);
  and (_11143_, _11142_, _05769_);
  or (_11144_, _11139_, _11143_);
  and (_11145_, _11144_, _05861_);
  nor (_11146_, _11145_, _11141_);
  and (_11147_, _05861_, _05855_);
  and (_11148_, _11107_, _05854_);
  nor (_11149_, _11148_, _11147_);
  and (_11150_, _11149_, _11146_);
  and (_11151_, _11115_, _11126_);
  nor (_11152_, _05860_, _05849_);
  not (_11153_, _11152_);
  and (_11154_, _11153_, _11151_);
  not (_11155_, _05853_);
  nor (_11156_, _11110_, _11139_);
  nor (_11157_, _11156_, _11155_);
  nor (_11158_, _11157_, _11154_);
  not (_11160_, _11107_);
  and (_11161_, _11108_, _11103_);
  nor (_11162_, _11161_, _11143_);
  nor (_11163_, _11162_, _11160_);
  nor (_11164_, _11161_, _11097_);
  nor (_11165_, _11164_, _11155_);
  nor (_11166_, _11165_, _11163_);
  and (_11167_, _11166_, _11158_);
  and (_11168_, _11167_, _11150_);
  nand (_11169_, _11168_, _11136_);
  and (_11170_, _11097_, _11107_);
  and (_11171_, _11115_, _11142_);
  and (_11172_, _11171_, _05850_);
  nor (_11173_, _11172_, _11170_);
  nor (_11174_, _11139_, _11122_);
  nor (_11176_, _11174_, _11160_);
  and (_11177_, _05854_, _05727_);
  and (_11178_, _11177_, _05853_);
  nor (_11179_, _11178_, _11176_);
  nand (_11180_, _11179_, _11173_);
  not (_11182_, _11171_);
  nor (_11183_, _11114_, _11182_);
  and (_11185_, _11116_, _05850_);
  and (_11186_, _11101_, _11143_);
  nor (_11187_, _11186_, _11185_);
  not (_11189_, _11187_);
  or (_11190_, _11189_, _11183_);
  or (_11191_, _11190_, _11180_);
  and (_11192_, _05880_, _05857_);
  and (_11193_, _05829_, _05810_);
  and (_11194_, _11193_, _11192_);
  or (_11195_, _11194_, _11101_);
  and (_11196_, _11195_, _11138_);
  and (_11197_, _11194_, _11096_);
  nand (_11198_, _05847_, _05769_);
  nor (_11199_, _11198_, _11105_);
  or (_11200_, _11199_, _11197_);
  and (_11201_, _05858_, _05788_);
  and (_11202_, _11201_, _05848_);
  and (_11203_, _05882_, _05857_);
  and (_11204_, _11203_, _11193_);
  or (_11206_, _11204_, _11202_);
  or (_11207_, _11206_, _11200_);
  or (_11208_, _11207_, _11196_);
  and (_11209_, _05853_, _05769_);
  and (_11210_, _11209_, _11105_);
  or (_11211_, _11109_, _11171_);
  or (_11212_, _11211_, _11097_);
  or (_11213_, _11212_, _11137_);
  and (_11214_, _11213_, _11101_);
  or (_11215_, _11214_, _11210_);
  or (_11216_, _11215_, _11208_);
  or (_11217_, _11216_, _11191_);
  or (_11218_, _11217_, _11169_);
  nor (_11219_, _11218_, _11133_);
  nor (_11221_, _11040_, _11038_);
  nor (_11222_, _11221_, _11041_);
  not (_11224_, _11222_);
  nor (_11225_, _11224_, _11219_);
  and (_11226_, _11151_, _05850_);
  nor (_11227_, _11226_, _11134_);
  and (_11228_, _11227_, _11187_);
  and (_11229_, _11228_, _11113_);
  and (_11230_, _11097_, _05847_);
  nor (_11231_, _11230_, _11197_);
  and (_11232_, _11231_, _11173_);
  and (_11233_, _11232_, _11179_);
  and (_11234_, _11233_, _11229_);
  not (_11235_, _11234_);
  nor (_11236_, _11235_, _11219_);
  not (_11237_, _11236_);
  nor (_11238_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_11239_, _11238_, _11038_);
  and (_11240_, _11239_, _11237_);
  and (_11241_, _11224_, _11219_);
  nor (_11242_, _11241_, _11225_);
  and (_11243_, _11242_, _11240_);
  nor (_11244_, _11243_, _11225_);
  not (_11245_, _11244_);
  and (_11246_, _11045_, _11042_);
  nor (_11247_, _11246_, _11046_);
  and (_11248_, _11247_, _11245_);
  and (_11249_, _11248_, _11095_);
  and (_11250_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_11251_, _11250_, _11054_);
  nand (_11252_, _11251_, _11092_);
  or (_11253_, _11251_, _11092_);
  and (_11254_, _11253_, _11252_);
  and (_11255_, _11254_, _11249_);
  and (_11256_, _11255_, _11091_);
  and (_11257_, _11256_, _11087_);
  and (_11258_, _11257_, _11084_);
  nor (_11259_, _11076_, _11075_);
  or (_11260_, _11259_, _11077_);
  and (_11261_, _11260_, _11258_);
  and (_11262_, _11261_, _11079_);
  and (_11263_, _11262_, _11073_);
  and (_11264_, _11263_, _11069_);
  and (_11265_, _11264_, _11065_);
  nor (_11266_, _11264_, _11065_);
  nor (_11267_, _11266_, _11265_);
  or (_11268_, _11267_, _09711_);
  or (_11269_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_11270_, rst, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_11271_, _11270_, _11269_);
  and (_11272_, _11271_, _11268_);
  and (_11273_, _06071_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_11274_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_11181_, _11274_, _11272_);
  and (_11275_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not (_11276_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_11277_, _06530_, _11276_);
  or (_11278_, _11277_, _11275_);
  and (_11184_, _11278_, _06071_);
  and (_11279_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11280_, _06530_, _09701_);
  or (_11281_, _11280_, _11279_);
  and (_11188_, _11281_, _06071_);
  and (_11282_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_11283_, _06530_, _05833_);
  or (_11284_, _11283_, _11282_);
  and (_11205_, _11284_, _06071_);
  not (_11286_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_11287_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_11288_, _11063_, _11287_);
  nor (_11289_, _11288_, _11286_);
  and (_11290_, _11288_, _11286_);
  nor (_11292_, _11290_, _11289_);
  not (_11293_, _11292_);
  nor (_11294_, _11063_, _11287_);
  or (_11295_, _11294_, _11288_);
  and (_11296_, _11295_, _11265_);
  and (_11297_, _11296_, _11293_);
  nor (_11298_, _11296_, _11293_);
  nor (_11299_, _11298_, _11297_);
  or (_11300_, _11299_, _09711_);
  or (_11301_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_11302_, _11301_, _11270_);
  and (_11304_, _11302_, _11300_);
  and (_11305_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_11220_, _11305_, _11304_);
  nor (_11307_, _11295_, _11265_);
  nor (_11308_, _11307_, _11296_);
  or (_11309_, _11308_, _09711_);
  or (_11310_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_11311_, _11310_, _11270_);
  and (_11312_, _11311_, _11309_);
  and (_11313_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_11223_, _11313_, _11312_);
  or (_11314_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_11315_, _06530_, _05737_);
  and (_11316_, _11315_, _06071_);
  and (_11285_, _11316_, _11314_);
  nor (_11317_, _11263_, _11069_);
  nor (_11318_, _11317_, _11264_);
  or (_11319_, _11318_, _09711_);
  or (_11320_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_11321_, _11320_, _11270_);
  and (_11322_, _11321_, _11319_);
  and (_11323_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_11291_, _11323_, _11322_);
  and (_11324_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_11325_, _06530_, _06958_);
  or (_11326_, _11325_, _11324_);
  and (_11303_, _11326_, _06071_);
  and (_11327_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_11328_, _06530_, _05862_);
  or (_11329_, _11328_, _11327_);
  and (_11306_, _11329_, _06071_);
  and (_11330_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_11331_, _06530_, _05693_);
  or (_11332_, _11331_, _11330_);
  and (_11339_, _11332_, _06071_);
  nor (_11333_, _06527_, _06231_);
  or (_11334_, _05811_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor (_11335_, _05718_, _10690_);
  nor (_11336_, _05696_, _10989_);
  or (_11337_, _11336_, _11335_);
  and (_11338_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11340_, _05711_, _05817_);
  nor (_11341_, _05705_, _05815_);
  or (_11342_, _11341_, _11340_);
  or (_11343_, _11342_, _11338_);
  or (_11344_, _11343_, _11337_);
  and (_11345_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_11346_, _11345_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_11347_, _11346_, _11344_);
  and (_11348_, _11347_, _06527_);
  and (_11349_, _11348_, _11334_);
  nor (_11350_, _11349_, _11333_);
  nor (_11373_, _11350_, rst);
  nor (_11351_, _06527_, _06224_);
  nor (_11352_, _05705_, _05789_);
  nor (_11353_, _05711_, _05791_);
  nor (_11354_, _11353_, _11352_);
  and (_11355_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_11356_, _05700_, _05793_);
  nor (_11357_, _11356_, _11355_);
  and (_11358_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_11359_, _05718_);
  and (_11360_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_11361_, _11360_, _11358_);
  and (_11362_, _11361_, _11357_);
  and (_11363_, _11362_, _11354_);
  nor (_11364_, _11363_, _09711_);
  nor (_11365_, _11364_, _11351_);
  nor (_11389_, _11365_, rst);
  nor (_11366_, _11236_, _05709_);
  nor (_11367_, _11219_, _05698_);
  and (_11368_, _11219_, _05698_);
  nor (_11369_, _11368_, _11367_);
  and (_11370_, _11369_, _11366_);
  nor (_11371_, _11369_, _11366_);
  nor (_11372_, _11371_, _11370_);
  or (_11374_, _11372_, _06528_);
  or (_11375_, _06527_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_11376_, _11375_, _11270_);
  and (_11393_, _11376_, _11374_);
  and (_11377_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_11378_, _11262_, _11073_);
  nor (_11379_, _11378_, _11263_);
  or (_11380_, _11379_, _09711_);
  or (_11381_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_11382_, _11381_, _11270_);
  and (_11383_, _11382_, _11380_);
  or (_11402_, _11383_, _11377_);
  and (_11384_, \oc8051_top_1.oc8051_decoder1.state [1], _05686_);
  and (_11385_, _11384_, _05685_);
  and (_11386_, _08740_, _08737_);
  nor (_11387_, _08746_, _11386_);
  and (_11388_, _11387_, _08736_);
  and (_11390_, _08714_, _08712_);
  and (_11391_, _08732_, _11390_);
  and (_11392_, _08710_, _08707_);
  and (_11394_, _08715_, _11392_);
  and (_11395_, _11394_, _08725_);
  and (_11396_, _11395_, _08732_);
  or (_11397_, _11396_, _11391_);
  nand (_11398_, _11397_, _11388_);
  not (_11399_, _08736_);
  and (_11400_, _08758_, _11399_);
  and (_11401_, _11400_, _08732_);
  and (_11403_, _11401_, _08728_);
  and (_11404_, _11387_, _11399_);
  and (_11405_, _11404_, _08728_);
  nor (_11406_, _11405_, _11403_);
  and (_11407_, _08746_, _11386_);
  and (_11408_, _11407_, _08736_);
  and (_11410_, _11408_, _08732_);
  and (_11411_, _08726_, _08753_);
  and (_11412_, _11411_, _11394_);
  and (_11413_, _11412_, _11410_);
  and (_11414_, _11388_, _08732_);
  and (_11415_, _11394_, _08726_);
  and (_11416_, _11415_, _11414_);
  nor (_11417_, _11416_, _11413_);
  and (_11418_, _11417_, _11406_);
  nand (_11419_, _11418_, _11398_);
  nand (_11420_, _11419_, _11385_);
  or (_11421_, _06526_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11422_, _08756_, _08721_);
  and (_11423_, _11422_, _11400_);
  and (_11424_, _11423_, _11421_);
  not (_11425_, _11424_);
  and (_11426_, _11384_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11427_, _11422_, _11404_);
  nand (_11428_, _11427_, _11426_);
  nand (_11429_, _11421_, _11405_);
  and (_11430_, _11429_, _11428_);
  and (_11431_, _11430_, _11425_);
  nand (_11433_, _11431_, _11420_);
  nor (_11434_, _06527_, _06080_);
  and (_11435_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11436_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_11438_, _05700_, _05754_);
  nor (_11439_, _11438_, _11436_);
  nor (_11441_, _05705_, _05749_);
  and (_11442_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_11444_, _11442_, _11441_);
  nor (_11445_, _05718_, _10995_);
  nor (_11446_, _05711_, _05760_);
  nor (_11447_, _11446_, _11445_);
  and (_11448_, _11447_, _11444_);
  and (_11449_, _11448_, _11439_);
  nor (_11450_, _11449_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11451_, _11450_, _11435_);
  nor (_11452_, _11451_, _06528_);
  nor (_11453_, _11452_, _11434_);
  and (_11454_, _11453_, _11433_);
  and (_11455_, _11431_, _11420_);
  nor (_11456_, _06527_, _06075_);
  nor (_11457_, _05705_, _05760_);
  nor (_11458_, _05711_, _05754_);
  nor (_11459_, _11458_, _11457_);
  nor (_11460_, _05696_, _10995_);
  nor (_11461_, _05700_, _05756_);
  nor (_11462_, _11461_, _11460_);
  and (_11463_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_11464_, _05718_, _05749_);
  nor (_11465_, _11464_, _11463_);
  and (_11466_, _11465_, _11462_);
  and (_11467_, _11466_, _11459_);
  nor (_11468_, _11467_, _09711_);
  nor (_11469_, _11468_, _11456_);
  and (_11470_, _11469_, _11455_);
  nor (_11471_, _11470_, _11454_);
  not (_11472_, _11471_);
  and (_11473_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_11474_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_11475_, _11474_);
  nor (_11476_, _06527_, _06258_);
  and (_11477_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11478_, _05696_, _06850_);
  and (_11479_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_11480_, _11479_, _11478_);
  nor (_11481_, _05705_, _05737_);
  and (_11482_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_11483_, _11482_, _11481_);
  and (_11484_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_11485_, _05711_, _05739_);
  nor (_11486_, _11485_, _11484_);
  and (_11487_, _11486_, _11483_);
  and (_11488_, _11487_, _11480_);
  nor (_11490_, _11488_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11491_, _11490_, _11477_);
  nor (_11492_, _11491_, _06528_);
  nor (_11493_, _11492_, _11476_);
  and (_11495_, _11493_, _11433_);
  nor (_11496_, _06527_, _06256_);
  nor (_11497_, _05705_, _05739_);
  and (_11498_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_11500_, _11498_, _11497_);
  and (_11501_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_11503_, _05700_, _05732_);
  nor (_11504_, _11503_, _11501_);
  and (_11505_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_11506_, _05718_, _05737_);
  nor (_11507_, _11506_, _11505_);
  and (_11508_, _11507_, _11504_);
  and (_11509_, _11508_, _11500_);
  nor (_11510_, _11509_, _09711_);
  nor (_11511_, _11510_, _11496_);
  and (_11512_, _11511_, _11455_);
  nor (_11513_, _11512_, _11495_);
  nand (_11514_, _11513_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_11515_, _11513_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_11516_, _11515_, _11514_);
  nor (_11517_, _06527_, _06277_);
  and (_11518_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11519_, _05696_, _06532_);
  and (_11520_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_11521_, _11520_, _11519_);
  nor (_11522_, _05705_, _05693_);
  and (_11523_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11524_, _11523_, _11522_);
  and (_11525_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_11526_, _05711_, _05716_);
  nor (_11527_, _11526_, _11525_);
  and (_11528_, _11527_, _11524_);
  and (_11529_, _11528_, _11521_);
  nor (_11530_, _11529_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11531_, _11530_, _11518_);
  nor (_11532_, _11531_, _06528_);
  nor (_11533_, _11532_, _11517_);
  and (_11534_, _11533_, _11433_);
  nor (_11535_, _06527_, _06279_);
  nor (_11536_, _05705_, _05716_);
  and (_11537_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_11538_, _11537_, _11536_);
  and (_11539_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_11540_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_11541_, _11540_, _11539_);
  nor (_11542_, _05718_, _05693_);
  nor (_11543_, _05700_, _05708_);
  nor (_11545_, _11543_, _11542_);
  and (_11546_, _11545_, _11541_);
  and (_11547_, _11546_, _11538_);
  nor (_11548_, _11547_, _09711_);
  nor (_11549_, _11548_, _11535_);
  and (_11550_, _11549_, _11455_);
  nor (_11551_, _11550_, _11534_);
  nor (_11552_, _11551_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_11553_, _11551_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_11554_, _06527_, _06148_);
  or (_11555_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05811_);
  nor (_11556_, _05718_, _09701_);
  nor (_11557_, _05696_, _06958_);
  or (_11558_, _11557_, _11556_);
  and (_11559_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11560_, _05705_, _05862_);
  nor (_11561_, _05711_, _05865_);
  or (_11562_, _11561_, _11560_);
  or (_11563_, _11562_, _11559_);
  or (_11564_, _11563_, _11558_);
  and (_11565_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_11566_, _11565_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_11567_, _11566_, _11564_);
  and (_11568_, _11567_, _06527_);
  and (_11569_, _11568_, _11555_);
  nor (_11570_, _11569_, _11554_);
  and (_11571_, _11570_, _11433_);
  and (_11572_, _11455_, _09713_);
  nor (_11573_, _11572_, _11571_);
  nand (_11574_, _11573_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_11575_, _06527_, _06167_);
  and (_11576_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11577_, _05696_, _11276_);
  and (_11578_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_11579_, _11578_, _11577_);
  nor (_11580_, _05705_, _05833_);
  and (_11581_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11582_, _11581_, _11580_);
  nor (_11583_, _05718_, _09022_);
  nor (_11584_, _05711_, _05835_);
  nor (_11585_, _11584_, _11583_);
  and (_11586_, _11585_, _11582_);
  and (_11587_, _11586_, _11579_);
  nor (_11588_, _11587_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11589_, _11588_, _11576_);
  nor (_11590_, _11589_, _06528_);
  nor (_11591_, _11590_, _11575_);
  and (_11592_, _11591_, _11433_);
  nor (_11593_, _06527_, _06169_);
  nor (_11594_, _05705_, _05835_);
  and (_11595_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_11596_, _11595_, _11594_);
  nor (_11597_, _05696_, _09022_);
  and (_11598_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_11600_, _11598_, _11597_);
  nor (_11601_, _05718_, _05833_);
  and (_11602_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11603_, _11602_, _11601_);
  and (_11604_, _11603_, _11600_);
  and (_11605_, _11604_, _11596_);
  nor (_11606_, _11605_, _09711_);
  nor (_11607_, _11606_, _11593_);
  and (_11608_, _11607_, _11455_);
  nor (_11609_, _11608_, _11592_);
  nor (_11610_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_11611_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_11612_, _11350_);
  or (_11613_, _11455_, _11612_);
  nor (_11614_, _06527_, _06233_);
  nor (_11615_, _05705_, _05817_);
  and (_11616_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11617_, _11616_, _11615_);
  nor (_11618_, _05696_, _10690_);
  and (_11619_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11620_, _11619_, _11618_);
  and (_11621_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_11622_, _05718_, _05815_);
  nor (_11623_, _11622_, _11621_);
  and (_11624_, _11623_, _11620_);
  and (_11625_, _11624_, _11617_);
  nor (_11626_, _11625_, _09711_);
  nor (_11627_, _11626_, _11614_);
  not (_11628_, _11627_);
  or (_11629_, _11628_, _11433_);
  nand (_11630_, _11629_, _11613_);
  or (_11631_, _11630_, _06241_);
  nor (_11632_, _06527_, _06214_);
  and (_11633_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11634_, _05801_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nor (_11635_, _05700_, _05791_);
  nor (_11636_, _11635_, _11634_);
  and (_11637_, _05706_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_11638_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_11639_, _11638_, _11637_);
  and (_11640_, _11359_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_11641_, _05711_, _05789_);
  nor (_11642_, _11641_, _11640_);
  and (_11643_, _11642_, _11639_);
  and (_11644_, _11643_, _11636_);
  nor (_11645_, _11644_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11646_, _11645_, _11633_);
  nor (_11647_, _11646_, _06528_);
  nor (_11648_, _11647_, _11632_);
  not (_11649_, _11648_);
  or (_11650_, _11649_, _11455_);
  not (_11651_, _11365_);
  or (_11652_, _11433_, _11651_);
  and (_11653_, _11652_, _11650_);
  nand (_11654_, _11653_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_11655_, _06527_, _06190_);
  and (_11656_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11657_, _05696_, _06962_);
  and (_11658_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_11659_, _11658_, _11657_);
  nor (_11660_, _05705_, _05782_);
  and (_11661_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_11662_, _11661_, _11660_);
  nor (_11663_, _05718_, _11005_);
  nor (_11664_, _05711_, _05773_);
  nor (_11665_, _11664_, _11663_);
  and (_11666_, _11665_, _11662_);
  and (_11667_, _11666_, _11659_);
  nor (_11668_, _11667_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11669_, _11668_, _11656_);
  nor (_11670_, _11669_, _06528_);
  nor (_11671_, _11670_, _11655_);
  not (_11672_, _11671_);
  or (_11673_, _11672_, _11455_);
  nor (_11674_, _06527_, _06188_);
  nor (_11675_, _05705_, _05773_);
  and (_11676_, _05778_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_11678_, _11676_, _11675_);
  nor (_11679_, _05696_, _11005_);
  and (_11680_, _05701_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_11681_, _11680_, _11679_);
  and (_11682_, _05714_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_11683_, _05718_, _05782_);
  nor (_11684_, _11683_, _11682_);
  and (_11685_, _11684_, _11681_);
  and (_11686_, _11685_, _11678_);
  nor (_11687_, _11686_, _09711_);
  nor (_11688_, _11687_, _11674_);
  not (_11689_, _11688_);
  or (_11690_, _11689_, _11433_);
  and (_11691_, _11690_, _11673_);
  and (_11693_, _11691_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_11694_, _11653_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_11695_, _11694_, _11654_);
  and (_11696_, _11695_, _11693_);
  not (_11697_, _11696_);
  nand (_11698_, _11697_, _11654_);
  nand (_11699_, _11630_, _06241_);
  and (_11700_, _11699_, _11631_);
  and (_11701_, _11700_, _11698_);
  not (_11702_, _11701_);
  nand (_11703_, _11702_, _11631_);
  nor (_11704_, _11703_, _11611_);
  nor (_11705_, _11704_, _11610_);
  or (_11706_, _11573_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_11707_, _11706_, _11574_);
  nand (_11708_, _11707_, _11705_);
  nand (_11709_, _11708_, _11574_);
  nor (_11710_, _11709_, _11553_);
  nor (_11711_, _11710_, _11552_);
  nand (_11713_, _11711_, _11516_);
  nand (_11714_, _11713_, _11514_);
  and (_11715_, _11714_, _11475_);
  or (_11716_, _11715_, _11473_);
  or (_11717_, _11716_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_11718_, _11717_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_11719_, _11718_, _06243_);
  or (_11721_, _11719_, _11472_);
  and (_11722_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_11723_, _11722_, _11716_);
  and (_11724_, _11723_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_11725_, _11724_, _11472_);
  and (_11726_, _11725_, _11721_);
  nand (_11727_, _11726_, _06172_);
  or (_11728_, _11726_, _06172_);
  and (_11729_, _11429_, _11420_);
  not (_11730_, _11385_);
  nor (_11731_, _08741_, _08736_);
  and (_11732_, _11731_, _08728_);
  and (_11733_, _08760_, _08764_);
  and (_11734_, _11733_, _08728_);
  or (_11735_, _11734_, _11732_);
  and (_11736_, _08748_, _11399_);
  and (_11737_, _11736_, _08732_);
  and (_11738_, _11737_, _08757_);
  and (_11739_, _11410_, _11390_);
  or (_11740_, _11739_, _11738_);
  nor (_11741_, _11740_, _11735_);
  or (_11742_, _11741_, _11730_);
  and (_11743_, _11742_, _11729_);
  not (_11744_, _11421_);
  and (_11745_, _11411_, _08717_);
  nor (_11746_, _11745_, _11423_);
  nor (_11747_, _11746_, _11744_);
  and (_11748_, _11738_, _11385_);
  nor (_11749_, _11748_, _11747_);
  nor (_11750_, _11749_, _11433_);
  nor (_11751_, _11750_, _11743_);
  and (_11752_, _11751_, _11728_);
  and (_11753_, _11752_, _11727_);
  not (_11754_, _07108_);
  or (_11755_, _07324_, _07297_);
  and (_11756_, _07323_, _07320_);
  nor (_11757_, _11756_, _11755_);
  and (_11758_, _11756_, _11755_);
  nor (_11759_, _11758_, _11757_);
  nor (_11760_, _11759_, _07531_);
  not (_11761_, _07296_);
  and (_11762_, _07531_, _11761_);
  or (_11763_, _11762_, _11760_);
  or (_11764_, _11763_, _11754_);
  not (_11765_, _07344_);
  or (_11766_, _07751_, _11765_);
  and (_11768_, _06731_, _06725_);
  or (_11769_, _11768_, _06716_);
  nor (_11770_, _11769_, _06732_);
  not (_11771_, _11770_);
  and (_11772_, _06699_, _06685_);
  nor (_11773_, _11772_, _06700_);
  nor (_11774_, _11773_, _06616_);
  not (_11775_, _11774_);
  or (_11776_, _07411_, _06166_);
  and (_11777_, _06352_, _06251_);
  and (_11778_, _06349_, _06305_);
  nor (_11779_, _11778_, _11777_);
  and (_11780_, _11779_, _11776_);
  and (_11781_, _11780_, _07940_);
  nor (_11782_, _06252_, _10897_);
  or (_11783_, _11782_, _06305_);
  nand (_11784_, _11783_, _07696_);
  and (_11785_, _11784_, _07937_);
  and (_11786_, _11785_, _07934_);
  and (_11787_, _11786_, _11781_);
  and (_11788_, _11787_, _11775_);
  and (_11789_, _11788_, _11771_);
  and (_11790_, _11789_, _11766_);
  and (_11791_, _11790_, _11764_);
  nor (_11792_, _11791_, _11428_);
  and (_11793_, _11732_, _11385_);
  not (_11794_, _11793_);
  and (_11795_, \oc8051_top_1.oc8051_decoder1.state [0], _05686_);
  not (_11796_, _11406_);
  and (_11797_, _11793_, _08746_);
  nor (_11798_, _11797_, _11796_);
  nor (_11799_, _11798_, _11795_);
  and (_11800_, _11799_, _11794_);
  and (_11801_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11802_, _11388_, _08764_);
  and (_11803_, _11802_, _08757_);
  nor (_11804_, _11803_, _11738_);
  and (_11805_, _08760_, _08732_);
  and (_11806_, _11805_, _08757_);
  not (_11807_, _11806_);
  and (_11808_, _11807_, _11804_);
  and (_11810_, _11394_, _08727_);
  and (_11811_, _11802_, _11810_);
  and (_11812_, _11733_, _11810_);
  nor (_11813_, _11812_, _11811_);
  and (_11814_, _11813_, _11808_);
  nor (_11815_, _11814_, _11744_);
  not (_11816_, _11815_);
  and (_11817_, _11811_, _05686_);
  and (_11818_, _11812_, _05686_);
  nor (_11819_, _11818_, _11817_);
  nor (_11821_, _11819_, _06526_);
  nor (_11822_, _11821_, _11793_);
  and (_11823_, _11822_, _11816_);
  nor (_11824_, _11823_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11825_, _11824_, _11801_);
  and (_11826_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11827_, _11428_);
  and (_11828_, _11737_, _11422_);
  not (_11829_, _11828_);
  and (_11830_, _11731_, _08746_);
  and (_11831_, _11830_, _08764_);
  and (_11833_, _11831_, _08757_);
  and (_11834_, _11831_, _11422_);
  nor (_11835_, _11834_, _11833_);
  and (_11836_, _11835_, _11829_);
  and (_11837_, _11414_, _08728_);
  not (_11838_, _11837_);
  and (_11839_, _11422_, _11414_);
  and (_11840_, _11408_, _08764_);
  and (_11841_, _11840_, _11422_);
  nor (_11842_, _11841_, _11839_);
  nand (_11843_, _11842_, _11838_);
  and (_11844_, _11831_, _11412_);
  and (_11845_, _11802_, _08728_);
  nor (_11846_, _11845_, _11844_);
  and (_11847_, _11412_, _11401_);
  nor (_11848_, _11847_, _11413_);
  nand (_11849_, _11848_, _11846_);
  nor (_11850_, _11849_, _11843_);
  and (_11851_, _11850_, _11836_);
  and (_11852_, _11736_, _08764_);
  and (_11853_, _11852_, _08757_);
  and (_11854_, _11852_, _11422_);
  nor (_11855_, _11854_, _11853_);
  and (_11856_, _11414_, _11412_);
  and (_11857_, _11733_, _11412_);
  nor (_11858_, _11857_, _11856_);
  and (_11859_, _11840_, _11412_);
  and (_11860_, _11408_, _08728_);
  nor (_11861_, _11860_, _11859_);
  and (_11862_, _11861_, _11858_);
  and (_11863_, _11862_, _11855_);
  and (_11864_, _11852_, _11412_);
  and (_11865_, _11422_, _11410_);
  nor (_11866_, _11865_, _11864_);
  and (_11867_, _11830_, _08732_);
  and (_11868_, _11867_, _08756_);
  and (_11869_, _11733_, _11422_);
  nor (_11870_, _11869_, _11868_);
  and (_11872_, _11870_, _11866_);
  and (_11873_, _11872_, _11863_);
  and (_11874_, _11395_, _08764_);
  and (_11875_, _11874_, _11388_);
  and (_11876_, _11802_, _11422_);
  nor (_11877_, _11876_, _11875_);
  nor (_11878_, _11867_, _11404_);
  not (_11879_, _11878_);
  and (_11880_, _11879_, _11412_);
  and (_11881_, _11805_, _11422_);
  nor (_11882_, _11881_, _11880_);
  and (_11883_, _11882_, _11877_);
  and (_11884_, _11400_, _08764_);
  and (_11885_, _11884_, _11412_);
  and (_11887_, _11412_, _08765_);
  nor (_11888_, _11887_, _11885_);
  nor (_11889_, _08732_, _08715_);
  and (_11890_, _11889_, _11388_);
  and (_11891_, _11805_, _11412_);
  nor (_11893_, _11891_, _11890_);
  and (_11894_, _11893_, _11888_);
  not (_11895_, _11427_);
  and (_11896_, _11895_, _11406_);
  and (_11897_, _11896_, _11894_);
  and (_11899_, _11897_, _11883_);
  and (_11900_, _11899_, _11873_);
  and (_11901_, _11900_, _11851_);
  nor (_11902_, _11901_, _11744_);
  nor (_11903_, _11902_, _11827_);
  and (_11904_, _11903_, _11794_);
  nor (_11905_, _11904_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11906_, _11905_, _11826_);
  and (_11907_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11908_, _11408_, _11395_);
  and (_11909_, _11805_, _11395_);
  nor (_11910_, _11909_, _11908_);
  or (_11911_, _11414_, _11400_);
  and (_11912_, _11911_, _11395_);
  nor (_11913_, _11912_, _11427_);
  and (_11914_, _11913_, _11910_);
  or (_11915_, _11879_, _11831_);
  and (_11916_, _11915_, _11395_);
  and (_11917_, _11733_, _11395_);
  and (_11918_, _11852_, _11395_);
  or (_11919_, _11918_, _11917_);
  and (_11920_, _11410_, _08728_);
  and (_11921_, _11395_, _08765_);
  or (_11922_, _11921_, _11920_);
  or (_11923_, _11922_, _11919_);
  nor (_11924_, _11923_, _11916_);
  and (_11925_, _11924_, _11914_);
  and (_11926_, _11925_, _11808_);
  nor (_11927_, _11926_, _11744_);
  nor (_11928_, _11799_, _11794_);
  nor (_11929_, _11928_, _11827_);
  not (_11930_, _11929_);
  nor (_11931_, _11930_, _11927_);
  nor (_11932_, _11931_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11933_, _11932_, _11907_);
  nor (_11934_, _11933_, _11906_);
  and (_11935_, _11934_, _11825_);
  and (_11936_, _06363_, _06012_);
  and (_11937_, _11936_, _06840_);
  not (_11938_, _11937_);
  nor (_11939_, _11938_, _07945_);
  and (_11940_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_11942_, _11940_, _11939_);
  and (_11943_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_11944_, _11938_, _06434_);
  nor (_11945_, _11944_, _11943_);
  and (_11946_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_11947_, _11938_, _09037_);
  nor (_11948_, _11947_, _11946_);
  nor (_11949_, _11937_, _05997_);
  and (_11950_, _11937_, _07978_);
  nor (_11951_, _11950_, _11949_);
  and (_11952_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_11953_, _11952_, _11948_);
  and (_11954_, _11953_, _11945_);
  and (_11955_, _11954_, _11942_);
  nor (_11956_, _11954_, _11942_);
  or (_11957_, _11956_, _11955_);
  and (_11958_, _11957_, _05899_);
  or (_11959_, _11958_, _06017_);
  and (_11960_, _11959_, _11938_);
  or (_11961_, _11960_, _11939_);
  and (_11962_, _11961_, _11935_);
  not (_11963_, _11962_);
  and (_11964_, _08985_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_11965_, _11964_, _10893_);
  not (_11966_, _11965_);
  and (_11967_, _11933_, _11825_);
  and (_11968_, _11967_, _11906_);
  and (_11969_, _11968_, _11966_);
  not (_11970_, _11933_);
  and (_11971_, _11970_, _11906_);
  and (_11972_, _11971_, _11825_);
  and (_11973_, _05923_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_11974_, _08991_, _06364_);
  nor (_11975_, _11974_, _11973_);
  and (_11976_, _11965_, _06378_);
  not (_11977_, _11976_);
  nor (_11978_, _11965_, _06378_);
  not (_11979_, _11978_);
  and (_11980_, _08721_, _06030_);
  and (_11981_, _08753_, _06004_);
  or (_11982_, _11981_, _11980_);
  nor (_11983_, _11982_, _09348_);
  and (_11984_, _11983_, _11979_);
  and (_11985_, _11984_, _11977_);
  and (_11986_, _11985_, _11975_);
  not (_11987_, _08991_);
  nor (_11989_, _11965_, _08721_);
  and (_11990_, _11989_, _11987_);
  and (_11991_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_11992_, _11965_, _08721_);
  and (_11993_, _11992_, _08991_);
  and (_11994_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_11995_, _11994_, _11991_);
  nor (_11996_, _11965_, _08753_);
  and (_11997_, _11996_, _08991_);
  and (_11998_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_11999_, _11965_, _08753_);
  and (_12000_, _11999_, _11987_);
  and (_12001_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_12002_, _12001_, _11998_);
  and (_12003_, _12002_, _11995_);
  and (_12004_, _11992_, _11987_);
  and (_12005_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_12006_, _11999_, _08991_);
  and (_12007_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_12008_, _12007_, _12005_);
  and (_12009_, _11996_, _11987_);
  and (_12010_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_12011_, _11989_, _08991_);
  and (_12013_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_12014_, _12013_, _12010_);
  and (_12015_, _12014_, _12008_);
  and (_12016_, _12015_, _12003_);
  nor (_12017_, _12016_, _11986_);
  not (_12019_, _07945_);
  and (_12020_, _11986_, _12019_);
  nor (_12021_, _12020_, _12017_);
  not (_12022_, _12021_);
  and (_12023_, _12022_, _11972_);
  not (_12024_, _11607_);
  nor (_12025_, _11970_, _11906_);
  and (_12026_, _12025_, _11825_);
  and (_12027_, _12026_, _12024_);
  or (_12028_, _12027_, _12023_);
  nor (_12029_, _12028_, _11969_);
  and (_12030_, _12029_, _11963_);
  nor (_12031_, _12030_, _06378_);
  and (_12032_, _12030_, _06378_);
  nor (_12033_, _12032_, _12031_);
  and (_12034_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_12035_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_12036_, _12035_, _12034_);
  and (_12037_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_12038_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_12039_, _12038_, _12037_);
  and (_12040_, _12039_, _12036_);
  and (_12041_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_12042_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_12043_, _12042_, _12041_);
  and (_12044_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_12045_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_12046_, _12045_, _12044_);
  and (_12047_, _12046_, _12043_);
  and (_12049_, _12047_, _12040_);
  nor (_12050_, _12049_, _11986_);
  and (_12051_, _11986_, _06360_);
  nor (_12052_, _12051_, _12050_);
  not (_12053_, _12052_);
  and (_12054_, _12053_, _11972_);
  not (_12055_, _12054_);
  nor (_12056_, _11938_, _06359_);
  nor (_12057_, _11938_, _06993_);
  and (_12058_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_12059_, _12058_, _12057_);
  and (_12060_, _12059_, _11955_);
  nor (_12061_, _11938_, _06609_);
  and (_12062_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_12063_, _12062_, _12061_);
  and (_12064_, _12063_, _12060_);
  nor (_12065_, _11938_, _09341_);
  and (_12066_, _11938_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_12067_, _12066_, _12065_);
  and (_12068_, _12067_, _12064_);
  nor (_12069_, _11937_, _05955_);
  nor (_12070_, _12069_, _12068_);
  and (_12071_, _12069_, _12068_);
  or (_12072_, _12071_, _12070_);
  nor (_12073_, _12072_, _05898_);
  or (_12074_, _12073_, _05959_);
  and (_12075_, _12074_, _11938_);
  or (_12076_, _12075_, _12056_);
  and (_12077_, _12076_, _11934_);
  not (_12078_, _12077_);
  not (_12079_, _11825_);
  not (_12080_, _11469_);
  and (_12081_, _12025_, _12080_);
  nor (_12082_, _12081_, _12079_);
  and (_12083_, _12082_, _12078_);
  and (_12084_, _12083_, _12055_);
  nor (_12085_, _12084_, _06807_);
  and (_12086_, _12084_, _06807_);
  nor (_12087_, _12086_, _12085_);
  nor (_12088_, _11971_, _11825_);
  not (_12090_, _11511_);
  and (_12091_, _12026_, _12090_);
  nor (_12092_, _12091_, _12088_);
  nor (_12093_, _12067_, _12064_);
  nor (_12094_, _12093_, _12068_);
  nor (_12095_, _12094_, _05898_);
  nor (_12096_, _12095_, _05944_);
  nor (_12097_, _12096_, _11937_);
  nor (_12098_, _12097_, _12065_);
  not (_12100_, _12098_);
  and (_12102_, _12100_, _11935_);
  and (_12103_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_12104_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_12105_, _12104_, _12103_);
  and (_12106_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_12107_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_12108_, _12107_, _12106_);
  and (_12109_, _12108_, _12105_);
  and (_12110_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_12112_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_12113_, _12112_, _12110_);
  and (_12114_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_12115_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_12116_, _12115_, _12114_);
  and (_12117_, _12116_, _12113_);
  and (_12118_, _12117_, _12109_);
  nor (_12119_, _12118_, _11986_);
  not (_12120_, _09341_);
  and (_12121_, _11986_, _12120_);
  nor (_12122_, _12121_, _12119_);
  not (_12123_, _12122_);
  and (_12124_, _12123_, _11972_);
  nor (_12125_, _12124_, _12102_);
  and (_12126_, _12125_, _12092_);
  nor (_12127_, _12126_, _06819_);
  and (_12128_, _12126_, _06819_);
  nor (_12129_, _12128_, _12127_);
  and (_12130_, _12129_, _12087_);
  not (_12131_, _11549_);
  and (_12132_, _12026_, _12131_);
  not (_12133_, _12025_);
  and (_12134_, _12088_, _12133_);
  nor (_12135_, _12134_, _12132_);
  nor (_12136_, _12063_, _12060_);
  nor (_12137_, _12136_, _12064_);
  nor (_12138_, _12137_, _05898_);
  nor (_12139_, _12138_, _05928_);
  nor (_12140_, _12139_, _11937_);
  nor (_12142_, _12140_, _12061_);
  not (_12143_, _12142_);
  and (_12144_, _12143_, _11935_);
  and (_12145_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_12146_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_12147_, _12146_, _12145_);
  and (_12148_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_12149_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_12150_, _12149_, _12148_);
  and (_12151_, _12150_, _12147_);
  and (_12152_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_12153_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_12154_, _12153_, _12152_);
  and (_12155_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_12156_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_12157_, _12156_, _12155_);
  and (_12158_, _12157_, _12154_);
  and (_12159_, _12158_, _12151_);
  nor (_12160_, _12159_, _11986_);
  not (_12161_, _06609_);
  and (_12162_, _11986_, _12161_);
  nor (_12163_, _12162_, _12160_);
  not (_12164_, _12163_);
  and (_12165_, _12164_, _11972_);
  nor (_12166_, _12165_, _12144_);
  and (_12167_, _12166_, _12135_);
  nor (_12168_, _12167_, _07767_);
  and (_12169_, _12167_, _07767_);
  nor (_12171_, _12169_, _12168_);
  not (_12172_, _09713_);
  and (_12173_, _12026_, _12172_);
  and (_12174_, _11968_, _11987_);
  nor (_12176_, _12174_, _12173_);
  and (_12177_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_12178_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_12180_, _12178_, _12177_);
  and (_12182_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_12183_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_12184_, _12183_, _12182_);
  and (_12185_, _12184_, _12180_);
  and (_12186_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_12187_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_12188_, _12187_, _12186_);
  and (_12189_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_12191_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_12192_, _12191_, _12189_);
  and (_12194_, _12192_, _12188_);
  and (_12195_, _12194_, _12185_);
  nor (_12196_, _12195_, _11986_);
  not (_12197_, _06993_);
  and (_12198_, _11986_, _12197_);
  nor (_12199_, _12198_, _12196_);
  not (_12201_, _12199_);
  and (_12202_, _12201_, _11972_);
  not (_12204_, _12202_);
  nor (_12205_, _12059_, _11955_);
  nor (_12207_, _12205_, _12060_);
  nor (_12208_, _12207_, _05898_);
  nor (_12209_, _12208_, _05902_);
  nor (_12210_, _12209_, _11937_);
  nor (_12212_, _12210_, _12057_);
  not (_12213_, _12212_);
  and (_12215_, _12213_, _11935_);
  and (_12216_, _11933_, _12079_);
  nor (_12218_, _12216_, _12215_);
  and (_12219_, _12218_, _12204_);
  and (_12221_, _12219_, _12176_);
  nor (_12222_, _12221_, _06364_);
  and (_12223_, _12221_, _06364_);
  nor (_12224_, _12223_, _12222_);
  and (_12225_, _12224_, _12171_);
  and (_12227_, _12225_, _12130_);
  and (_12228_, _12227_, _12033_);
  nor (_12230_, _06805_, _06013_);
  and (_12231_, _12230_, _12228_);
  and (_12233_, _12231_, _11800_);
  not (_12234_, _12233_);
  nor (_12236_, _11747_, _11827_);
  not (_12237_, _12236_);
  not (_12238_, _07792_);
  not (_12239_, _11799_);
  not (_12240_, _07687_);
  nor (_12241_, _06689_, _06687_);
  and (_12242_, _12241_, _11773_);
  nor (_12243_, _11793_, _08039_);
  and (_12244_, _12243_, _12242_);
  and (_12245_, _12244_, _12240_);
  and (_12246_, _12245_, _12239_);
  and (_12247_, _12246_, _07612_);
  and (_12248_, _12247_, _07368_);
  and (_12249_, _12248_, _12238_);
  not (_12250_, _12249_);
  nor (_12251_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_12252_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_12253_, _12252_, _12251_);
  nor (_12255_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_12256_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_12257_, _12256_, _12255_);
  and (_12258_, _12257_, _12253_);
  and (_12259_, _12258_, _11928_);
  not (_12260_, _12259_);
  and (_12262_, _11800_, _06118_);
  and (_12263_, _11797_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_12264_, _12263_, _12262_);
  and (_12266_, _12264_, _12260_);
  and (_12267_, _12266_, _12250_);
  and (_12268_, _11405_, _08764_);
  or (_12269_, _12268_, _11403_);
  and (_12270_, _11732_, _08764_);
  nor (_12271_, _12270_, _12269_);
  not (_12272_, _12271_);
  nor (_12273_, _12272_, _12267_);
  and (_12274_, _11405_, _08732_);
  nor (_12275_, _12274_, _11739_);
  and (_12276_, _11732_, _08732_);
  not (_12277_, _12276_);
  and (_12278_, _12277_, _11417_);
  and (_12279_, _12278_, _12275_);
  and (_12280_, _12279_, _11398_);
  and (_12282_, _12280_, _12267_);
  nor (_12283_, _12282_, _12273_);
  nor (_12284_, _11738_, _11734_);
  and (_12285_, _12284_, _11895_);
  not (_12286_, _12285_);
  nor (_12288_, _12286_, _12283_);
  nor (_12289_, _12288_, _11730_);
  nor (_12291_, _12289_, _12237_);
  not (_12292_, _08941_);
  and (_12294_, _11928_, _12292_);
  nor (_12295_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_12296_, _12295_, _08985_);
  and (_12297_, _12296_, _10935_);
  not (_12298_, _12297_);
  and (_12299_, _12298_, _11797_);
  nor (_12301_, _12299_, _12294_);
  not (_12302_, _12301_);
  nor (_12304_, _12302_, _12291_);
  and (_12305_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_12306_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_12307_, _12306_, _12305_);
  and (_12308_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_12309_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_12310_, _12309_, _12308_);
  and (_12311_, _12310_, _12307_);
  and (_12312_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_12313_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_12314_, _12313_, _12312_);
  and (_12316_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_12317_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_12318_, _12317_, _12316_);
  and (_12319_, _12318_, _12314_);
  and (_12320_, _12319_, _12311_);
  nor (_12321_, _12320_, _11986_);
  and (_12322_, _11986_, _07978_);
  nor (_12323_, _12322_, _12321_);
  not (_12324_, _12323_);
  and (_12325_, _12324_, _11972_);
  and (_12326_, _12026_, _11689_);
  nor (_12328_, _12326_, _12325_);
  nor (_12329_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_12330_, _12329_, _11952_);
  nor (_12332_, _12330_, _05898_);
  nor (_12333_, _12332_, _05998_);
  nor (_12335_, _12333_, _11937_);
  nor (_12336_, _12335_, _11950_);
  not (_12337_, _12336_);
  and (_12338_, _12337_, _11935_);
  and (_12339_, _11968_, _08753_);
  nor (_12340_, _12339_, _12338_);
  and (_12341_, _12340_, _12328_);
  and (_12343_, _12341_, _06030_);
  nor (_12344_, _12341_, _06030_);
  or (_12346_, _12344_, _12343_);
  nor (_12347_, _12346_, _06827_);
  and (_12348_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_12349_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_12350_, _12349_, _12348_);
  and (_12351_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_12352_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_12353_, _12352_, _12351_);
  and (_12354_, _12353_, _12350_);
  and (_12355_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_12356_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_12357_, _12356_, _12355_);
  and (_12359_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_12360_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_12362_, _12360_, _12359_);
  and (_12363_, _12362_, _12357_);
  and (_12364_, _12363_, _12354_);
  nor (_12365_, _12364_, _11986_);
  and (_12366_, _11986_, _11023_);
  nor (_12368_, _12366_, _12365_);
  not (_12369_, _12368_);
  and (_12370_, _12369_, _11972_);
  and (_12371_, _11971_, _12079_);
  nor (_12372_, _11952_, _11948_);
  nor (_12374_, _12372_, _11953_);
  nor (_12375_, _12374_, _05898_);
  nor (_12376_, _12375_, _05985_);
  nor (_12377_, _12376_, _11937_);
  nor (_12378_, _12377_, _11947_);
  not (_12379_, _12378_);
  and (_12380_, _12379_, _11935_);
  or (_12381_, _12380_, _12371_);
  and (_12382_, _12026_, _11651_);
  and (_12383_, _11968_, _08725_);
  or (_12384_, _12383_, _12382_);
  or (_12385_, _12384_, _12381_);
  nor (_12386_, _12385_, _12370_);
  nor (_12387_, _12386_, _05993_);
  and (_12388_, _12386_, _05993_);
  nor (_12389_, _12388_, _12387_);
  nor (_12390_, _11953_, _11945_);
  nor (_12391_, _12390_, _11954_);
  nor (_12393_, _12391_, _05898_);
  nor (_12394_, _12393_, _05972_);
  nor (_12395_, _12394_, _11937_);
  nor (_12397_, _12395_, _11944_);
  not (_12398_, _12397_);
  and (_12399_, _12398_, _11935_);
  not (_12400_, _12399_);
  and (_12401_, _11968_, _11392_);
  and (_12402_, _12000_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_12403_, _11990_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_12404_, _12403_, _12402_);
  and (_12405_, _12009_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_12406_, _12004_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_12407_, _12406_, _12405_);
  and (_12408_, _12407_, _12404_);
  and (_12409_, _12006_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_12410_, _12011_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_12411_, _12410_, _12409_);
  and (_12412_, _11997_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_12413_, _11993_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_12414_, _12413_, _12412_);
  and (_12416_, _12414_, _12411_);
  and (_12417_, _12416_, _12408_);
  nor (_12418_, _12417_, _11986_);
  and (_12419_, _11986_, _06435_);
  nor (_12420_, _12419_, _12418_);
  not (_12421_, _12420_);
  and (_12422_, _12421_, _11972_);
  and (_12423_, _12026_, _11628_);
  or (_12424_, _12423_, _12422_);
  nor (_12425_, _12424_, _12401_);
  and (_12426_, _12425_, _12400_);
  nor (_12427_, _12426_, _05981_);
  and (_12428_, _12426_, _05981_);
  nor (_12429_, _12428_, _12427_);
  nor (_12430_, _12429_, _12389_);
  and (_12431_, _12430_, _12347_);
  and (_12432_, _12431_, _12228_);
  nor (_12433_, _05967_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_12434_, _12433_, _12432_);
  not (_12435_, _12434_);
  and (_12436_, _12435_, _12304_);
  and (_12437_, _12436_, _12234_);
  not (_12438_, _11748_);
  and (_12439_, _07494_, _07479_);
  not (_12441_, _12439_);
  and (_12442_, _07495_, _06715_);
  and (_12443_, _12442_, _12441_);
  not (_12444_, _12443_);
  and (_12445_, _07920_, _07344_);
  not (_12446_, _12445_);
  nor (_12447_, _07442_, _06302_);
  and (_12449_, _07573_, _06660_);
  nor (_12450_, _12449_, _06120_);
  nor (_12451_, _12450_, _12447_);
  and (_12452_, _12451_, _06701_);
  nor (_12453_, _12451_, _06701_);
  nor (_12454_, _12453_, _12452_);
  and (_12455_, _12454_, _06145_);
  and (_12456_, _06701_, _06349_);
  nor (_12457_, _06187_, _06128_);
  and (_12458_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_12459_, _12458_, _12457_);
  or (_12460_, _12459_, _06779_);
  nor (_12462_, _12460_, _12456_);
  not (_12463_, _12462_);
  nor (_12464_, _12463_, _12455_);
  and (_12465_, _12464_, _12446_);
  and (_12466_, _12465_, _12444_);
  nor (_12467_, _12466_, _12438_);
  and (_12469_, _11750_, _11743_);
  and (_12470_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_12472_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12473_, _12472_, _12470_);
  and (_12474_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12475_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12476_, _12475_, _12474_);
  and (_12477_, _12476_, _11722_);
  and (_12478_, _12477_, _12473_);
  and (_12479_, _12478_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12480_, _12478_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12481_, _12480_, _12479_);
  and (_12482_, _12481_, _12469_);
  and (_12483_, _12024_, _11424_);
  and (_12484_, _11749_, _11455_);
  and (_12485_, _12484_, _11743_);
  and (_12486_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_12487_, _12486_, _12483_);
  or (_12488_, _12487_, _12482_);
  nor (_12489_, _12488_, _12467_);
  nand (_12491_, _12489_, _12437_);
  or (_12492_, _12491_, _11792_);
  or (_12493_, _12492_, _11753_);
  not (_12494_, _06530_);
  and (_12495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12498_, _12497_, _12495_);
  and (_12499_, _12498_, _11250_);
  and (_12500_, _12499_, _12494_);
  and (_12501_, _12500_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12503_, _12502_, _12501_);
  nor (_12504_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12505_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_12506_, _12505_, _12504_);
  or (_12507_, _12506_, _12437_);
  and (_12508_, _12507_, _06071_);
  and (_11409_, _12508_, _12493_);
  nor (_11432_, _12368_, rst);
  or (_12509_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  nand (_12510_, _06530_, _10995_);
  and (_12511_, _12510_, _06071_);
  and (_11437_, _12511_, _12509_);
  or (_12512_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_12513_, _06530_, _05739_);
  and (_12514_, _12513_, _06071_);
  and (_11440_, _12514_, _12512_);
  and (_11443_, _08725_, _06071_);
  nor (_12515_, _06993_, _06996_);
  and (_12516_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_12517_, _12516_, _06390_);
  or (_12518_, _12517_, _12515_);
  or (_12519_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_12520_, _12519_, _06071_);
  and (_11489_, _12520_, _12518_);
  or (_12521_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_12522_, _06530_, _05693_);
  and (_12523_, _12522_, _06071_);
  and (_11494_, _12523_, _12521_);
  and (_12524_, _06071_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_12525_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_12527_, _11874_, _11731_);
  or (_12528_, _12527_, _11908_);
  or (_12529_, _11879_, _11852_);
  and (_12530_, _12529_, _11810_);
  or (_12531_, _12530_, _12528_);
  and (_12532_, _08761_, _08764_);
  and (_12533_, _11831_, _11810_);
  or (_12534_, _12533_, _11844_);
  and (_12535_, _11805_, _08728_);
  or (_12536_, _12535_, _12534_);
  or (_12537_, _12536_, _12532_);
  or (_12538_, _12537_, _12531_);
  or (_12539_, _11864_, _11859_);
  or (_12540_, _12539_, _11834_);
  and (_12541_, _11889_, _11736_);
  and (_12542_, _11889_, _11407_);
  or (_12543_, _12542_, _12541_);
  or (_12544_, _12543_, _11854_);
  or (_12545_, _12544_, _12540_);
  not (_12546_, _11398_);
  and (_12547_, _11805_, _11810_);
  and (_12548_, _11810_, _11414_);
  and (_12549_, _11810_, _08765_);
  or (_12550_, _12549_, _12548_);
  or (_12551_, _12550_, _12547_);
  or (_12552_, _12551_, _12546_);
  or (_12553_, _12552_, _12545_);
  or (_12555_, _12553_, _12538_);
  and (_12556_, _12555_, _08775_);
  or (_11499_, _12556_, _12525_);
  and (_12558_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _06071_);
  and (_11502_, _12558_, _05811_);
  and (_12559_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_12561_, _08865_, _06609_);
  or (_12562_, _12561_, _12559_);
  and (_11544_, _12562_, _06071_);
  and (_12563_, _08254_, word_in[0]);
  nand (_12564_, _08174_, _09175_);
  or (_12565_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_12566_, _12565_, _12564_);
  and (_12567_, _12566_, _08196_);
  or (_12568_, _12567_, _08184_);
  nand (_12569_, _08174_, _09726_);
  or (_12570_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_12571_, _12570_, _12569_);
  and (_12572_, _12571_, _08221_);
  nand (_12573_, _08174_, _09936_);
  or (_12574_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_12575_, _12574_, _12573_);
  and (_12576_, _12575_, _08200_);
  nand (_12577_, _08174_, _09476_);
  or (_12578_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_12579_, _12578_, _12577_);
  and (_12580_, _12579_, _08208_);
  or (_12581_, _12580_, _12576_);
  or (_12582_, _12581_, _12572_);
  or (_12583_, _12582_, _12568_);
  nand (_12584_, _08174_, _10161_);
  or (_12585_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_12586_, _12585_, _12584_);
  and (_12587_, _12586_, _08196_);
  or (_12588_, _12587_, _08281_);
  nand (_12589_, _08174_, _10589_);
  or (_12590_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12591_, _12590_, _12589_);
  and (_12592_, _12591_, _08221_);
  nand (_12593_, _08174_, _10795_);
  or (_12594_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12595_, _12594_, _12593_);
  and (_12596_, _12595_, _08200_);
  nand (_12597_, _08174_, _10371_);
  or (_12598_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_12599_, _12598_, _12597_);
  and (_12601_, _12599_, _08208_);
  or (_12602_, _12601_, _12596_);
  or (_12603_, _12602_, _12592_);
  or (_12604_, _12603_, _12588_);
  and (_12605_, _12604_, _12583_);
  and (_12606_, _12605_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12606_, _12563_);
  and (_12607_, _08254_, word_in[1]);
  nand (_12608_, _08174_, _09490_);
  or (_12609_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_12610_, _12609_, _12608_);
  and (_12611_, _12610_, _08208_);
  or (_12612_, _12611_, _08184_);
  nand (_12613_, _08174_, _09740_);
  or (_12614_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_12615_, _12614_, _12613_);
  and (_12616_, _12615_, _08221_);
  nand (_12617_, _08174_, _09950_);
  or (_12618_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_12619_, _12618_, _12617_);
  and (_12620_, _12619_, _08200_);
  nand (_12621_, _08174_, _09197_);
  or (_12622_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_12623_, _12622_, _12621_);
  and (_12625_, _12623_, _08196_);
  or (_12626_, _12625_, _12620_);
  or (_12627_, _12626_, _12616_);
  or (_12628_, _12627_, _12612_);
  nand (_12629_, _08174_, _10387_);
  or (_12630_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_12631_, _12630_, _12629_);
  and (_12632_, _12631_, _08208_);
  or (_12633_, _12632_, _08281_);
  nand (_12634_, _08174_, _10809_);
  or (_12635_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_12636_, _12635_, _12634_);
  and (_12637_, _12636_, _08200_);
  nand (_12638_, _08174_, _10606_);
  or (_12639_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_12640_, _12639_, _12638_);
  and (_12641_, _12640_, _08221_);
  or (_12642_, _12641_, _12637_);
  nand (_12643_, _08174_, _10177_);
  or (_12644_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_12645_, _12644_, _12643_);
  and (_12646_, _12645_, _08196_);
  or (_12647_, _12646_, _12642_);
  or (_12648_, _12647_, _12633_);
  and (_12649_, _12648_, _12628_);
  and (_12650_, _12649_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12650_, _12607_);
  and (_12651_, _08254_, word_in[2]);
  nand (_12652_, _08174_, _09502_);
  or (_12653_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_12654_, _12653_, _12652_);
  and (_12655_, _12654_, _08208_);
  or (_12656_, _12655_, _08184_);
  nand (_12657_, _08174_, _09752_);
  or (_12658_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_12659_, _12658_, _12657_);
  and (_12660_, _12659_, _08221_);
  nand (_12661_, _08174_, _09965_);
  or (_12662_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_12663_, _12662_, _12661_);
  and (_12664_, _12663_, _08200_);
  nand (_12665_, _08174_, _09208_);
  or (_12666_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_12667_, _12666_, _12665_);
  and (_12668_, _12667_, _08196_);
  or (_12669_, _12668_, _12664_);
  or (_12670_, _12669_, _12660_);
  or (_12671_, _12670_, _12656_);
  nand (_12672_, _08174_, _10399_);
  or (_12673_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_12674_, _12673_, _12672_);
  and (_12675_, _12674_, _08208_);
  or (_12676_, _12675_, _08281_);
  nand (_12677_, _08174_, _10820_);
  or (_12678_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_12679_, _12678_, _12677_);
  and (_12680_, _12679_, _08200_);
  nand (_12681_, _08174_, _10619_);
  or (_12682_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_12683_, _12682_, _12681_);
  and (_12684_, _12683_, _08221_);
  or (_12685_, _12684_, _12680_);
  nand (_12686_, _08174_, _10195_);
  or (_12687_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_12688_, _12687_, _12686_);
  and (_12689_, _12688_, _08196_);
  or (_12690_, _12689_, _12685_);
  or (_12691_, _12690_, _12676_);
  and (_12692_, _12691_, _12671_);
  and (_12693_, _12692_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12693_, _12651_);
  and (_12695_, _08254_, word_in[3]);
  nand (_12696_, _08174_, _09513_);
  or (_12697_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_12698_, _12697_, _12696_);
  and (_12699_, _12698_, _08208_);
  or (_12700_, _12699_, _08184_);
  nand (_12701_, _08174_, _09764_);
  or (_12702_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_12703_, _12702_, _12701_);
  and (_12704_, _12703_, _08221_);
  nand (_12705_, _08174_, _09976_);
  or (_12706_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_12707_, _12706_, _12705_);
  and (_12708_, _12707_, _08200_);
  nand (_12709_, _08174_, _09258_);
  or (_12710_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_12711_, _12710_, _12709_);
  and (_12712_, _12711_, _08196_);
  or (_12713_, _12712_, _12708_);
  or (_12714_, _12713_, _12704_);
  or (_12715_, _12714_, _12700_);
  nand (_12716_, _08174_, _10412_);
  or (_12717_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_12718_, _12717_, _12716_);
  and (_12719_, _12718_, _08208_);
  or (_12720_, _12719_, _08281_);
  nand (_12721_, _08174_, _10838_);
  or (_12722_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_12723_, _12722_, _12721_);
  and (_12724_, _12723_, _08200_);
  nand (_12725_, _08174_, _10631_);
  or (_12726_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_12727_, _12726_, _12725_);
  and (_12728_, _12727_, _08221_);
  or (_12729_, _12728_, _12724_);
  nand (_12730_, _08174_, _10208_);
  or (_12731_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_12732_, _12731_, _12730_);
  and (_12733_, _12732_, _08196_);
  or (_12734_, _12733_, _12729_);
  or (_12735_, _12734_, _12720_);
  and (_12736_, _12735_, _12715_);
  and (_12737_, _12736_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _12737_, _12695_);
  and (_12738_, _08254_, word_in[4]);
  nand (_12739_, _08174_, _09275_);
  or (_12740_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_12741_, _12740_, _12739_);
  and (_12742_, _12741_, _08196_);
  or (_12743_, _12742_, _08184_);
  nand (_12744_, _08174_, _09776_);
  or (_12745_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_12746_, _12745_, _12744_);
  and (_12747_, _12746_, _08221_);
  nand (_12748_, _08174_, _09991_);
  or (_12749_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_12750_, _12749_, _12748_);
  and (_12751_, _12750_, _08200_);
  nand (_12752_, _08174_, _09525_);
  or (_12753_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_12754_, _12753_, _12752_);
  and (_12755_, _12754_, _08208_);
  or (_12756_, _12755_, _12751_);
  or (_12757_, _12756_, _12747_);
  or (_12758_, _12757_, _12743_);
  nand (_12759_, _08174_, _10220_);
  or (_12760_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_12761_, _12760_, _12759_);
  and (_12762_, _12761_, _08196_);
  or (_12763_, _12762_, _08281_);
  nand (_12764_, _08174_, _10643_);
  or (_12765_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_12766_, _12765_, _12764_);
  and (_12767_, _12766_, _08221_);
  nand (_12768_, _08174_, _10850_);
  or (_12769_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_12770_, _12769_, _12768_);
  and (_12771_, _12770_, _08200_);
  nand (_12772_, _08174_, _10425_);
  or (_12773_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_12774_, _12773_, _12772_);
  and (_12775_, _12774_, _08208_);
  or (_12776_, _12775_, _12771_);
  or (_12777_, _12776_, _12767_);
  or (_12778_, _12777_, _12763_);
  and (_12779_, _12778_, _12758_);
  and (_12780_, _12779_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _12780_, _12738_);
  and (_12781_, _08254_, word_in[5]);
  nand (_12782_, _08174_, _09295_);
  or (_12783_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_12784_, _12783_, _12782_);
  and (_12785_, _12784_, _08196_);
  or (_12786_, _12785_, _08184_);
  nand (_12787_, _08174_, _09787_);
  or (_12788_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_12789_, _12788_, _12787_);
  and (_12790_, _12789_, _08221_);
  nand (_12791_, _08174_, _10008_);
  or (_12792_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_12793_, _12792_, _12791_);
  and (_12794_, _12793_, _08200_);
  nand (_12795_, _08174_, _09538_);
  or (_12796_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_12797_, _12796_, _12795_);
  and (_12798_, _12797_, _08208_);
  or (_12799_, _12798_, _12794_);
  or (_12800_, _12799_, _12790_);
  or (_12801_, _12800_, _12786_);
  nand (_12802_, _08174_, _10232_);
  or (_12803_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_12804_, _12803_, _12802_);
  and (_12805_, _12804_, _08196_);
  or (_12806_, _12805_, _08281_);
  nand (_12807_, _08174_, _10654_);
  or (_12808_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_12809_, _12808_, _12807_);
  and (_12810_, _12809_, _08221_);
  nand (_12811_, _08174_, _10862_);
  or (_12812_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_12813_, _12812_, _12811_);
  and (_12814_, _12813_, _08200_);
  nand (_12815_, _08174_, _10441_);
  or (_12816_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_12817_, _12816_, _12815_);
  and (_12818_, _12817_, _08208_);
  or (_12819_, _12818_, _12814_);
  or (_12820_, _12819_, _12810_);
  or (_12821_, _12820_, _12806_);
  and (_12822_, _12821_, _12801_);
  and (_12823_, _12822_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _12823_, _12781_);
  and (_12824_, _08254_, word_in[6]);
  nand (_12825_, _08174_, _09313_);
  or (_12826_, _08174_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_12827_, _12826_, _12825_);
  and (_12828_, _12827_, _08196_);
  or (_12829_, _12828_, _08184_);
  nand (_12830_, _08174_, _09800_);
  or (_12831_, _08174_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_12832_, _12831_, _12830_);
  and (_12833_, _12832_, _08221_);
  nand (_12834_, _08174_, _10019_);
  or (_12835_, _08174_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_12836_, _12835_, _12834_);
  and (_12837_, _12836_, _08200_);
  nand (_12838_, _08174_, _09550_);
  or (_12839_, _08174_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_12840_, _12839_, _12838_);
  and (_12841_, _12840_, _08208_);
  or (_12842_, _12841_, _12837_);
  or (_12843_, _12842_, _12833_);
  or (_12844_, _12843_, _12829_);
  nand (_12845_, _08174_, _10244_);
  or (_12846_, _08174_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_12847_, _12846_, _12845_);
  and (_12848_, _12847_, _08196_);
  or (_12849_, _12848_, _08281_);
  nand (_12850_, _08174_, _10667_);
  or (_12851_, _08174_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_12852_, _12851_, _12850_);
  and (_12853_, _12852_, _08221_);
  nand (_12854_, _08174_, _10874_);
  or (_12855_, _08174_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_12856_, _12855_, _12854_);
  and (_12857_, _12856_, _08200_);
  nand (_12858_, _08174_, _10454_);
  or (_12859_, _08174_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_12860_, _12859_, _12858_);
  and (_12861_, _12860_, _08208_);
  or (_12862_, _12861_, _12857_);
  or (_12863_, _12862_, _12853_);
  or (_12864_, _12863_, _12849_);
  and (_12865_, _12864_, _12844_);
  and (_12866_, _12865_, _08253_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _12866_, _12824_);
  and (_12867_, _08357_, word_in[8]);
  nand (_12868_, _08174_, _09369_);
  or (_12869_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_12870_, _12869_, _12868_);
  and (_12871_, _12870_, _08359_);
  nand (_12872_, _08174_, _09047_);
  or (_12873_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_12874_, _12873_, _12872_);
  and (_12875_, _12874_, _08358_);
  or (_12876_, _12875_, _12871_);
  and (_12877_, _12876_, _08321_);
  nand (_12878_, _08174_, _10269_);
  or (_12879_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_12880_, _12879_, _12878_);
  and (_12881_, _12880_, _08359_);
  nand (_12882_, _08174_, _10050_);
  or (_12883_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_12884_, _12883_, _12882_);
  and (_12885_, _12884_, _08358_);
  or (_12886_, _12885_, _12881_);
  and (_12887_, _12886_, _08323_);
  nand (_12888_, _08174_, _09825_);
  or (_12889_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_12890_, _12889_, _12888_);
  and (_12891_, _12890_, _08359_);
  nand (_12892_, _08174_, _09593_);
  or (_12893_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _08358_);
  or (_12896_, _12895_, _12891_);
  and (_12897_, _12896_, _08346_);
  nand (_12898_, _08174_, _10700_);
  or (_12899_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_12900_, _12899_, _12898_);
  and (_12901_, _12900_, _08359_);
  nand (_12902_, _08174_, _10484_);
  or (_12903_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_12904_, _12903_, _12902_);
  and (_12905_, _12904_, _08358_);
  or (_12906_, _12905_, _12901_);
  and (_12908_, _12906_, _08350_);
  or (_12909_, _12908_, _12897_);
  or (_12910_, _12909_, _12887_);
  nor (_12911_, _12910_, _12877_);
  nor (_12912_, _12911_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _12912_, _12867_);
  and (_12913_, _08357_, word_in[9]);
  nand (_12914_, _08174_, _09386_);
  or (_12915_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_12916_, _12915_, _12914_);
  and (_12918_, _12916_, _08359_);
  nand (_12919_, _08174_, _09078_);
  or (_12920_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_12921_, _12920_, _12919_);
  and (_12922_, _12921_, _08358_);
  or (_12923_, _12922_, _12918_);
  and (_12924_, _12923_, _08321_);
  nand (_12925_, _08174_, _10285_);
  or (_12926_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_12927_, _12926_, _12925_);
  and (_12928_, _12927_, _08359_);
  nand (_12929_, _08174_, _10066_);
  or (_12930_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _08358_);
  or (_12933_, _12932_, _12928_);
  and (_12934_, _12933_, _08323_);
  nand (_12935_, _08174_, _09841_);
  or (_12936_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_12937_, _12936_, _12935_);
  and (_12938_, _12937_, _08359_);
  nand (_12939_, _08174_, _09611_);
  or (_12940_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_12941_, _12940_, _12939_);
  and (_12942_, _12941_, _08358_);
  or (_12943_, _12942_, _12938_);
  and (_12944_, _12943_, _08346_);
  nand (_12945_, _08174_, _10712_);
  or (_12946_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_12947_, _12946_, _12945_);
  and (_12948_, _12947_, _08359_);
  nand (_12949_, _08174_, _10501_);
  or (_12950_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _08358_);
  or (_12953_, _12952_, _12948_);
  and (_12954_, _12953_, _08350_);
  or (_12955_, _12954_, _12944_);
  or (_12956_, _12955_, _12934_);
  nor (_12957_, _12956_, _12924_);
  nor (_12958_, _12957_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _12958_, _12913_);
  and (_12959_, _08357_, word_in[10]);
  nand (_12960_, _08174_, _09400_);
  or (_12961_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_12962_, _12961_, _12960_);
  and (_12963_, _12962_, _08359_);
  nand (_12964_, _08174_, _09093_);
  or (_12965_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_12966_, _12965_, _12964_);
  and (_12967_, _12966_, _08358_);
  or (_12968_, _12967_, _12963_);
  and (_12969_, _12968_, _08321_);
  nand (_12970_, _08174_, _10298_);
  or (_12971_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_12972_, _12971_, _12970_);
  and (_12973_, _12972_, _08359_);
  nand (_12974_, _08174_, _10079_);
  or (_12975_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_12976_, _12975_, _12974_);
  and (_12977_, _12976_, _08358_);
  or (_12978_, _12977_, _12973_);
  and (_12979_, _12978_, _08323_);
  nand (_12980_, _08174_, _09853_);
  or (_12981_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_12982_, _12981_, _12980_);
  and (_12983_, _12982_, _08359_);
  nand (_12984_, _08174_, _09623_);
  or (_12985_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_12986_, _12985_, _12984_);
  and (_12987_, _12986_, _08358_);
  or (_12988_, _12987_, _12983_);
  and (_12989_, _12988_, _08346_);
  nand (_12990_, _08174_, _10724_);
  or (_12991_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_12992_, _12991_, _12990_);
  and (_12993_, _12992_, _08359_);
  nand (_12994_, _08174_, _10513_);
  or (_12995_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_12996_, _12995_, _12994_);
  and (_12998_, _12996_, _08358_);
  or (_12999_, _12998_, _12993_);
  and (_13000_, _12999_, _08350_);
  or (_13001_, _13000_, _12989_);
  or (_13002_, _13001_, _12979_);
  nor (_13003_, _13002_, _12969_);
  nor (_13004_, _13003_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13004_, _12959_);
  and (_13005_, _08357_, word_in[11]);
  nand (_13006_, _08174_, _09413_);
  or (_13007_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_13008_, _13007_, _13006_);
  and (_13009_, _13008_, _08359_);
  nand (_13010_, _08174_, _09105_);
  or (_13011_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_13012_, _13011_, _13010_);
  and (_13013_, _13012_, _08358_);
  or (_13014_, _13013_, _13009_);
  and (_13015_, _13014_, _08321_);
  nand (_13016_, _08174_, _10310_);
  or (_13017_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_13018_, _13017_, _13016_);
  and (_13019_, _13018_, _08359_);
  nand (_13020_, _08174_, _10095_);
  or (_13021_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_13022_, _13021_, _13020_);
  and (_13023_, _13022_, _08358_);
  or (_13024_, _13023_, _13019_);
  and (_13025_, _13024_, _08323_);
  nand (_13026_, _08174_, _09865_);
  or (_13027_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _08359_);
  nand (_13030_, _08174_, _09636_);
  or (_13031_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_13032_, _13031_, _13030_);
  and (_13033_, _13032_, _08358_);
  or (_13035_, _13033_, _13029_);
  and (_13036_, _13035_, _08346_);
  nand (_13037_, _08174_, _10736_);
  or (_13038_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_13039_, _13038_, _13037_);
  and (_13040_, _13039_, _08359_);
  nand (_13041_, _08174_, _10525_);
  or (_13042_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_13043_, _13042_, _13041_);
  and (_13044_, _13043_, _08358_);
  or (_13045_, _13044_, _13040_);
  and (_13046_, _13045_, _08350_);
  or (_13047_, _13046_, _13036_);
  or (_13048_, _13047_, _13025_);
  nor (_13049_, _13048_, _13015_);
  nor (_13050_, _13049_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13050_, _13005_);
  and (_13051_, _08357_, word_in[12]);
  nand (_13052_, _08174_, _09424_);
  or (_13053_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_13054_, _13053_, _13052_);
  and (_13055_, _13054_, _08359_);
  nand (_13057_, _08174_, _09120_);
  or (_13058_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_13059_, _13058_, _13057_);
  and (_13060_, _13059_, _08358_);
  or (_13061_, _13060_, _13055_);
  and (_13062_, _13061_, _08321_);
  nand (_13063_, _08174_, _10323_);
  or (_13064_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_13065_, _13064_, _13063_);
  and (_13066_, _13065_, _08359_);
  nand (_13067_, _08174_, _10110_);
  or (_13068_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_13069_, _13068_, _13067_);
  and (_13070_, _13069_, _08358_);
  or (_13071_, _13070_, _13066_);
  and (_13072_, _13071_, _08323_);
  nand (_13073_, _08174_, _09878_);
  or (_13074_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_13075_, _13074_, _13073_);
  and (_13076_, _13075_, _08359_);
  nand (_13077_, _08174_, _09648_);
  or (_13078_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_13079_, _13078_, _13077_);
  and (_13080_, _13079_, _08358_);
  or (_13081_, _13080_, _13076_);
  and (_13082_, _13081_, _08346_);
  nand (_13083_, _08174_, _10747_);
  or (_13084_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_13086_, _13084_, _13083_);
  and (_13087_, _13086_, _08359_);
  nand (_13088_, _08174_, _10537_);
  or (_13089_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_13090_, _13089_, _13088_);
  and (_13091_, _13090_, _08358_);
  or (_13092_, _13091_, _13087_);
  and (_13093_, _13092_, _08350_);
  or (_13094_, _13093_, _13082_);
  or (_13095_, _13094_, _13072_);
  nor (_13096_, _13095_, _13062_);
  nor (_13097_, _13096_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13097_, _13051_);
  and (_13099_, _08357_, word_in[13]);
  nand (_13100_, _08174_, _09435_);
  or (_13101_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_13102_, _13101_, _13100_);
  and (_13103_, _13102_, _08359_);
  nand (_13104_, _08174_, _09131_);
  or (_13105_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _08358_);
  or (_13108_, _13107_, _13103_);
  and (_13109_, _13108_, _08321_);
  nand (_13111_, _08174_, _10334_);
  or (_13112_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_13113_, _13112_, _13111_);
  and (_13114_, _13113_, _08359_);
  nand (_13115_, _08174_, _10121_);
  or (_13116_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_13117_, _13116_, _13115_);
  and (_13118_, _13117_, _08358_);
  or (_13119_, _13118_, _13114_);
  and (_13120_, _13119_, _08323_);
  nand (_13121_, _08174_, _09891_);
  or (_13122_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_13123_, _13122_, _13121_);
  and (_13124_, _13123_, _08359_);
  nand (_13125_, _08174_, _09661_);
  or (_13126_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_13127_, _13126_, _13125_);
  and (_13128_, _13127_, _08358_);
  or (_13129_, _13128_, _13124_);
  and (_13130_, _13129_, _08346_);
  nand (_13131_, _08174_, _10761_);
  or (_13132_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_13133_, _13132_, _13131_);
  and (_13134_, _13133_, _08359_);
  nand (_13135_, _08174_, _10549_);
  or (_13136_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_13137_, _13136_, _13135_);
  and (_13138_, _13137_, _08358_);
  or (_13139_, _13138_, _13134_);
  and (_13140_, _13139_, _08350_);
  or (_13141_, _13140_, _13130_);
  or (_13142_, _13141_, _13120_);
  nor (_13143_, _13142_, _13109_);
  nor (_13144_, _13143_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13144_, _13099_);
  and (_13145_, _08357_, word_in[14]);
  nand (_13146_, _08174_, _09448_);
  or (_13147_, _08174_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_13148_, _13147_, _13146_);
  and (_13149_, _13148_, _08359_);
  nand (_13150_, _08174_, _09144_);
  or (_13151_, _08174_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_13152_, _13151_, _13150_);
  and (_13153_, _13152_, _08358_);
  or (_13154_, _13153_, _13149_);
  and (_13155_, _13154_, _08321_);
  nand (_13156_, _08174_, _10346_);
  or (_13157_, _08174_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_13158_, _13157_, _13156_);
  and (_13159_, _13158_, _08359_);
  nand (_13160_, _08174_, _10134_);
  or (_13161_, _08174_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_13162_, _13161_, _13160_);
  and (_13163_, _13162_, _08358_);
  or (_13164_, _13163_, _13159_);
  and (_13165_, _13164_, _08323_);
  nand (_13166_, _08174_, _09910_);
  or (_13167_, _08174_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_13168_, _13167_, _13166_);
  and (_13169_, _13168_, _08359_);
  nand (_13170_, _08174_, _09673_);
  or (_13171_, _08174_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_13172_, _13171_, _13170_);
  and (_13173_, _13172_, _08358_);
  or (_13174_, _13173_, _13169_);
  and (_13175_, _13174_, _08346_);
  nand (_13176_, _08174_, _10773_);
  or (_13177_, _08174_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_13178_, _13177_, _13176_);
  and (_13179_, _13178_, _08359_);
  nand (_13180_, _08174_, _10561_);
  or (_13181_, _08174_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_13182_, _13181_, _13180_);
  and (_13183_, _13182_, _08358_);
  or (_13184_, _13183_, _13179_);
  and (_13185_, _13184_, _08350_);
  or (_13186_, _13185_, _13175_);
  or (_13187_, _13186_, _13165_);
  nor (_13188_, _13187_, _13155_);
  nor (_13189_, _13188_, _08357_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13189_, _13145_);
  and (_13190_, _08450_, word_in[16]);
  and (_13191_, _12579_, _08196_);
  and (_13192_, _12566_, _08200_);
  or (_13193_, _13192_, _13191_);
  and (_13194_, _12575_, _08221_);
  and (_13195_, _12571_, _08208_);
  or (_13196_, _13195_, _13194_);
  or (_13197_, _13196_, _13193_);
  or (_13198_, _13197_, _08419_);
  and (_13199_, _12595_, _08221_);
  and (_13200_, _12599_, _08196_);
  or (_13201_, _13200_, _13199_);
  and (_13202_, _12591_, _08208_);
  and (_13203_, _12586_, _08200_);
  or (_13204_, _13203_, _13202_);
  or (_13205_, _13204_, _13201_);
  or (_13207_, _13205_, _08460_);
  nand (_13208_, _13207_, _13198_);
  nor (_13209_, _13208_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13209_, _13190_);
  and (_13210_, _08450_, word_in[17]);
  and (_13211_, _12623_, _08200_);
  and (_13212_, _12610_, _08196_);
  or (_13213_, _13212_, _13211_);
  and (_13214_, _12615_, _08208_);
  and (_13215_, _12619_, _08221_);
  or (_13216_, _13215_, _13214_);
  or (_13217_, _13216_, _13213_);
  or (_13218_, _13217_, _08419_);
  and (_13219_, _12636_, _08221_);
  and (_13220_, _12631_, _08196_);
  or (_13221_, _13220_, _13219_);
  and (_13222_, _12640_, _08208_);
  and (_13223_, _12645_, _08200_);
  or (_13224_, _13223_, _13222_);
  or (_13225_, _13224_, _13221_);
  or (_13226_, _13225_, _08460_);
  nand (_13227_, _13226_, _13218_);
  nor (_13228_, _13227_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13228_, _13210_);
  and (_13229_, _08450_, word_in[18]);
  and (_13230_, _12663_, _08221_);
  and (_13231_, _12654_, _08196_);
  or (_13232_, _13231_, _13230_);
  and (_13233_, _12659_, _08208_);
  and (_13234_, _12667_, _08200_);
  or (_13235_, _13234_, _13233_);
  or (_13236_, _13235_, _13232_);
  or (_13237_, _13236_, _08419_);
  and (_13238_, _12674_, _08196_);
  and (_13239_, _12688_, _08200_);
  or (_13240_, _13239_, _13238_);
  and (_13241_, _12679_, _08221_);
  and (_13242_, _12683_, _08208_);
  or (_13243_, _13242_, _13241_);
  or (_13244_, _13243_, _13240_);
  or (_13245_, _13244_, _08460_);
  nand (_13247_, _13245_, _13237_);
  nor (_13248_, _13247_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13248_, _13229_);
  and (_13249_, _08450_, word_in[19]);
  and (_13250_, _12707_, _08221_);
  and (_13251_, _12698_, _08196_);
  or (_13252_, _13251_, _13250_);
  and (_13253_, _12703_, _08208_);
  and (_13254_, _12711_, _08200_);
  or (_13255_, _13254_, _13253_);
  or (_13256_, _13255_, _13252_);
  or (_13257_, _13256_, _08419_);
  and (_13258_, _12723_, _08221_);
  and (_13259_, _12718_, _08196_);
  or (_13260_, _13259_, _13258_);
  and (_13261_, _12727_, _08208_);
  and (_13262_, _12732_, _08200_);
  or (_13263_, _13262_, _13261_);
  or (_13264_, _13263_, _13260_);
  or (_13265_, _13264_, _08460_);
  nand (_13266_, _13265_, _13257_);
  nor (_13267_, _13266_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13267_, _13249_);
  and (_13268_, _08450_, word_in[20]);
  and (_13269_, _12750_, _08221_);
  and (_13270_, _12754_, _08196_);
  or (_13271_, _13270_, _13269_);
  and (_13272_, _12746_, _08208_);
  and (_13273_, _12741_, _08200_);
  or (_13274_, _13273_, _13272_);
  or (_13275_, _13274_, _13271_);
  or (_13276_, _13275_, _08419_);
  and (_13277_, _12770_, _08221_);
  and (_13278_, _12774_, _08196_);
  or (_13279_, _13278_, _13277_);
  and (_13280_, _12766_, _08208_);
  and (_13282_, _12761_, _08200_);
  or (_13283_, _13282_, _13280_);
  or (_13284_, _13283_, _13279_);
  or (_13285_, _13284_, _08460_);
  nand (_13286_, _13285_, _13276_);
  nor (_13287_, _13286_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13287_, _13268_);
  and (_13288_, _08450_, word_in[21]);
  and (_13290_, _12793_, _08221_);
  and (_13291_, _12797_, _08196_);
  or (_13292_, _13291_, _13290_);
  and (_13293_, _12789_, _08208_);
  and (_13294_, _12784_, _08200_);
  or (_13295_, _13294_, _13293_);
  or (_13296_, _13295_, _13292_);
  or (_13297_, _13296_, _08419_);
  and (_13298_, _12817_, _08196_);
  and (_13299_, _12804_, _08200_);
  or (_13300_, _13299_, _13298_);
  and (_13301_, _12813_, _08221_);
  and (_13302_, _12809_, _08208_);
  or (_13303_, _13302_, _13301_);
  or (_13304_, _13303_, _13300_);
  or (_13305_, _13304_, _08460_);
  nand (_13306_, _13305_, _13297_);
  nor (_13307_, _13306_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13307_, _13288_);
  and (_13308_, _08450_, word_in[22]);
  and (_13309_, _12836_, _08221_);
  and (_13310_, _12840_, _08196_);
  or (_13311_, _13310_, _13309_);
  and (_13312_, _12832_, _08208_);
  and (_13313_, _12827_, _08200_);
  or (_13314_, _13313_, _13312_);
  or (_13315_, _13314_, _13311_);
  or (_13316_, _13315_, _08419_);
  and (_13317_, _12860_, _08196_);
  and (_13318_, _12847_, _08200_);
  or (_13319_, _13318_, _13317_);
  and (_13320_, _12856_, _08221_);
  and (_13321_, _12852_, _08208_);
  or (_13322_, _13321_, _13320_);
  or (_13323_, _13322_, _13319_);
  or (_13325_, _13323_, _08460_);
  nand (_13326_, _13325_, _13316_);
  nor (_13327_, _13326_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13327_, _13308_);
  or (_13329_, _11830_, _08748_);
  and (_13330_, _13329_, _11889_);
  and (_13331_, _11830_, _11395_);
  and (_13332_, _11852_, _11415_);
  or (_13333_, _13332_, _13331_);
  or (_13334_, _13333_, _13330_);
  and (_13335_, _11810_, _08750_);
  and (_13337_, _11867_, _11415_);
  or (_13338_, _13337_, _13335_);
  and (_13339_, _11737_, _11810_);
  and (_13340_, _11805_, _11415_);
  or (_13341_, _13340_, _13339_);
  or (_13342_, _13341_, _13338_);
  or (_13343_, _13342_, _13334_);
  and (_13344_, _11404_, _08757_);
  and (_13345_, _11400_, _08757_);
  or (_13346_, _13345_, _13344_);
  or (_13347_, _13346_, _12536_);
  or (_13348_, _13347_, _13343_);
  nor (_13349_, _11878_, _08715_);
  and (_13350_, _11404_, _11395_);
  and (_13351_, _11391_, _08758_);
  and (_13352_, _13351_, _08736_);
  or (_13353_, _13352_, _13350_);
  or (_13354_, _11410_, _11400_);
  and (_13355_, _13354_, _11810_);
  or (_13356_, _13355_, _13353_);
  or (_13357_, _13356_, _13349_);
  or (_13358_, _11921_, _11887_);
  and (_13360_, _11415_, _11404_);
  or (_13361_, _13360_, _12549_);
  or (_13362_, _13361_, _13358_);
  or (_13364_, _11918_, _11909_);
  or (_13365_, _13364_, _11803_);
  or (_13367_, _13365_, _13362_);
  or (_13368_, _13367_, _13357_);
  or (_13370_, _13368_, _13348_);
  and (_13372_, _13370_, _06527_);
  and (_13373_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_13375_, _08732_, _11390_);
  and (_13376_, _13375_, _08749_);
  and (_13377_, _13376_, _08754_);
  and (_13378_, _08741_, _08736_);
  and (_13379_, _13378_, _08746_);
  and (_13380_, _13379_, _08757_);
  or (_13381_, _13380_, _08767_);
  or (_13382_, _13381_, _13377_);
  not (_13383_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_13384_, _11795_, _13383_);
  and (_13385_, _13384_, _13382_);
  or (_13386_, _13385_, _13373_);
  or (_13387_, _13386_, _13372_);
  and (_11599_, _13387_, _06071_);
  and (_13389_, _08508_, word_in[24]);
  and (_13390_, _12884_, _08359_);
  and (_13391_, _12880_, _08358_);
  or (_13393_, _13391_, _13390_);
  and (_13394_, _13393_, _08482_);
  and (_13395_, _12874_, _08359_);
  and (_13396_, _12870_, _08358_);
  or (_13397_, _13396_, _13395_);
  and (_13398_, _13397_, _08480_);
  and (_13399_, _12894_, _08359_);
  and (_13400_, _12890_, _08358_);
  or (_13401_, _13400_, _13399_);
  and (_13402_, _13401_, _08517_);
  and (_13403_, _12904_, _08359_);
  and (_13404_, _12900_, _08358_);
  or (_13405_, _13404_, _13403_);
  and (_13406_, _13405_, _08522_);
  or (_13407_, _13406_, _13402_);
  or (_13408_, _13407_, _13398_);
  nor (_13409_, _13408_, _13394_);
  nor (_13410_, _13409_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13410_, _13389_);
  and (_13411_, _08508_, word_in[25]);
  and (_13412_, _12931_, _08359_);
  and (_13414_, _12927_, _08358_);
  or (_13415_, _13414_, _13412_);
  and (_13417_, _13415_, _08482_);
  and (_13418_, _12921_, _08359_);
  and (_13419_, _12916_, _08358_);
  or (_13420_, _13419_, _13418_);
  and (_13421_, _13420_, _08480_);
  and (_13422_, _12941_, _08359_);
  and (_13423_, _12937_, _08358_);
  or (_13425_, _13423_, _13422_);
  and (_13426_, _13425_, _08517_);
  and (_13428_, _12951_, _08359_);
  and (_13429_, _12947_, _08358_);
  or (_13431_, _13429_, _13428_);
  and (_13432_, _13431_, _08522_);
  or (_13434_, _13432_, _13426_);
  or (_13435_, _13434_, _13421_);
  nor (_13437_, _13435_, _13417_);
  nor (_13438_, _13437_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13438_, _13411_);
  and (_13440_, _08508_, word_in[26]);
  and (_13442_, _12966_, _08359_);
  and (_13443_, _12962_, _08358_);
  or (_13444_, _13443_, _13442_);
  and (_13445_, _13444_, _08480_);
  and (_13446_, _12976_, _08359_);
  and (_13447_, _12972_, _08358_);
  or (_13448_, _13447_, _13446_);
  and (_13449_, _13448_, _08482_);
  and (_13450_, _12986_, _08359_);
  and (_13451_, _12982_, _08358_);
  or (_13452_, _13451_, _13450_);
  and (_13453_, _13452_, _08517_);
  and (_13454_, _12996_, _08359_);
  and (_13455_, _12992_, _08358_);
  or (_13456_, _13455_, _13454_);
  and (_13458_, _13456_, _08522_);
  or (_13459_, _13458_, _13453_);
  or (_13460_, _13459_, _13449_);
  nor (_13462_, _13460_, _13445_);
  nor (_13463_, _13462_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13463_, _13440_);
  and (_13465_, _08508_, word_in[27]);
  and (_13466_, _13012_, _08359_);
  and (_13467_, _13008_, _08358_);
  or (_13468_, _13467_, _13466_);
  and (_13469_, _13468_, _08480_);
  and (_13470_, _13022_, _08359_);
  and (_13471_, _13018_, _08358_);
  or (_13472_, _13471_, _13470_);
  and (_13473_, _13472_, _08482_);
  and (_13474_, _13032_, _08359_);
  and (_13476_, _13028_, _08358_);
  or (_13477_, _13476_, _13474_);
  and (_13479_, _13477_, _08517_);
  and (_13480_, _13043_, _08359_);
  and (_13481_, _13039_, _08358_);
  or (_13482_, _13481_, _13480_);
  and (_13483_, _13482_, _08522_);
  or (_13484_, _13483_, _13479_);
  or (_13485_, _13484_, _13473_);
  nor (_13486_, _13485_, _13469_);
  nor (_13488_, _13486_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13488_, _13465_);
  and (_13489_, _08508_, word_in[28]);
  and (_13490_, _13069_, _08359_);
  and (_13491_, _13065_, _08358_);
  or (_13492_, _13491_, _13490_);
  and (_13493_, _13492_, _08482_);
  and (_13494_, _13059_, _08359_);
  and (_13495_, _13054_, _08358_);
  or (_13496_, _13495_, _13494_);
  and (_13498_, _13496_, _08480_);
  and (_13499_, _13079_, _08359_);
  and (_13500_, _13075_, _08358_);
  or (_13501_, _13500_, _13499_);
  and (_13503_, _13501_, _08517_);
  and (_13504_, _13090_, _08359_);
  and (_13506_, _13086_, _08358_);
  or (_13507_, _13506_, _13504_);
  and (_13509_, _13507_, _08522_);
  or (_13510_, _13509_, _13503_);
  or (_13511_, _13510_, _13498_);
  nor (_13512_, _13511_, _13493_);
  nor (_13513_, _13512_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13513_, _13489_);
  and (_13514_, _08508_, word_in[29]);
  and (_13515_, _13117_, _08359_);
  and (_13516_, _13113_, _08358_);
  or (_13518_, _13516_, _13515_);
  and (_13519_, _13518_, _08482_);
  and (_13521_, _13106_, _08359_);
  and (_13522_, _13102_, _08358_);
  or (_13523_, _13522_, _13521_);
  and (_13524_, _13523_, _08480_);
  and (_13525_, _13127_, _08359_);
  and (_13526_, _13123_, _08358_);
  or (_13527_, _13526_, _13525_);
  and (_13528_, _13527_, _08517_);
  and (_13529_, _13137_, _08359_);
  and (_13530_, _13133_, _08358_);
  or (_13531_, _13530_, _13529_);
  and (_13532_, _13531_, _08522_);
  or (_13533_, _13532_, _13528_);
  or (_13534_, _13533_, _13524_);
  nor (_13535_, _13534_, _13519_);
  nor (_13537_, _13535_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13537_, _13514_);
  and (_13538_, _08508_, word_in[30]);
  and (_13539_, _13162_, _08359_);
  and (_13540_, _13158_, _08358_);
  or (_13541_, _13540_, _13539_);
  and (_13543_, _13541_, _08482_);
  and (_13544_, _13152_, _08359_);
  and (_13546_, _13148_, _08358_);
  or (_13547_, _13546_, _13544_);
  and (_13549_, _13547_, _08480_);
  and (_13550_, _13172_, _08359_);
  and (_13551_, _13168_, _08358_);
  or (_13552_, _13551_, _13550_);
  and (_13553_, _13552_, _08517_);
  and (_13554_, _13182_, _08359_);
  and (_13555_, _13178_, _08358_);
  or (_13556_, _13555_, _13554_);
  and (_13557_, _13556_, _08522_);
  or (_13558_, _13557_, _13553_);
  or (_13559_, _13558_, _13549_);
  nor (_13560_, _13559_, _13543_);
  nor (_13562_, _13560_, _08508_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13562_, _13538_);
  and (_13564_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08003_);
  and (_13566_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_13567_, _13566_, _13564_);
  and (_11677_, _13567_, _06071_);
  nor (_11692_, _11627_, rst);
  nor (_11712_, _11688_, rst);
  or (_13569_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_13570_, _06530_, _05760_);
  and (_13572_, _13570_, _06071_);
  and (_11720_, _13572_, _13569_);
  nand (_13574_, _06376_, _06386_);
  or (_13576_, _09347_, _13574_);
  and (_13577_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_13578_, _07978_, _06966_);
  or (_13579_, _06391_, _06381_);
  and (_13580_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_13582_, _13580_, _13579_);
  or (_13583_, _13582_, _13578_);
  or (_13584_, _13583_, _13577_);
  and (_11767_, _13584_, _06071_);
  or (_13585_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand (_13586_, _06530_, _05862_);
  and (_13587_, _13586_, _06071_);
  and (_11809_, _13587_, _13585_);
  and (_13588_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_13589_, _12197_, _06369_);
  or (_13590_, _13589_, _13588_);
  and (_11820_, _13590_, _06071_);
  nor (_13592_, _11242_, _11240_);
  nor (_13593_, _13592_, _11243_);
  or (_13594_, _13593_, _09711_);
  or (_13595_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_13597_, _13595_, _11270_);
  and (_13598_, _13597_, _13594_);
  and (_13599_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_11832_, _13599_, _13598_);
  nor (_11871_, _11607_, rst);
  nand (_13602_, _10978_, _08053_);
  or (_13603_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_13604_, _13603_, _06071_);
  and (_11886_, _13604_, _13602_);
  and (_13606_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_13608_, _12120_, _07979_);
  or (_13609_, _13608_, _13606_);
  and (_11892_, _13609_, _06071_);
  or (_13611_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_13613_, _06530_, _05782_);
  and (_13614_, _13613_, _06071_);
  and (_11898_, _13614_, _13611_);
  and (_13616_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_13617_, _11239_, _11237_);
  nor (_13618_, _13617_, _11240_);
  or (_13619_, _13618_, _09711_);
  or (_13620_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_13621_, _13620_, _11270_);
  and (_13623_, _13621_, _13619_);
  or (_11941_, _13623_, _13616_);
  and (_13625_, _11422_, _11401_);
  and (_13627_, _11745_, _08732_);
  or (_13628_, _13627_, _13625_);
  and (_13629_, _11396_, _08748_);
  or (_13630_, _13629_, _11875_);
  and (_13631_, _11860_, _08764_);
  or (_13632_, _11408_, _11400_);
  and (_13633_, _13632_, _11395_);
  or (_13634_, _13633_, _13631_);
  or (_13635_, _13634_, _13630_);
  or (_13636_, _13635_, _13628_);
  and (_13637_, _13636_, _11421_);
  and (_13638_, _13628_, _11385_);
  and (_13639_, _13379_, _08764_);
  and (_13640_, _13639_, _11810_);
  or (_13641_, _13640_, _11811_);
  and (_13642_, _13641_, _13384_);
  or (_13643_, _13642_, _13638_);
  or (_13644_, _13643_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_13645_, _13644_, _13637_);
  or (_13646_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05686_);
  and (_13647_, _13646_, _06071_);
  and (_11988_, _13647_, _13645_);
  and (_13648_, _12161_, _06369_);
  not (_13649_, _06376_);
  or (_13650_, _06394_, _13649_);
  nor (_13651_, _06387_, _06390_);
  or (_13652_, _13651_, _13650_);
  and (_13653_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or (_13654_, _13653_, _13648_);
  and (_12012_, _13654_, _06071_);
  and (_13655_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_13656_, _11023_, _06369_);
  or (_13657_, _13656_, _13655_);
  and (_12018_, _13657_, _06071_);
  and (_13658_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_13659_, _06611_, _06434_);
  or (_13660_, _13659_, _13658_);
  and (_12048_, _13660_, _06071_);
  or (_13661_, _11254_, _11249_);
  nor (_13662_, _11255_, _09711_);
  and (_13663_, _13662_, _13661_);
  nor (_13664_, _09710_, _06153_);
  nor (_13665_, _13664_, _13663_);
  or (_13666_, _13665_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand (_13667_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_13668_, _13667_, _13666_);
  nor (_12089_, _13668_, rst);
  and (_13669_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_13670_, _11023_, _06966_);
  and (_13671_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_13672_, _13671_, _13579_);
  or (_13673_, _13672_, _13670_);
  or (_13674_, _13673_, _13669_);
  and (_12099_, _13674_, _06071_);
  and (_13675_, _13576_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_13676_, _07945_, _06967_);
  and (_13677_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_13678_, _13677_, _13579_);
  or (_13679_, _13678_, _13676_);
  or (_13680_, _13679_, _13675_);
  and (_12101_, _13680_, _06071_);
  and (_13681_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_13682_, _11260_, _11258_);
  nor (_13683_, _13682_, _11261_);
  or (_13684_, _13683_, _09711_);
  or (_13685_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_13687_, _13685_, _11270_);
  and (_13688_, _13687_, _13684_);
  or (_12111_, _13688_, _13681_);
  nor (_13689_, _11257_, _11084_);
  nor (_13690_, _13689_, _11258_);
  or (_13691_, _13690_, _09711_);
  or (_13692_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_13693_, _13692_, _11270_);
  and (_13694_, _13693_, _13691_);
  and (_13695_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_12141_, _13695_, _13694_);
  and (_12170_, _08753_, _06071_);
  and (_13696_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_13697_, _11256_, _11087_);
  nor (_13698_, _13697_, _11257_);
  or (_13699_, _13698_, _09711_);
  or (_13700_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_13701_, _13700_, _11270_);
  and (_13702_, _13701_, _13699_);
  or (_12175_, _13702_, _13696_);
  nor (_12179_, _11493_, rst);
  not (_13703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_13704_, _13703_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_13705_, _13704_, _07885_);
  nor (_13706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_13707_, _13706_, _13705_);
  or (_13708_, _13707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_13709_, _06026_, _05923_);
  and (_13710_, _13709_, _10946_);
  and (_13711_, _13710_, _06806_);
  or (_13712_, _13711_, _13708_);
  and (_13713_, _08799_, _06383_);
  or (_13714_, _06383_, _07907_);
  nand (_13715_, _13714_, _13711_);
  or (_13716_, _13715_, _13713_);
  and (_13717_, _13716_, _13712_);
  and (_13718_, _09248_, _06821_);
  or (_13719_, _13718_, _13717_);
  nand (_13720_, _13718_, _07977_);
  and (_13721_, _13720_, _06071_);
  and (_12181_, _13721_, _13719_);
  and (_13722_, _07104_, _06805_);
  and (_13723_, _13722_, _06840_);
  nand (_13724_, _13723_, _09341_);
  or (_13725_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_13726_, _13725_, _06071_);
  and (_12190_, _13726_, _13724_);
  nand (_13727_, _13723_, _09037_);
  or (_13728_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_13729_, _13728_, _06071_);
  and (_12193_, _13729_, _13727_);
  and (_13730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_13731_, _13730_, _07885_);
  and (_13732_, _07902_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_13733_, _13732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_13734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_13735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_13736_, _13735_, _13734_);
  and (_13737_, _13736_, _13733_);
  nor (_13738_, _13737_, _13731_);
  and (_13739_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  not (_13740_, _13738_);
  and (_13741_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_13742_, _13741_, _13739_);
  and (_13743_, _06380_, _06012_);
  and (_13744_, _13743_, _06821_);
  or (_13745_, _13744_, _13742_);
  not (_13746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand (_13747_, _13746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand (_13748_, _13747_, _07902_);
  nand (_13749_, _13748_, _13744_);
  and (_13750_, _13749_, _13745_);
  and (_12200_, _13750_, _06071_);
  and (_13751_, _06362_, _06027_);
  and (_13752_, _13751_, _06821_);
  and (_13753_, _13752_, _07885_);
  and (_13754_, _13753_, _12019_);
  and (_13755_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_13756_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_13757_, _13756_, _13755_);
  nor (_13758_, _13757_, _13744_);
  and (_13759_, _13752_, _07902_);
  not (_13760_, _13759_);
  nor (_13761_, _13760_, _06434_);
  or (_13762_, _13761_, _13758_);
  or (_13763_, _13762_, _13754_);
  and (_12203_, _13763_, _06071_);
  or (_13764_, _13737_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not (_13765_, _13731_);
  not (_13766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand (_13767_, _13737_, _13766_);
  and (_13769_, _13767_, _13765_);
  and (_13770_, _13769_, _13764_);
  nor (_13771_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_13772_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_13774_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_13776_, _13774_, _13772_);
  and (_13777_, _13776_, _13771_);
  not (_13778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_13779_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_13780_, _13779_, _13778_);
  and (_13781_, _13780_, _13766_);
  and (_13782_, _13781_, _13777_);
  nor (_13783_, _13782_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_13784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_13785_, _13784_, _13783_);
  and (_13786_, _13785_, _13731_);
  nor (_13788_, _13786_, _13770_);
  nor (_13789_, _13788_, _13752_);
  and (_13790_, _13753_, _07978_);
  or (_13791_, _13790_, _13789_);
  and (_12206_, _13791_, _06071_);
  and (_13792_, _13733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_13793_, _13792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_13794_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_13796_, _13794_, _13733_);
  nor (_13797_, _13796_, _13793_);
  nor (_13798_, _13752_, rst);
  and (_12211_, _13798_, _13797_);
  or (_13799_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_13800_, _06530_, _05716_);
  and (_13802_, _13800_, _06071_);
  and (_12214_, _13802_, _13799_);
  and (_13803_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_13804_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_13805_, _13804_, _13803_);
  and (_12217_, _13805_, _06071_);
  nor (_13806_, _11255_, _11091_);
  nor (_13807_, _13806_, _11256_);
  or (_13808_, _13807_, _09711_);
  or (_13809_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_13810_, _13809_, _11270_);
  and (_13811_, _13810_, _13808_);
  and (_13812_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_12220_, _13812_, _13811_);
  not (_13813_, _12167_);
  nor (_13814_, _12126_, _13813_);
  not (_13815_, _12084_);
  and (_13816_, _13815_, _12221_);
  and (_13817_, _13816_, _13814_);
  and (_13818_, _12386_, _12341_);
  not (_13819_, _12030_);
  and (_13820_, _12426_, _13819_);
  and (_13821_, _13820_, _13818_);
  and (_13822_, _13821_, _13817_);
  nor (_13823_, _12426_, _12030_);
  and (_13824_, _13823_, _13818_);
  and (_13825_, _13824_, _13817_);
  nor (_13826_, _13825_, _13822_);
  not (_13827_, _12341_);
  and (_13828_, _12386_, _13827_);
  and (_13829_, _13828_, _13823_);
  and (_13830_, _13829_, _13817_);
  nor (_13831_, _12386_, _13827_);
  and (_13832_, _13820_, _13831_);
  and (_13833_, _13832_, _13817_);
  nor (_13835_, _13833_, _13830_);
  and (_13836_, _13835_, _13826_);
  and (_13837_, _12126_, _13815_);
  and (_13838_, _12221_, _12167_);
  and (_13839_, _13838_, _13837_);
  and (_13840_, _13821_, _13839_);
  nor (_13842_, _12386_, _12341_);
  and (_13843_, _13842_, _13820_);
  and (_13844_, _13843_, _13817_);
  nor (_13845_, _13844_, _13840_);
  not (_13846_, _12221_);
  and (_13847_, _13837_, _13813_);
  and (_13848_, _13847_, _13846_);
  not (_13849_, _12426_);
  and (_13850_, _13842_, _13849_);
  and (_13851_, _13850_, _12030_);
  and (_13852_, _13851_, _13848_);
  and (_13853_, _13847_, _12221_);
  and (_13854_, _13853_, _13821_);
  nor (_13856_, _13854_, _13852_);
  and (_13857_, _13856_, _13845_);
  and (_13858_, _13857_, _13836_);
  and (_13860_, _13843_, _13839_);
  and (_13861_, _13828_, _13820_);
  and (_13863_, _13861_, _13839_);
  nor (_13864_, _13863_, _13860_);
  and (_13865_, _13832_, _13839_);
  and (_13866_, _13829_, _13839_);
  nor (_13867_, _13866_, _13865_);
  and (_13869_, _13867_, _13864_);
  and (_13870_, _13824_, _13839_);
  and (_13871_, _13851_, _13839_);
  nor (_13872_, _13871_, _13870_);
  nor (_13873_, _12221_, _13813_);
  and (_13874_, _13873_, _13837_);
  and (_13875_, _13874_, _13821_);
  and (_13876_, _13861_, _13874_);
  nor (_13877_, _13876_, _13875_);
  and (_13878_, _13877_, _13872_);
  and (_13879_, _13878_, _13869_);
  and (_13880_, _13879_, _13858_);
  and (_13881_, _12426_, _12030_);
  and (_13882_, _13818_, _13881_);
  nor (_13883_, _12084_, _12221_);
  and (_13884_, _13883_, _13814_);
  and (_13885_, _13884_, _13882_);
  and (_13886_, _13882_, _12221_);
  nor (_13887_, _12126_, _12167_);
  and (_13888_, _13887_, _13815_);
  and (_13889_, _13888_, _13886_);
  nor (_13890_, _13889_, _13885_);
  nand (_13891_, _13882_, _13837_);
  and (_13892_, _13881_, _13839_);
  and (_13893_, _13892_, _13831_);
  and (_13894_, _13842_, _13881_);
  and (_13895_, _13894_, _13839_);
  nor (_13896_, _13895_, _13893_);
  and (_13897_, _13828_, _13892_);
  and (_13898_, _13882_, _13846_);
  and (_13899_, _13888_, _13898_);
  nor (_13900_, _13899_, _13897_);
  and (_13901_, _13900_, _13896_);
  and (_13902_, _13901_, _13891_);
  and (_13903_, _13902_, _13890_);
  and (_13904_, _13903_, _13880_);
  and (_13905_, _13889_, _07823_);
  not (_13906_, _12295_);
  and (_13907_, _13885_, _13906_);
  nor (_13908_, _13907_, _13905_);
  nand (_13909_, _13895_, _07429_);
  and (_13910_, _13909_, _13908_);
  nor (_13911_, _13910_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_13912_, _13911_);
  and (_13913_, _13889_, _07766_);
  not (_13914_, _10946_);
  nor (_13915_, _13850_, _13914_);
  and (_13916_, _13915_, _12228_);
  nor (_13917_, _13916_, _13913_);
  and (_13918_, _13917_, _12435_);
  and (_13919_, _13918_, _13912_);
  not (_13920_, _13919_);
  nor (_13921_, _13920_, _13904_);
  not (_13922_, _13921_);
  and (_13923_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_13924_, _13893_, _07429_);
  not (_13925_, _13924_);
  nand (_13926_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand (_13927_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_13928_, _13927_, _13926_);
  nand (_13929_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_13930_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_13931_, _13930_, _13929_);
  and (_13932_, _13931_, _13928_);
  nand (_13933_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_13934_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_13935_, _13934_, _13933_);
  nand (_13936_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand (_13937_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_13938_, _13937_, _13936_);
  and (_13939_, _13938_, _13935_);
  and (_13940_, _13939_, _13932_);
  nand (_13942_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_13943_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_13944_, _13943_, _13942_);
  nand (_13945_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand (_13946_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_13947_, _13946_, _13945_);
  and (_13948_, _13947_, _13944_);
  nand (_13949_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand (_13950_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_13951_, _13950_, _13949_);
  nand (_13952_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_13953_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_13954_, _13953_, _13952_);
  and (_13955_, _13954_, _13951_);
  and (_13956_, _13955_, _13948_);
  and (_13957_, _13956_, _13940_);
  nand (_13958_, _13897_, _11961_);
  nand (_13959_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_13960_, _13959_, _13958_);
  nand (_13961_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand (_13962_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_13963_, _13962_, _13961_);
  and (_13964_, _13963_, _13960_);
  and (_13966_, _13898_, _13847_);
  and (_13967_, _11399_, _11390_);
  and (_13968_, _13967_, _08746_);
  nor (_13969_, _13968_, _11918_);
  nor (_13970_, _11885_, _11739_);
  nor (_13971_, _13331_, _12541_);
  and (_13972_, _13971_, _13970_);
  and (_13973_, _13972_, _13969_);
  and (_13974_, _13973_, _11866_);
  not (_13975_, _11855_);
  and (_13976_, _11400_, _11395_);
  nor (_13977_, _13976_, _13975_);
  not (_13978_, _11870_);
  nor (_13979_, _13337_, _13978_);
  and (_13980_, _13979_, _13977_);
  and (_13981_, _13980_, _13974_);
  and (_13982_, _13981_, _11851_);
  nor (_13983_, _13982_, _11744_);
  nor (_13985_, _13983_, p3_in[3]);
  not (_13986_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_13987_, _13983_, _13986_);
  nor (_13988_, _13987_, _13985_);
  nand (_13990_, _13988_, _13966_);
  and (_13991_, _13853_, _13882_);
  nor (_13993_, _13983_, p2_in[3]);
  not (_13994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_13996_, _13983_, _13994_);
  nor (_13997_, _13996_, _13993_);
  nand (_13998_, _13997_, _13991_);
  and (_13999_, _13998_, _13990_);
  and (_14000_, _13882_, _13839_);
  nor (_14002_, _13983_, p0_in[3]);
  not (_14003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_14004_, _13983_, _14003_);
  nor (_14005_, _14004_, _14002_);
  nand (_14006_, _14005_, _14000_);
  and (_14007_, _13874_, _13882_);
  nor (_00002_, _13983_, p1_in[3]);
  not (_00003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00004_, _13983_, _00003_);
  nor (_00005_, _00004_, _00002_);
  nand (_00006_, _00005_, _14007_);
  and (_00007_, _00006_, _14006_);
  and (_00008_, _00007_, _13999_);
  and (_00009_, _00008_, _13964_);
  nand (_00010_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_00011_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00012_, _00011_, _00010_);
  and (_00013_, _00012_, _00009_);
  nand (_00015_, _00013_, _13957_);
  nand (_00016_, _00015_, _13919_);
  nand (_00017_, _00016_, _13925_);
  or (_00018_, _00017_, _13923_);
  nand (_00019_, _13924_, _11791_);
  and (_00020_, _00019_, _06071_);
  and (_12226_, _00020_, _00018_);
  and (_00021_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00022_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_00023_, _00022_, _00021_);
  and (_12229_, _00023_, _06071_);
  and (_00024_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_00025_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_00026_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_00027_, _00026_, _00025_);
  and (_00028_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_00029_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_00030_, _00029_, _00028_);
  or (_00031_, _00030_, _00027_);
  and (_00032_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_00033_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_00034_, _00033_, _00032_);
  and (_00035_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_00036_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00037_, _00036_, _00035_);
  or (_00038_, _00037_, _00034_);
  or (_00039_, _00038_, _00031_);
  and (_00040_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00041_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_00042_, _00041_, _00040_);
  and (_00043_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00044_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00045_, _00044_, _00043_);
  or (_00046_, _00045_, _00042_);
  and (_00047_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_00048_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_00049_, _00048_, _00047_);
  and (_00050_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00051_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_00052_, _00051_, _00050_);
  or (_00053_, _00052_, _00049_);
  or (_00054_, _00053_, _00046_);
  or (_00055_, _00054_, _00039_);
  and (_00056_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00057_, _13897_, _12398_);
  or (_00058_, _00057_, _00056_);
  and (_00059_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00060_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00061_, _00060_, _00059_);
  or (_00062_, _00061_, _00058_);
  or (_00063_, _13983_, p0_in[2]);
  not (_00064_, _13983_);
  or (_00065_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_00066_, _00065_, _00063_);
  and (_00067_, _00066_, _14000_);
  or (_00068_, _13983_, p1_in[2]);
  or (_00069_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_00070_, _00069_, _00068_);
  and (_00071_, _00070_, _14007_);
  or (_00072_, _00071_, _00067_);
  or (_00073_, _13983_, p3_in[2]);
  or (_00074_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_00075_, _00074_, _00073_);
  and (_00076_, _00075_, _13966_);
  or (_00077_, _13983_, p2_in[2]);
  or (_00078_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_00079_, _00078_, _00077_);
  and (_00080_, _00079_, _13991_);
  or (_00081_, _00080_, _00076_);
  or (_00082_, _00081_, _00072_);
  or (_00083_, _00082_, _00062_);
  and (_00084_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00085_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_00086_, _00085_, _00084_);
  or (_00087_, _00086_, _00083_);
  or (_00088_, _00087_, _00055_);
  and (_00089_, _00088_, _13919_);
  or (_00090_, _00089_, _13924_);
  or (_00091_, _00090_, _00024_);
  or (_00092_, _13925_, _07564_);
  and (_00093_, _00092_, _06071_);
  and (_12232_, _00093_, _00091_);
  and (_00094_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_00095_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_00096_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_00097_, _00096_, _00095_);
  and (_00098_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_00099_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_00100_, _00099_, _00098_);
  or (_00101_, _00100_, _00097_);
  and (_00102_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_00103_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_00104_, _00103_, _00102_);
  and (_00105_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00106_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_00107_, _00106_, _00105_);
  or (_00108_, _00107_, _00104_);
  or (_00109_, _00108_, _00101_);
  and (_00110_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00111_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00112_, _00111_, _00110_);
  and (_00113_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00114_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00115_, _00114_, _00113_);
  or (_00116_, _00115_, _00112_);
  and (_00117_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_00118_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_00119_, _00118_, _00117_);
  and (_00120_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00121_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_00122_, _00121_, _00120_);
  or (_00123_, _00122_, _00119_);
  or (_00124_, _00123_, _00116_);
  or (_00125_, _00124_, _00109_);
  and (_00126_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00127_, _13897_, _12379_);
  or (_00128_, _00127_, _00126_);
  and (_00129_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00130_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00131_, _00130_, _00129_);
  or (_00132_, _00131_, _00128_);
  or (_00133_, _13983_, p0_in[1]);
  or (_00134_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_00135_, _00134_, _00133_);
  and (_00136_, _00135_, _14000_);
  or (_00137_, _13983_, p1_in[1]);
  or (_00138_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_00139_, _00138_, _00137_);
  and (_00140_, _00139_, _14007_);
  or (_00141_, _00140_, _00136_);
  or (_00142_, _13983_, p2_in[1]);
  or (_00143_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_00144_, _00143_, _00142_);
  and (_00145_, _00144_, _13991_);
  or (_00146_, _13983_, p3_in[1]);
  or (_00147_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_00148_, _00147_, _00146_);
  and (_00149_, _00148_, _13966_);
  or (_00150_, _00149_, _00145_);
  or (_00151_, _00150_, _00141_);
  or (_00152_, _00151_, _00132_);
  and (_00153_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00154_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_00155_, _00154_, _00153_);
  or (_00156_, _00155_, _00152_);
  or (_00157_, _00156_, _00125_);
  and (_00158_, _00157_, _13919_);
  or (_00159_, _00158_, _13924_);
  or (_00160_, _00159_, _00094_);
  nand (_00161_, _13924_, _08110_);
  and (_00162_, _00161_, _06071_);
  and (_12235_, _00162_, _00160_);
  or (_00163_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_00164_, _06530_, _05749_);
  and (_00165_, _00164_, _06071_);
  and (_12254_, _00165_, _00163_);
  or (_00166_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  nand (_00167_, _06530_, _11276_);
  and (_00168_, _00167_, _06071_);
  and (_12261_, _00168_, _00166_);
  nand (_00169_, _13924_, _08053_);
  and (_00170_, _00169_, _06071_);
  nand (_00171_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_00172_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_00173_, _00172_, _00171_);
  nand (_00174_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_00175_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_00176_, _00175_, _00174_);
  and (_00177_, _00176_, _00173_);
  nand (_00178_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_00179_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_00180_, _00179_, _00178_);
  nand (_00181_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_00182_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00183_, _00182_, _00181_);
  and (_00184_, _00183_, _00180_);
  and (_00185_, _00184_, _00177_);
  nand (_00187_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_00188_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00189_, _00188_, _00187_);
  nand (_00190_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_00191_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00192_, _00191_, _00190_);
  and (_00193_, _00192_, _00189_);
  nand (_00194_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_00195_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_00196_, _00195_, _00194_);
  nand (_00197_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00198_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_00199_, _00198_, _00197_);
  and (_00200_, _00199_, _00196_);
  and (_00201_, _00200_, _00193_);
  and (_00202_, _00201_, _00185_);
  nand (_00203_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_00204_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00205_, _00204_, _00203_);
  nand (_00206_, _13897_, _12337_);
  nand (_00207_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00208_, _00207_, _00206_);
  and (_00209_, _00208_, _00205_);
  nor (_00210_, _13983_, p2_in[0]);
  not (_00211_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_00212_, _13983_, _00211_);
  nor (_00213_, _00212_, _00210_);
  nand (_00214_, _00213_, _13991_);
  nor (_00215_, _13983_, p3_in[0]);
  not (_00216_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_00217_, _13983_, _00216_);
  nor (_00218_, _00217_, _00215_);
  nand (_00219_, _00218_, _13966_);
  and (_00220_, _00219_, _00214_);
  nor (_00221_, _13983_, p0_in[0]);
  not (_00222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_00223_, _13983_, _00222_);
  nor (_00224_, _00223_, _00221_);
  nand (_00225_, _00224_, _14000_);
  nor (_00226_, _13983_, p1_in[0]);
  not (_00227_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_00228_, _13983_, _00227_);
  nor (_00229_, _00228_, _00226_);
  nand (_00230_, _00229_, _14007_);
  and (_00231_, _00230_, _00225_);
  and (_00232_, _00231_, _00220_);
  and (_00233_, _00232_, _00209_);
  nand (_00234_, _08811_, _07872_);
  or (_00235_, _08811_, _07872_);
  nand (_00236_, _00235_, _00234_);
  or (_00237_, _07772_, _07715_);
  and (_00238_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_00239_, _06006_, _06161_);
  nor (_00240_, _00239_, _10928_);
  nor (_00241_, _00240_, _08806_);
  nor (_00242_, _00241_, _00238_);
  and (_00243_, _00242_, _07830_);
  nand (_00244_, _00243_, _00237_);
  and (_00245_, _07823_, _07746_);
  not (_00246_, _00245_);
  and (_00247_, _00246_, _00244_);
  or (_00248_, _00247_, _08952_);
  nand (_00249_, _00247_, _08952_);
  and (_00250_, _00249_, _00248_);
  nand (_00251_, _00250_, _00236_);
  or (_00252_, _00250_, _00236_);
  nand (_00253_, _00252_, _00251_);
  or (_00254_, _08110_, _07772_);
  and (_00255_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not (_00256_, _06362_);
  nor (_00257_, _06803_, _00256_);
  nor (_00259_, _06362_, _06226_);
  nor (_00260_, _00259_, _00257_);
  nor (_00261_, _00260_, _08806_);
  nor (_00262_, _00261_, _00255_);
  and (_00263_, _00262_, _07830_);
  nand (_00265_, _00263_, _00254_);
  and (_00266_, _08169_, _07823_);
  not (_00267_, _00266_);
  and (_00268_, _00267_, _00265_);
  or (_00269_, _00268_, _08964_);
  nand (_00270_, _00268_, _08964_);
  nand (_00271_, _00270_, _00269_);
  and (_00272_, _07773_, _07564_);
  and (_00273_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_00274_, _07754_);
  nor (_00275_, _00274_, _06803_);
  nor (_00276_, _07754_, _06237_);
  or (_00277_, _00276_, _00275_);
  and (_00278_, _00277_, _08805_);
  or (_00279_, _00278_, _00273_);
  or (_00280_, _00279_, _07823_);
  or (_00281_, _00280_, _00272_);
  or (_00282_, _07830_, _07594_);
  and (_00283_, _00282_, _00281_);
  or (_00284_, _11791_, _07772_);
  and (_00285_, _08941_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00286_, _07105_, _08799_);
  nor (_00287_, _07105_, _06183_);
  nor (_00288_, _00287_, _00286_);
  nor (_00289_, _00288_, _08806_);
  nor (_00290_, _00289_, _00285_);
  and (_00291_, _00290_, _07830_);
  and (_00292_, _00291_, _00284_);
  and (_00293_, _12466_, _07823_);
  or (_00294_, _00293_, _00292_);
  nand (_00295_, _00294_, _00283_);
  or (_00296_, _00294_, _00283_);
  and (_00297_, _00296_, _00295_);
  nand (_00298_, _00297_, _00271_);
  or (_00299_, _00297_, _00271_);
  nand (_00300_, _00299_, _00298_);
  nand (_00301_, _00300_, _00253_);
  or (_00302_, _00300_, _00253_);
  nand (_00303_, _00302_, _00301_);
  nand (_00304_, _00303_, _13885_);
  nand (_00305_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00306_, _00305_, _00304_);
  and (_00307_, _00306_, _00233_);
  and (_00308_, _00307_, _00202_);
  nor (_00309_, _00308_, _13920_);
  nand (_00310_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_00311_, _00310_, _13925_);
  or (_00312_, _00311_, _00309_);
  and (_12265_, _00312_, _00170_);
  nor (_12281_, _12323_, rst);
  nor (_12287_, _12122_, rst);
  nor (_12290_, _11511_, rst);
  nor (_00313_, _11248_, _11095_);
  nor (_00314_, _00313_, _11249_);
  or (_00315_, _00314_, _09711_);
  or (_00317_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00318_, _00317_, _11270_);
  and (_00319_, _00318_, _00315_);
  and (_00320_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_12293_, _00320_, _00319_);
  nor (_12300_, _11570_, rst);
  or (_00322_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_00323_, _00322_, _13711_);
  nand (_00324_, _00256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_00325_, _00324_, _13711_);
  or (_00326_, _00325_, _00257_);
  and (_00327_, _00326_, _00323_);
  or (_00328_, _00327_, _13718_);
  nand (_00329_, _13718_, _09037_);
  and (_00330_, _00329_, _06071_);
  and (_12303_, _00330_, _00328_);
  nand (_00331_, _13723_, _06434_);
  or (_00332_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_00333_, _00332_, _06071_);
  and (_12315_, _00333_, _00331_);
  nor (_00334_, _11723_, _11471_);
  nor (_00335_, _11718_, _11472_);
  or (_00336_, _00335_, _00334_);
  nand (_00337_, _00336_, _06243_);
  or (_00338_, _00336_, _06243_);
  and (_00339_, _00338_, _00337_);
  and (_00340_, _00339_, _11751_);
  and (_00341_, _11827_, _07564_);
  and (_00342_, _11748_, _07594_);
  and (_00343_, _11628_, _11424_);
  and (_00344_, _12469_, _05768_);
  and (_00345_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_00346_, _00345_, _00344_);
  or (_00347_, _00346_, _00343_);
  nor (_00348_, _00347_, _00342_);
  nand (_00349_, _00348_, _12437_);
  or (_00350_, _00349_, _00341_);
  or (_00351_, _00350_, _00340_);
  and (_00352_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00353_, _00352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00354_, _00353_, _12503_);
  or (_00355_, _00354_, _12437_);
  and (_00356_, _00355_, _06071_);
  and (_12327_, _00356_, _00351_);
  and (_00357_, _13753_, _12197_);
  and (_00358_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_00360_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_00361_, _00360_, _00358_);
  nor (_00362_, _00361_, _13744_);
  nor (_00363_, _13760_, _07945_);
  or (_00364_, _00363_, _00362_);
  or (_00365_, _00364_, _00357_);
  and (_12331_, _00365_, _06071_);
  not (_00366_, _07643_);
  or (_00367_, _12485_, _11748_);
  and (_00368_, _00367_, _00366_);
  nor (_00369_, _11428_, _11053_);
  and (_00370_, _12469_, _12131_);
  nor (_00371_, _11533_, _11425_);
  or (_00372_, _00371_, _00370_);
  or (_00373_, _00372_, _00369_);
  not (_00374_, _11709_);
  or (_00375_, _11552_, _11553_);
  or (_00376_, _00375_, _00374_);
  nand (_00377_, _00375_, _00374_);
  and (_00378_, _00377_, _11751_);
  and (_00379_, _00378_, _00376_);
  or (_00380_, _00379_, _00373_);
  nor (_00381_, _00380_, _00368_);
  nand (_00382_, _00381_, _12437_);
  and (_00383_, _11250_, _08178_);
  and (_00384_, _00383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00385_, _00383_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00386_, _00385_, _00384_);
  or (_00387_, _00386_, _12437_);
  and (_00389_, _00387_, _06071_);
  and (_12334_, _00389_, _00382_);
  nor (_00390_, _11261_, _11079_);
  nor (_00391_, _00390_, _11262_);
  or (_00392_, _00391_, _09711_);
  or (_00394_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00395_, _00394_, _11270_);
  and (_00396_, _00395_, _00392_);
  and (_00397_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_12342_, _00397_, _00396_);
  nor (_00398_, _11247_, _11245_);
  nor (_00399_, _00398_, _11248_);
  or (_00400_, _00399_, _09711_);
  or (_00401_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00402_, _00401_, _11270_);
  and (_00403_, _00402_, _00400_);
  and (_00404_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_12345_, _00404_, _00403_);
  nor (_00405_, _11236_, _06528_);
  nand (_00406_, _00405_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00407_, _00405_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00408_, _00407_, _11270_);
  and (_12358_, _00408_, _00406_);
  and (_00409_, _07011_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00410_, _00409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12361_, _00410_, _06071_);
  nor (_12367_, _11648_, rst);
  nor (_00411_, _13796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_00412_, _13796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_00413_, _00412_, _00411_);
  and (_12373_, _00413_, _13798_);
  and (_00414_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _08003_);
  and (_00415_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00416_, _00415_, _00414_);
  and (_12392_, _00416_, _06071_);
  or (_00417_, _08992_, rxd_i);
  nand (_00418_, _00417_, _07903_);
  or (_00419_, _07904_, _07889_);
  and (_00420_, _00419_, _00418_);
  not (_00421_, _07886_);
  nand (_00422_, _07910_, _00421_);
  or (_00423_, _00422_, _00420_);
  and (_12396_, _00423_, _06560_);
  not (_00424_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_00425_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_00426_, _00425_, _00424_);
  and (_00427_, _00426_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_00428_, _00425_, _00424_);
  or (_00429_, _00428_, _00426_);
  nand (_00431_, _00429_, _06071_);
  nor (_12415_, _00431_, _00427_);
  or (_00432_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_00434_, _00425_, rst);
  and (_12440_, _00434_, _00432_);
  nor (_12448_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  not (_00435_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_00436_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_00437_, _07885_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00438_, _00437_, _00436_);
  nor (_00439_, _00438_, _00435_);
  and (_00440_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_00441_, _00440_, _00439_);
  or (_00442_, _00441_, _13711_);
  or (_00443_, _07754_, _00435_);
  nand (_00444_, _00443_, _13711_);
  or (_00445_, _00444_, _00275_);
  and (_00446_, _00445_, _00442_);
  or (_00447_, _00446_, _13718_);
  nand (_00448_, _13718_, _06434_);
  and (_00449_, _00448_, _06071_);
  and (_12461_, _00449_, _00447_);
  nand (_00450_, _13723_, _07945_);
  or (_00451_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_00452_, _00451_, _06071_);
  and (_12468_, _00452_, _00450_);
  and (_00453_, _13753_, _12161_);
  and (_00454_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_00455_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_00456_, _00455_, _00454_);
  nor (_00457_, _00456_, _13744_);
  nor (_00458_, _13760_, _06993_);
  or (_00459_, _00458_, _00457_);
  or (_00460_, _00459_, _00453_);
  and (_12471_, _00460_, _06071_);
  or (_00461_, _11719_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_00462_, _00461_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_00463_, _00462_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_00464_, _00463_, _11471_);
  and (_00465_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00466_, _00465_, _11722_);
  and (_00467_, _00466_, _11716_);
  and (_00468_, _00467_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_00469_, _00468_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_00471_, _00469_, _11472_);
  and (_00472_, _00471_, _00464_);
  nor (_00473_, _00472_, _06261_);
  and (_00474_, _00472_, _06261_);
  or (_00476_, _00474_, _00473_);
  and (_00477_, _00476_, _11751_);
  and (_00478_, _11827_, _07425_);
  and (_00479_, _11748_, _07520_);
  and (_00480_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00481_, _00480_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00482_, _00481_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_00483_, _00481_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_00484_, _00483_, _00482_);
  and (_00485_, _00484_, _12469_);
  and (_00486_, _12090_, _11424_);
  and (_00487_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_00488_, _00487_, _00486_);
  or (_00489_, _00488_, _00485_);
  or (_00490_, _00489_, _00479_);
  nor (_00491_, _00490_, _00478_);
  nand (_00492_, _00491_, _12437_);
  or (_00493_, _00492_, _00477_);
  and (_00494_, _00352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00495_, _00494_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00496_, _00495_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_00497_, _00496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00498_, _00497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_00499_, _00497_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00500_, _00499_, _00498_);
  or (_00501_, _00500_, _12437_);
  and (_00502_, _00501_, _06071_);
  and (_12490_, _00502_, _00493_);
  and (_00504_, _00462_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_00505_, _00504_, _00464_);
  or (_00506_, _00468_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00507_, _00506_, _00469_);
  or (_00508_, _00507_, _11471_);
  and (_00509_, _00508_, _11751_);
  and (_00510_, _00509_, _00505_);
  nor (_00511_, _11428_, _07643_);
  nor (_00512_, _12438_, _07673_);
  nor (_00513_, _00480_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00514_, _00513_, _00481_);
  and (_00515_, _00514_, _12469_);
  and (_00516_, _12131_, _11424_);
  or (_00517_, _00516_, _00515_);
  and (_00518_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_00519_, _00518_, _00517_);
  nor (_00520_, _00519_, _00512_);
  nand (_00521_, _00520_, _12437_);
  or (_00522_, _00521_, _00511_);
  or (_00523_, _00522_, _00510_);
  nor (_00524_, _00496_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00525_, _00524_, _00497_);
  or (_00526_, _00525_, _12437_);
  and (_00527_, _00526_, _06071_);
  and (_12496_, _00527_, _00523_);
  and (_00528_, _00467_, _11472_);
  nor (_00529_, _11721_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00530_, _00529_, _00528_);
  nand (_00532_, _00530_, _06151_);
  or (_00533_, _00530_, _06151_);
  and (_00534_, _00533_, _00532_);
  and (_00535_, _00534_, _11751_);
  nor (_00536_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00537_, _00536_, _00480_);
  and (_00538_, _00537_, _12469_);
  nor (_00539_, _11428_, _07715_);
  nor (_00540_, _12438_, _07746_);
  and (_00541_, _11424_, _12172_);
  and (_00542_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_00543_, _00542_, _00541_);
  or (_00544_, _00543_, _00540_);
  or (_00545_, _00544_, _00539_);
  nor (_00546_, _00545_, _00538_);
  nand (_00547_, _00546_, _12437_);
  or (_00548_, _00547_, _00535_);
  nor (_00549_, _12505_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00550_, _00549_, _00496_);
  or (_00551_, _00550_, _12437_);
  and (_00552_, _00551_, _06071_);
  and (_12526_, _00552_, _00548_);
  nor (_00553_, _07881_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_00554_, _00553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_00555_, _00553_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_00556_, _00555_, _06071_);
  and (_12554_, _00556_, _00554_);
  not (_00557_, _13718_);
  and (_00558_, _13711_, _07105_);
  and (_00559_, _00558_, _06803_);
  nor (_00560_, _00558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_00561_, _00560_, _00559_);
  nand (_00562_, _00561_, _00557_);
  nand (_00564_, _13718_, _07945_);
  and (_00565_, _00564_, _06071_);
  and (_12557_, _00565_, _00562_);
  and (_00566_, _13753_, _12120_);
  and (_00567_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_00568_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_00569_, _00568_, _00567_);
  nor (_00570_, _00569_, _13744_);
  nor (_00571_, _13760_, _06609_);
  or (_00573_, _00571_, _00570_);
  or (_00575_, _00573_, _00566_);
  and (_12560_, _00575_, _06071_);
  not (_00576_, _13711_);
  or (_00577_, _00576_, _10936_);
  and (_00578_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_00579_, _00578_, _13718_);
  nor (_00580_, _10930_, _08993_);
  or (_00581_, _00580_, _10928_);
  and (_00582_, _00581_, _13711_);
  or (_00583_, _00582_, _00579_);
  nand (_00584_, _13718_, _06993_);
  and (_00585_, _00584_, _06071_);
  and (_12600_, _00585_, _00583_);
  nor (_00586_, _09341_, _06611_);
  and (_00587_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_00588_, _00587_, _00586_);
  and (_12624_, _00588_, _06071_);
  nand (_00589_, _11791_, _10978_);
  or (_00590_, _10978_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00591_, _00590_, _06071_);
  and (_12694_, _00591_, _00589_);
  nor (_12907_, _11931_, rst);
  not (_00593_, _07715_);
  and (_00594_, _00367_, _00593_);
  or (_00595_, _11707_, _11705_);
  and (_00596_, _11751_, _11708_);
  and (_00597_, _00596_, _00595_);
  and (_00598_, _12469_, _12172_);
  nor (_00599_, _11570_, _11425_);
  and (_00600_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00601_, _00600_, _00599_);
  or (_00602_, _00601_, _00598_);
  or (_00603_, _00602_, _00597_);
  nor (_00604_, _00603_, _00594_);
  nand (_00605_, _00604_, _12437_);
  nor (_00606_, _08180_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00607_, _00606_, _00383_);
  or (_00608_, _00607_, _12437_);
  and (_00609_, _00608_, _06071_);
  and (_13034_, _00609_, _00605_);
  or (_00610_, _12437_, _08181_);
  and (_00611_, _00610_, _06071_);
  not (_00612_, _11791_);
  and (_00613_, _00367_, _00612_);
  or (_00614_, _11610_, _11611_);
  not (_00615_, _00614_);
  nand (_00616_, _00615_, _11703_);
  or (_00617_, _00615_, _11703_);
  and (_00619_, _00617_, _11751_);
  and (_00620_, _00619_, _00616_);
  nor (_00622_, _11591_, _11425_);
  and (_00623_, _12469_, _12024_);
  or (_00624_, _00623_, _00622_);
  or (_00625_, _00624_, _00620_);
  or (_00626_, _00625_, _00613_);
  nand (_00627_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_00628_, _00627_, _12437_);
  or (_00629_, _00628_, _00626_);
  and (_13056_, _00629_, _00611_);
  or (_00630_, _12437_, _08192_);
  and (_00631_, _00630_, _06071_);
  and (_00632_, _00367_, _07564_);
  or (_00633_, _11700_, _11698_);
  and (_00634_, _11751_, _11702_);
  and (_00635_, _00634_, _00633_);
  nor (_00636_, _11428_, _08177_);
  and (_00637_, _11424_, _11612_);
  and (_00638_, _12469_, _11628_);
  or (_00639_, _00638_, _00637_);
  or (_00640_, _00639_, _00636_);
  or (_00642_, _00640_, _00635_);
  nor (_00643_, _00642_, _00632_);
  nand (_00644_, _00643_, _12437_);
  and (_13085_, _00644_, _00631_);
  not (_00645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00646_, _12437_, _11428_);
  nor (_00647_, _00646_, _00645_);
  and (_00648_, _11649_, _11424_);
  and (_00649_, _12469_, _11651_);
  or (_00650_, _00649_, _00648_);
  or (_00651_, _11695_, _11693_);
  and (_00652_, _11751_, _11697_);
  and (_00653_, _00652_, _00651_);
  or (_00654_, _00653_, _00650_);
  not (_00655_, _08110_);
  and (_00656_, _00367_, _00655_);
  or (_00657_, _00656_, _00654_);
  and (_00658_, _00657_, _12437_);
  or (_00659_, _00658_, _00647_);
  and (_13098_, _00659_, _06071_);
  not (_00660_, _08053_);
  and (_00661_, _00367_, _00660_);
  or (_00662_, _11691_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_00663_, _11693_);
  and (_00664_, _11751_, _00663_);
  and (_00665_, _00664_, _00662_);
  and (_00666_, _11827_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00667_, _11672_, _11424_);
  and (_00668_, _12469_, _11689_);
  or (_00669_, _00668_, _00667_);
  or (_00670_, _00669_, _00666_);
  or (_00671_, _00670_, _00665_);
  nor (_00672_, _00671_, _00661_);
  nand (_00673_, _00672_, _12437_);
  or (_00674_, _12437_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00675_, _00674_, _06071_);
  and (_13110_, _00675_, _00673_);
  or (_00676_, _07819_, _07757_);
  or (_00677_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00678_, _00677_, _06071_);
  and (_13206_, _00678_, _00676_);
  and (_00679_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_00680_, _07819_, _07530_);
  or (_00681_, _00680_, _00679_);
  or (_00682_, _00681_, _07429_);
  or (_00683_, _07870_, _07433_);
  and (_00684_, _00683_, _06071_);
  and (_13246_, _00684_, _00682_);
  and (_00685_, _00367_, _07425_);
  or (_00686_, _11711_, _11516_);
  and (_00687_, _11751_, _11713_);
  and (_00688_, _00687_, _00686_);
  nor (_00689_, _11428_, _11052_);
  and (_00690_, _12469_, _12090_);
  nor (_00691_, _11493_, _11425_);
  or (_00692_, _00691_, _00690_);
  or (_00693_, _00692_, _00689_);
  or (_00694_, _00693_, _00688_);
  nor (_00695_, _00694_, _00685_);
  nand (_00696_, _00695_, _12437_);
  and (_00697_, _00384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00698_, _00384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, _12437_);
  and (_00701_, _00700_, _06071_);
  and (_13281_, _00701_, _00696_);
  and (_00702_, _11716_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_00703_, _00702_, _11471_);
  and (_00704_, _11717_, _11471_);
  nor (_00705_, _00704_, _00703_);
  and (_00706_, _00705_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_00707_, _00705_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_00708_, _00707_, _11751_);
  nor (_00709_, _00708_, _00706_);
  nor (_00710_, _11428_, _08110_);
  nor (_00711_, _12438_, _08169_);
  and (_00712_, _11424_, _11651_);
  and (_00713_, _12469_, _05747_);
  or (_00714_, _00713_, _00712_);
  and (_00715_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00716_, _00715_, _00714_);
  or (_00717_, _00716_, _00711_);
  nor (_00718_, _00717_, _00710_);
  nand (_00719_, _00718_, _12437_);
  or (_00720_, _00719_, _00709_);
  nor (_00721_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_00722_, _00721_, _00352_);
  or (_00723_, _00722_, _12437_);
  and (_00724_, _00723_, _06071_);
  and (_13289_, _00724_, _00720_);
  and (_00726_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_00727_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00729_, _00727_, _06510_);
  or (_00730_, _06486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_00731_, _06499_, _06445_);
  and (_00732_, _00731_, _00730_);
  or (_00733_, _00732_, _06474_);
  and (_00734_, _00733_, _00729_);
  or (_00735_, _00734_, _00726_);
  and (_00736_, _06505_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00737_, _00736_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_00738_, _00737_, _06071_);
  and (_13324_, _00738_, _00735_);
  nor (_00739_, _11428_, _08053_);
  nand (_00740_, _11716_, _06193_);
  or (_00741_, _11716_, _06193_);
  and (_00742_, _00741_, _00740_);
  and (_00743_, _00742_, _11471_);
  and (_00744_, _00703_, _11717_);
  or (_00745_, _00744_, _00743_);
  and (_00746_, _00745_, _11751_);
  and (_00747_, _11748_, _08139_);
  and (_00748_, _12469_, _05726_);
  and (_00749_, _11689_, _11424_);
  and (_00750_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00751_, _00750_, _00749_);
  nor (_00752_, _00751_, _00748_);
  nand (_00753_, _00752_, _12437_);
  or (_00754_, _00753_, _00747_);
  or (_00755_, _00754_, _00746_);
  or (_00756_, _00755_, _00739_);
  nor (_00757_, _12500_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00758_, _00757_, _12501_);
  or (_00759_, _00758_, _12437_);
  and (_00760_, _00759_, _06071_);
  and (_13328_, _00760_, _00756_);
  and (_00761_, _07105_, _06027_);
  and (_00762_, _00761_, _06840_);
  nand (_00763_, _00762_, _09341_);
  not (_00764_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_00765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00764_);
  not (_00766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00767_, _00766_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_00768_, t1_i);
  and (_00769_, _00768_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00770_, _00769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_00771_, _00770_, _00767_);
  and (_00772_, _00771_, _00765_);
  and (_00773_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00774_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00775_, _00774_, _00773_);
  and (_00776_, _00775_, _00772_);
  and (_00777_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00779_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00780_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00782_, _00780_, _00779_);
  not (_00783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00784_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00785_);
  nor (_00787_, _00786_, _00784_);
  and (_00788_, _09244_, _06012_);
  and (_00789_, _06840_, _00788_);
  nor (_00790_, _00789_, _00787_);
  and (_00791_, _00790_, _00782_);
  not (_00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00793_, _00790_, _00792_);
  and (_00794_, _06840_, _06032_);
  and (_00795_, _00794_, _06027_);
  and (_00796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00797_, _00796_, _00778_);
  and (_00798_, _00797_, _00784_);
  nand (_00799_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00800_, _00799_, _00795_);
  or (_00801_, _00800_, _00793_);
  or (_00802_, _00801_, _00791_);
  or (_00803_, _00762_, _00802_);
  and (_00804_, _00803_, _06071_);
  and (_13336_, _00804_, _00763_);
  and (_00805_, _00367_, _07819_);
  nor (_00806_, _11453_, _11425_);
  and (_00807_, _12469_, _12080_);
  or (_00808_, _00807_, _00806_);
  or (_00809_, _11473_, _11474_);
  not (_00810_, _00809_);
  nand (_00811_, _00810_, _11714_);
  or (_00812_, _00810_, _11714_);
  and (_00813_, _00812_, _11751_);
  and (_00814_, _00813_, _00811_);
  or (_00815_, _00814_, _00808_);
  or (_00816_, _00815_, _00805_);
  or (_00817_, _11428_, _11051_);
  nand (_00818_, _00817_, _12437_);
  or (_00819_, _00818_, _00816_);
  nor (_00820_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00821_, _00820_, _12500_);
  or (_00822_, _00821_, _12437_);
  and (_00823_, _00822_, _06071_);
  and (_13359_, _00823_, _00819_);
  nand (_00824_, _00762_, _06993_);
  and (_00825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_00827_, _00825_, _00789_);
  not (_00828_, _00827_);
  and (_00829_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00830_, _00780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00831_, _00830_, _00784_);
  and (_00832_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_00833_, _00825_);
  nor (_00834_, _00776_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_00835_, _00834_, _00777_);
  and (_00836_, _00835_, _00833_);
  nor (_00837_, _00836_, _00832_);
  nor (_00838_, _00837_, _00789_);
  or (_00839_, _00838_, _00829_);
  or (_00840_, _00839_, _00762_);
  and (_00841_, _00840_, _06071_);
  and (_13363_, _00841_, _00824_);
  and (_00842_, _00774_, _00772_);
  and (_00843_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_00844_, _00843_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00845_, _00844_, _00776_);
  and (_00846_, _00845_, _00827_);
  and (_00847_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_00848_, _00847_, _00846_);
  nand (_00849_, _00831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00850_, _00849_, _00789_);
  or (_00851_, _00850_, _00762_);
  or (_00852_, _00851_, _00848_);
  nand (_00853_, _00762_, _07945_);
  and (_00854_, _00853_, _06071_);
  and (_13366_, _00854_, _00852_);
  nor (_00855_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00856_, _00855_, _00843_);
  nand (_00857_, _00856_, _00827_);
  or (_00858_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00859_, _00858_, _00857_);
  and (_00860_, _07106_, _06027_);
  nand (_00861_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00862_, _00861_, _00795_);
  or (_00863_, _00862_, _00860_);
  or (_00865_, _00863_, _00859_);
  nand (_00866_, _00860_, _06434_);
  and (_00867_, _00866_, _06071_);
  and (_13369_, _00867_, _00865_);
  and (_00868_, _06435_, _06369_);
  or (_00869_, _06438_, _06394_);
  and (_00870_, _00869_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or (_00871_, _00870_, _00868_);
  and (_13371_, _00871_, _06071_);
  nand (_00873_, _00762_, _06609_);
  nor (_00874_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00875_, _00874_, _00778_);
  and (_00876_, _00875_, _00790_);
  not (_00877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00878_, _00790_, _00877_);
  nand (_00879_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_00880_, _00879_, _00795_);
  or (_00881_, _00880_, _00878_);
  or (_00882_, _00881_, _00876_);
  or (_00883_, _00882_, _00762_);
  and (_00884_, _00883_, _06071_);
  and (_13374_, _00884_, _00873_);
  and (_00885_, _00828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00887_, _00775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00889_, _00888_, _00796_);
  and (_00890_, _00889_, _00887_);
  and (_00891_, _00890_, _00784_);
  and (_00892_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00893_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00894_, _00893_, _00892_);
  and (_00895_, _00894_, _00833_);
  nor (_00896_, _00895_, _00891_);
  nor (_00898_, _00896_, _00789_);
  or (_00899_, _00898_, _00860_);
  or (_00900_, _00899_, _00885_);
  nand (_00901_, _00762_, _07977_);
  and (_00902_, _00901_, _06071_);
  and (_13388_, _00902_, _00900_);
  nor (_00903_, _00892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00904_, _00903_, _00842_);
  nand (_00905_, _00904_, _00827_);
  or (_00906_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00907_, _00906_, _00905_);
  nand (_00908_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00909_, _00908_, _00795_);
  or (_00910_, _00909_, _00860_);
  or (_00911_, _00910_, _00907_);
  nand (_00912_, _00762_, _09037_);
  and (_00913_, _00912_, _06071_);
  and (_13392_, _00913_, _00911_);
  not (_00914_, _00762_);
  not (_00915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_00916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00917_, _00916_, _00777_);
  and (_00918_, _00797_, _00786_);
  nor (_00919_, _00918_, _00917_);
  and (_00920_, _00919_, _00915_);
  nor (_00921_, _00919_, _00915_);
  nor (_00922_, _00921_, _00920_);
  nor (_00923_, _00922_, _00789_);
  and (_00924_, _00789_, _07977_);
  or (_00925_, _00924_, _00923_);
  nand (_00926_, _00925_, _00914_);
  nand (_00927_, _00762_, _00915_);
  and (_00928_, _00927_, _06071_);
  and (_13413_, _00928_, _00926_);
  nand (_00929_, _00789_, _09037_);
  or (_00930_, _00921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_00931_, _00921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00932_, _00931_, _00930_);
  or (_00933_, _00932_, _00789_);
  and (_00934_, _00933_, _00914_);
  and (_00935_, _00934_, _00929_);
  and (_00936_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00937_, _00936_, _00935_);
  and (_13416_, _00937_, _06071_);
  nand (_00938_, _00789_, _07945_);
  and (_00939_, _00887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00940_, _00939_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00941_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00942_, _00941_, _00940_);
  and (_00943_, _00942_, _00916_);
  and (_00944_, _00889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00945_, _00944_, _00939_);
  and (_00946_, _00945_, _00772_);
  and (_00947_, _00946_, _00786_);
  nor (_00948_, _00947_, _00943_);
  and (_00949_, _00948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00950_, _00948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00951_, _00950_, _00949_);
  or (_00952_, _00951_, _00789_);
  and (_00953_, _00952_, _00914_);
  and (_00954_, _00953_, _00938_);
  and (_00955_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00956_, _00955_, _00954_);
  and (_13424_, _00956_, _06071_);
  nand (_00957_, _00789_, _06609_);
  and (_00958_, _00946_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00959_, _00958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00960_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_00961_, _00786_);
  and (_00962_, _00890_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00963_, _00962_, _00941_);
  and (_00964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_00965_, _00964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00966_, _00965_, _00963_);
  nor (_00967_, _00966_, _00961_);
  and (_00968_, _00967_, _00960_);
  and (_00969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00970_, _00942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00971_, _00970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00972_, _00971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_00973_, _00916_);
  and (_00974_, _00965_, _00942_);
  nor (_00975_, _00974_, _00973_);
  and (_00976_, _00975_, _00972_);
  or (_00977_, _00976_, _00969_);
  or (_00978_, _00977_, _00968_);
  or (_00979_, _00978_, _00789_);
  and (_00980_, _00979_, _00914_);
  and (_00981_, _00980_, _00957_);
  and (_00982_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00983_, _00982_, _00981_);
  and (_13427_, _00983_, _06071_);
  nand (_00984_, _00789_, _06993_);
  or (_00985_, _00958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_00986_, _00959_, _00961_);
  and (_00987_, _00986_, _00985_);
  and (_00988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_00989_, _00970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_00990_, _00971_, _00973_);
  and (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00988_);
  or (_00993_, _00992_, _00987_);
  or (_00994_, _00993_, _00789_);
  and (_00995_, _00994_, _00914_);
  and (_00996_, _00995_, _00984_);
  and (_00997_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00998_, _00997_, _00996_);
  and (_13430_, _00998_, _06071_);
  not (_01000_, _00795_);
  and (_01001_, _00931_, _01000_);
  or (_01003_, _01001_, _00860_);
  and (_01004_, _01003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_01005_, _01000_, _06434_);
  or (_01007_, _00931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_01008_, _01007_, _00795_);
  nor (_01010_, _01008_, _01005_);
  nor (_01011_, _01010_, _00860_);
  or (_01012_, _01011_, _01004_);
  and (_13433_, _01012_, _06071_);
  and (_01014_, _09576_, _06381_);
  and (_01016_, _13574_, _06011_);
  nand (_01017_, _06392_, _06011_);
  or (_01018_, _01017_, _01016_);
  and (_01020_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_01021_, _01020_, _01014_);
  and (_13436_, _01021_, _06071_);
  not (_01022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_01023_, t0_i);
  and (_01025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01023_);
  nor (_01027_, _01025_, _01022_);
  not (_01029_, _01027_);
  not (_01030_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_01031_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_01032_, _01031_, _01030_);
  and (_01033_, _01032_, _01029_);
  not (_01034_, _01033_);
  and (_01035_, _06840_, _06028_);
  nor (_01037_, _01035_, _01034_);
  or (_01038_, _01037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_01040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_01043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_01044_, _01043_, _01041_);
  and (_01046_, _01044_, _01040_);
  and (_01047_, _01046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_01050_, _01047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01053_, _01051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01055_, _01054_, _01050_);
  and (_01057_, _01033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_01058_, _01057_, _01055_);
  or (_01060_, _01058_, _01035_);
  and (_01061_, _01060_, _01038_);
  and (_01062_, _07754_, _06027_);
  and (_01063_, _01062_, _06840_);
  or (_01064_, _01063_, _01061_);
  nand (_01065_, _01063_, _07977_);
  and (_01066_, _01065_, _06071_);
  and (_13439_, _01066_, _01064_);
  nor (_01068_, _10945_, _06026_);
  and (_01069_, _01068_, _05923_);
  and (_01070_, _01069_, _06807_);
  and (_01072_, _01070_, _06806_);
  and (_01074_, _01072_, _06383_);
  or (_01076_, _01074_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01077_, _01076_, _09250_);
  nand (_01079_, _01074_, _06803_);
  and (_01080_, _01079_, _01077_);
  and (_01081_, _09249_, _07978_);
  or (_01082_, _01081_, _01080_);
  and (_13441_, _01082_, _06071_);
  nor (_01084_, _01057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_01085_, _01057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_01087_, _01085_, _01084_);
  and (_01088_, _01050_, _01033_);
  and (_01089_, _01088_, _01053_);
  and (_01090_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_01091_, _01090_, _01087_);
  nor (_01092_, _01091_, _01035_);
  and (_01093_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_01094_, _01093_, _01092_);
  or (_01095_, _01094_, _01063_);
  nand (_01096_, _01063_, _09037_);
  and (_01097_, _01096_, _06071_);
  and (_13457_, _01097_, _01095_);
  not (_01098_, _01063_);
  and (_01099_, _01044_, _01033_);
  and (_01100_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_01101_, _01100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_01102_, _01101_, _01099_);
  and (_01103_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_01104_, _01103_, _01102_);
  nor (_01105_, _01104_, _01035_);
  and (_01106_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_01107_, _01106_, _01105_);
  and (_01108_, _01107_, _01098_);
  nor (_01109_, _01098_, _07945_);
  or (_01110_, _01109_, _01108_);
  and (_13461_, _01110_, _06071_);
  nor (_01111_, _01085_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_01112_, _01111_, _01100_);
  and (_01113_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_01114_, _01113_, _01112_);
  nor (_01115_, _01114_, _01035_);
  and (_01116_, _01035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_01117_, _01116_, _01115_);
  and (_01118_, _01117_, _01098_);
  nor (_01119_, _01098_, _06434_);
  or (_01120_, _01119_, _01118_);
  and (_13464_, _01120_, _06071_);
  or (_01121_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01122_, _01121_, _06071_);
  or (_01123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_01124_, _01123_, _06453_);
  or (_01125_, _01124_, _06459_);
  and (_01126_, _06463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01127_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01128_, _06467_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01129_, _01128_, _06470_);
  and (_01130_, _01129_, _01127_);
  nand (_01131_, _09237_, _06470_);
  nand (_01132_, _01131_, _06458_);
  or (_01133_, _01132_, _01130_);
  and (_01134_, _01133_, _01125_);
  and (_01136_, _09237_, _06452_);
  or (_01137_, _01136_, _01134_);
  and (_01139_, _01137_, _06474_);
  and (_01140_, _01123_, _06491_);
  or (_01141_, _01140_, _06498_);
  and (_01142_, _09237_, _06483_);
  not (_01143_, _06497_);
  and (_01144_, _06480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_01146_, _01144_, _06483_);
  and (_01147_, _06478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01148_, _01147_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01150_, _01148_, _01146_);
  or (_01151_, _01150_, _01143_);
  or (_01153_, _01151_, _01142_);
  and (_01155_, _01153_, _01141_);
  nand (_01156_, _09237_, _06490_);
  nand (_01158_, _01156_, _06519_);
  or (_01159_, _01158_, _01155_);
  or (_01160_, _06519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_01161_, _01160_, _01159_);
  and (_01163_, _01161_, _06564_);
  or (_01164_, _01163_, _01139_);
  or (_01165_, _01164_, _06508_);
  and (_13475_, _01165_, _01122_);
  nor (_01166_, _06562_, _06508_);
  not (_01167_, _01166_);
  and (_01168_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_01169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_01170_, _01126_, _01169_);
  nand (_01171_, _01170_, _01129_);
  or (_01172_, _09226_, _06471_);
  and (_01173_, _01172_, _01171_);
  or (_01174_, _01173_, _06457_);
  not (_01176_, _06455_);
  not (_01177_, _06457_);
  or (_01178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01179_, _01178_, _01177_);
  and (_01181_, _01179_, _01176_);
  and (_01182_, _01181_, _01174_);
  and (_01183_, _09226_, _06455_);
  or (_01184_, _01183_, _06452_);
  or (_01185_, _01184_, _01182_);
  or (_01186_, _01178_, _06453_);
  and (_01187_, _01186_, _06474_);
  and (_01188_, _01187_, _01185_);
  or (_01190_, _01178_, _06491_);
  and (_01192_, _06519_, _06564_);
  or (_01193_, _01147_, _01169_);
  nand (_01194_, _01193_, _01146_);
  or (_01195_, _09226_, _06484_);
  and (_01197_, _01195_, _01194_);
  or (_01198_, _01197_, _06494_);
  not (_01200_, _06496_);
  not (_01201_, _06494_);
  or (_01203_, _01178_, _01201_);
  and (_01204_, _01203_, _01200_);
  and (_01205_, _01204_, _01198_);
  and (_01206_, _09226_, _06496_);
  or (_01207_, _01206_, _06490_);
  or (_01208_, _01207_, _01205_);
  and (_01209_, _01208_, _01192_);
  and (_01210_, _01209_, _01190_);
  or (_01211_, _01210_, _01188_);
  and (_01212_, _01211_, _06509_);
  or (_01213_, _01212_, _01168_);
  and (_13478_, _01213_, _06071_);
  and (_01214_, _06395_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_01215_, _09576_, _06368_);
  or (_01216_, _01215_, _01214_);
  and (_13487_, _01216_, _06071_);
  nand (_01217_, _00789_, _09341_);
  and (_01218_, _00974_, _00916_);
  and (_01219_, _00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_01220_, _01219_, _00786_);
  nor (_01221_, _01220_, _01218_);
  and (_01222_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_01223_, _01221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_01225_, _01223_, _01222_);
  or (_01226_, _01225_, _00789_);
  and (_01227_, _01226_, _00914_);
  and (_01228_, _01227_, _01217_);
  and (_01229_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_01230_, _01229_, _01228_);
  and (_13497_, _01230_, _06071_);
  nand (_01231_, _01063_, _06609_);
  nor (_01232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_01233_, _01232_);
  and (_01234_, _01099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01235_, _01234_, _01233_);
  not (_01237_, _01235_);
  nor (_01238_, _01237_, _01035_);
  and (_01239_, _01238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_01240_, _01238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_01241_, _01240_, _01239_);
  nand (_01242_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_01243_, _01242_, _01035_);
  or (_01244_, _01243_, _01241_);
  or (_01245_, _01244_, _01063_);
  and (_01246_, _01245_, _06071_);
  and (_13502_, _01246_, _01231_);
  nand (_01248_, _01063_, _09341_);
  not (_01249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_01250_, _01035_, _01249_);
  and (_01251_, _01232_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_01252_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_01253_, _01252_, _01251_);
  and (_01254_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_01255_, _01254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_01256_, _01047_, _01033_);
  and (_01257_, _01256_, _01233_);
  or (_01258_, _01257_, _01035_);
  and (_01259_, _01258_, _01255_);
  or (_01260_, _01259_, _01253_);
  and (_01261_, _01260_, _01250_);
  or (_01262_, _01261_, _01063_);
  and (_01263_, _01262_, _06071_);
  and (_13505_, _01263_, _01248_);
  nand (_01264_, _01063_, _06993_);
  not (_01265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand (_01266_, _01035_, _01265_);
  and (_01267_, _01089_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_01268_, _01099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_01269_, _01268_, _01234_);
  or (_01270_, _01269_, _01267_);
  or (_01271_, _01270_, _01035_);
  and (_01272_, _01271_, _01266_);
  or (_01273_, _01272_, _01063_);
  and (_01274_, _01273_, _06071_);
  and (_13508_, _01274_, _01264_);
  nor (_01276_, _06508_, _06474_);
  or (_01277_, _01276_, _06445_);
  nand (_01279_, _00727_, _06562_);
  and (_01280_, _01279_, _06071_);
  and (_13517_, _01280_, _01277_);
  and (_13520_, _07336_, _06071_);
  not (_01281_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nor (_01282_, _01166_, _01281_);
  or (_01283_, _06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01284_, _01283_, _06453_);
  and (_01285_, _01284_, _06474_);
  and (_01286_, _06467_, _06445_);
  nor (_01287_, _01286_, _06470_);
  and (_01288_, _06463_, _06445_);
  or (_01290_, _01288_, _01281_);
  nand (_01291_, _01290_, _01287_);
  or (_01293_, _09225_, _06471_);
  and (_01294_, _01293_, _01291_);
  or (_01295_, _01294_, _06457_);
  or (_01296_, _01283_, _01177_);
  and (_01297_, _01296_, _01176_);
  and (_01298_, _01297_, _01295_);
  and (_01300_, _09225_, _06455_);
  or (_01301_, _01300_, _06452_);
  or (_01302_, _01301_, _01298_);
  and (_01303_, _01302_, _01285_);
  or (_01304_, _06494_, _06484_);
  and (_01305_, _01304_, _01200_);
  or (_01307_, _01305_, _09225_);
  and (_01308_, _06480_, _06445_);
  nor (_01309_, _01308_, _06483_);
  and (_01310_, _06478_, _06445_);
  nor (_01311_, _01310_, _01281_);
  nor (_01312_, _01311_, _01143_);
  nand (_01313_, _01312_, _01309_);
  and (_01314_, _01313_, _01307_);
  or (_01315_, _01314_, _06490_);
  or (_01316_, _06496_, _01201_);
  and (_01318_, _01316_, _06491_);
  or (_01319_, _01318_, _01283_);
  and (_01320_, _01319_, _01192_);
  and (_01321_, _01320_, _01315_);
  or (_01322_, _01321_, _01303_);
  and (_01323_, _01322_, _06509_);
  or (_01324_, _01323_, _01282_);
  and (_13536_, _01324_, _06071_);
  and (_01325_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_01326_, _06445_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01327_, _01326_, _06453_);
  or (_01329_, _01327_, _06459_);
  or (_01330_, _01288_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01331_, _01330_, _01287_);
  nand (_01332_, _09236_, _06470_);
  nand (_01333_, _01332_, _06458_);
  or (_01334_, _01333_, _01331_);
  and (_01335_, _01334_, _01329_);
  and (_01336_, _09236_, _06452_);
  or (_01337_, _01336_, _01335_);
  and (_01338_, _01337_, _06474_);
  and (_01339_, _06497_, _06483_);
  or (_01340_, _01339_, _06490_);
  and (_01341_, _01340_, _09236_);
  or (_01342_, _01326_, _06497_);
  and (_01343_, _01342_, _06491_);
  or (_01344_, _01310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01345_, _01344_, _01309_);
  or (_01346_, _01345_, _01143_);
  and (_01347_, _01346_, _01343_);
  or (_01349_, _01347_, _01341_);
  and (_01350_, _01349_, _01192_);
  or (_01351_, _01350_, _01338_);
  and (_01352_, _01351_, _06509_);
  or (_01353_, _01352_, _01325_);
  and (_13542_, _01353_, _06071_);
  nand (_01354_, _01035_, _09341_);
  and (_01355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_01356_, _01355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01357_, _01356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01358_, _01357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01360_, _01358_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01361_, _01360_, _01234_);
  nand (_01362_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_01363_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01364_, _01363_, _01232_);
  and (_01365_, _01364_, _01362_);
  and (_01366_, _01360_, _01088_);
  or (_01368_, _01366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_01369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _01369_);
  and (_01371_, _01358_, _01088_);
  and (_01372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01373_, _01372_, _01371_);
  not (_01374_, _01373_);
  and (_01375_, _01374_, _01370_);
  and (_01376_, _01375_, _01368_);
  not (_01377_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01378_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_01379_, _01378_, _01357_);
  and (_01380_, _01379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_01381_, _01380_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_01382_, _01381_, _01377_);
  or (_01383_, _01382_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_01384_, _01372_);
  or (_01385_, _01381_, _01384_);
  and (_01386_, _01385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01387_, _01386_, _01383_);
  or (_01388_, _01387_, _01376_);
  or (_01389_, _01388_, _01365_);
  or (_01390_, _01389_, _01035_);
  and (_01391_, _01390_, _01098_);
  and (_01392_, _01391_, _01354_);
  and (_01393_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_01394_, _01393_, _01392_);
  and (_13545_, _01394_, _06071_);
  nand (_01395_, _01035_, _06609_);
  or (_01396_, _01370_, _01053_);
  and (_01397_, _01371_, _01369_);
  nor (_01398_, _01397_, _01377_);
  and (_01399_, _01397_, _01377_);
  or (_01400_, _01399_, _01398_);
  and (_01401_, _01400_, _01396_);
  and (_01402_, _01378_, _01358_);
  or (_01403_, _01402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_01405_, _01402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01406_, _01405_, _01404_);
  and (_01407_, _01406_, _01403_);
  and (_01409_, _01358_, _01234_);
  or (_01410_, _01409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_01411_, _01361_, _01233_);
  and (_01412_, _01411_, _01410_);
  or (_01413_, _01412_, _01407_);
  or (_01414_, _01413_, _01401_);
  or (_01415_, _01414_, _01035_);
  and (_01416_, _01415_, _01098_);
  and (_01417_, _01416_, _01395_);
  and (_01418_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_01419_, _01418_, _01417_);
  and (_13548_, _01419_, _06071_);
  nand (_01420_, _01035_, _09037_);
  and (_01421_, _01088_, _01369_);
  and (_01422_, _01421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01423_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_01424_, _01422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_01425_, _01424_, _01396_);
  and (_01426_, _01425_, _01423_);
  not (_01427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_01428_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01429_, _01428_, _01427_);
  and (_01430_, _01355_, _01234_);
  nor (_01431_, _01430_, _01233_);
  and (_01432_, _01431_, _01429_);
  and (_01433_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_01434_, _01433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_01435_, _01378_, _01355_);
  not (_01436_, _01435_);
  and (_01437_, _01436_, _01404_);
  and (_01438_, _01437_, _01434_);
  or (_01439_, _01438_, _01432_);
  or (_01440_, _01439_, _01426_);
  or (_01441_, _01440_, _01035_);
  and (_01443_, _01441_, _01420_);
  or (_01444_, _01443_, _01063_);
  nand (_01445_, _01063_, _01427_);
  and (_01446_, _01445_, _06071_);
  and (_13561_, _01446_, _01444_);
  nand (_01447_, _01035_, _06434_);
  or (_01448_, _01430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01449_, _01356_, _01234_);
  nor (_01450_, _01449_, _01233_);
  and (_01451_, _01450_, _01448_);
  and (_01452_, _01355_, _01088_);
  or (_01453_, _01452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01454_, _01356_, _01088_);
  not (_01455_, _01454_);
  and (_01456_, _01455_, _01370_);
  and (_01457_, _01456_, _01453_);
  and (_01458_, _01435_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_01459_, _01458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01460_, _01378_, _01356_);
  nand (_01462_, _01460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01463_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01465_, _01463_, _01459_);
  or (_01466_, _01465_, _01457_);
  or (_01467_, _01466_, _01451_);
  or (_01468_, _01467_, _01035_);
  and (_01469_, _01468_, _01098_);
  and (_01470_, _01469_, _01447_);
  and (_01471_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_01472_, _01471_, _01470_);
  and (_13563_, _01472_, _06071_);
  and (_01473_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01474_, _01473_, _01166_);
  and (_13565_, _01474_, _06071_);
  nor (_01475_, _06478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01476_, _01475_, _06480_);
  or (_01477_, _01476_, _06483_);
  and (_01478_, _01477_, _01201_);
  or (_01479_, _01478_, _06496_);
  and (_01480_, _01479_, _06491_);
  and (_01481_, _01480_, _01192_);
  and (_01482_, _06474_, _06453_);
  nor (_01483_, _06463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01484_, _01483_, _06467_);
  or (_01485_, _01484_, _06470_);
  and (_01486_, _01485_, _01177_);
  or (_01487_, _01486_, _06455_);
  and (_01488_, _01487_, _01482_);
  or (_01489_, _01488_, _06508_);
  or (_01490_, _01489_, _01481_);
  or (_01491_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01492_, _01491_, _06071_);
  and (_13568_, _01492_, _01490_);
  nand (_01493_, _01035_, _07945_);
  and (_01494_, _01454_, _01369_);
  or (_01495_, _01494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_01496_, _01494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01497_, _01496_, _01495_);
  and (_01498_, _01497_, _01396_);
  or (_01499_, _01449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01500_, _01357_, _01234_);
  nor (_01502_, _01500_, _01233_);
  and (_01503_, _01502_, _01499_);
  or (_01504_, _01460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_01506_, _01379_);
  and (_01507_, _01506_, _01404_);
  and (_01508_, _01507_, _01504_);
  or (_01509_, _01508_, _01503_);
  or (_01510_, _01509_, _01498_);
  or (_01511_, _01510_, _01035_);
  and (_01513_, _01511_, _01098_);
  and (_01514_, _01513_, _01493_);
  and (_01516_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_01518_, _01516_, _01514_);
  and (_13571_, _01518_, _06071_);
  and (_13573_, _10924_, _06508_);
  nand (_01519_, _01035_, _06993_);
  and (_01521_, _01357_, _01088_);
  or (_01522_, _01521_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_01523_, _01371_);
  and (_01524_, _01523_, _01370_);
  and (_01525_, _01524_, _01522_);
  or (_01526_, _01500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_01527_, _01409_, _01233_);
  and (_01528_, _01527_, _01526_);
  or (_01529_, _01380_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01530_, _01381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01531_, _01530_, _01529_);
  or (_01532_, _01531_, _01528_);
  or (_01533_, _01532_, _01525_);
  or (_01534_, _01533_, _01035_);
  and (_01535_, _01534_, _01098_);
  and (_01536_, _01535_, _01519_);
  and (_01537_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_01538_, _01537_, _01536_);
  and (_13575_, _01538_, _06071_);
  and (_01539_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01540_, _01539_, _01166_);
  and (_13581_, _01540_, _06071_);
  nand (_01541_, _01035_, _07977_);
  or (_01542_, _01421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_01543_, _01422_);
  and (_01544_, _01543_, _01396_);
  and (_01545_, _01544_, _01542_);
  or (_01546_, _01234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01547_, _01428_, _01232_);
  and (_01548_, _01547_, _01546_);
  or (_01549_, _01378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_01550_, _01433_);
  and (_01551_, _01550_, _01404_);
  and (_01552_, _01551_, _01549_);
  or (_01553_, _01552_, _01548_);
  or (_01554_, _01553_, _01545_);
  or (_01555_, _01554_, _01035_);
  and (_01556_, _01555_, _01541_);
  or (_01557_, _01556_, _01063_);
  or (_01558_, _01098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01559_, _01558_, _06071_);
  and (_13591_, _01559_, _01557_);
  and (_13596_, _11017_, _06508_);
  and (_01560_, _13743_, _06840_);
  nand (_01561_, _01560_, _07977_);
  or (_01562_, _01560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01563_, _01562_, _06071_);
  and (_13600_, _01563_, _01561_);
  nor (_01564_, _06481_, _06488_);
  nand (_01565_, _06517_, _01564_);
  nor (_01566_, _01565_, _06474_);
  and (_01567_, _06508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_01568_, _06508_, _06470_);
  nor (_01569_, _01568_, _06450_);
  not (_01570_, _06468_);
  and (_01571_, _01570_, _06459_);
  and (_01573_, _01571_, _01569_);
  or (_01574_, _01573_, _01567_);
  or (_01576_, _01574_, _01566_);
  and (_13601_, _01576_, _06071_);
  and (_01577_, _12019_, _06369_);
  and (_01578_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_01579_, _01578_, _01577_);
  and (_13605_, _01579_, _06071_);
  and (_01581_, _13751_, _06840_);
  or (_01582_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_01583_, _01582_, _06071_);
  nand (_01584_, _01581_, _06434_);
  and (_13607_, _01584_, _01583_);
  or (_01585_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_01586_, _06530_, _05833_);
  and (_01587_, _01586_, _06071_);
  and (_13610_, _01587_, _01585_);
  or (_01588_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_01589_, _01588_, _06071_);
  nand (_01590_, _01581_, _07945_);
  and (_13612_, _01590_, _01589_);
  nand (_01591_, _01560_, _09037_);
  or (_01592_, _01560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01593_, _01592_, _06071_);
  and (_13615_, _01593_, _01591_);
  or (_01594_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_01595_, _01594_, _06071_);
  nand (_01596_, _01581_, _06609_);
  and (_13622_, _01596_, _01595_);
  or (_01597_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_01598_, _01597_, _06071_);
  nand (_01599_, _01581_, _09341_);
  and (_13624_, _01599_, _01598_);
  or (_01600_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_01601_, _01600_, _06071_);
  nand (_01602_, _01581_, _06993_);
  and (_13626_, _01602_, _01601_);
  and (_01603_, _12120_, _06369_);
  and (_01604_, _13652_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_01605_, _01604_, _01603_);
  and (_13686_, _01605_, _06071_);
  nor (_01606_, _05937_, _05923_);
  and (_01607_, _01606_, _06820_);
  and (_01608_, _01607_, _13722_);
  and (_01609_, _13710_, _10943_);
  not (_01610_, _01609_);
  or (_01611_, _01610_, _10936_);
  and (_01612_, _01611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01613_, _01612_, _01608_);
  nor (_01614_, _10930_, _06479_);
  or (_01615_, _01614_, _10928_);
  and (_01617_, _01615_, _01609_);
  or (_01619_, _01617_, _01613_);
  nand (_01621_, _01608_, _06993_);
  and (_01622_, _01621_, _06071_);
  and (_13768_, _01622_, _01619_);
  not (_01623_, _01608_);
  and (_01625_, _01609_, _07105_);
  or (_01626_, _01625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_01627_, _01626_, _01623_);
  nand (_01628_, _01625_, _06803_);
  and (_01629_, _01628_, _01627_);
  nor (_01630_, _01623_, _07945_);
  or (_01631_, _01630_, _01629_);
  and (_13773_, _01631_, _06071_);
  nor (_01632_, _07753_, _06361_);
  or (_01633_, _01610_, _01632_);
  and (_01634_, _01633_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01635_, _01634_, _01608_);
  and (_01636_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_01637_, _01636_, _00275_);
  and (_01638_, _01637_, _01609_);
  or (_01639_, _01638_, _01635_);
  nand (_01640_, _01608_, _06434_);
  and (_01641_, _01640_, _06071_);
  and (_13775_, _01641_, _01639_);
  and (_13787_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  and (_01643_, _01609_, _08801_);
  or (_01644_, _01643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_01645_, _01644_, _01623_);
  nand (_01646_, _01643_, _06803_);
  and (_01647_, _01646_, _01645_);
  nor (_01649_, _01623_, _09341_);
  or (_01650_, _01649_, _01647_);
  and (_13795_, _01650_, _06071_);
  and (_01652_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_01653_, _11023_, _06610_);
  or (_01654_, _01653_, _01652_);
  and (_13801_, _01654_, _06071_);
  and (_01655_, _10948_, _06362_);
  or (_01656_, _01655_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_01657_, _01656_, _10953_);
  nand (_01659_, _01655_, _06803_);
  and (_01660_, _01659_, _01657_);
  nor (_01661_, _10953_, _09037_);
  or (_01662_, _01661_, _01660_);
  and (_13834_, _01662_, _06071_);
  and (_01664_, _10948_, _06383_);
  and (_01665_, _01664_, _06803_);
  nor (_01666_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_01667_, _01666_, _01665_);
  nand (_01668_, _01667_, _10953_);
  nand (_01669_, _10952_, _07977_);
  and (_01670_, _01669_, _06071_);
  and (_13841_, _01670_, _01668_);
  and (_01671_, _10948_, _08801_);
  and (_01672_, _01671_, _06803_);
  nor (_01674_, _01671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01675_, _01674_, _01672_);
  nand (_01676_, _01675_, _10953_);
  nand (_01677_, _10952_, _09341_);
  and (_01678_, _01677_, _06071_);
  and (_13855_, _01678_, _01676_);
  or (_01680_, _05993_, _05981_);
  nand (_01681_, _01680_, _10948_);
  and (_01682_, _01681_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01683_, _01682_, _10952_);
  or (_01684_, _06005_, _05981_);
  and (_01685_, _01684_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_01686_, _01685_, _08943_);
  and (_01687_, _01686_, _10948_);
  or (_01688_, _01687_, _01683_);
  nand (_01689_, _10952_, _06609_);
  and (_01690_, _01689_, _06071_);
  and (_13859_, _01690_, _01688_);
  not (_01691_, _10948_);
  or (_01692_, _01691_, _10936_);
  and (_01693_, _01692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_01694_, _01693_, _10952_);
  nor (_01695_, _10930_, _06464_);
  or (_01696_, _01695_, _10928_);
  and (_01697_, _01696_, _10948_);
  or (_01698_, _01697_, _01694_);
  nand (_01699_, _10952_, _06993_);
  and (_01700_, _01699_, _06071_);
  and (_13862_, _01700_, _01698_);
  and (_01701_, _10948_, _07105_);
  or (_01702_, _01701_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01703_, _01702_, _10953_);
  nand (_01704_, _01701_, _06803_);
  and (_01706_, _01704_, _01703_);
  nor (_01707_, _10953_, _07945_);
  or (_01708_, _01707_, _01706_);
  and (_13868_, _01708_, _06071_);
  nor (_13941_, _12084_, rst);
  nand (_13965_, _12397_, _06071_);
  nor (_13984_, _12098_, rst);
  nor (_13989_, _12142_, rst);
  nor (_13992_, _12212_, rst);
  and (_13995_, _11961_, _06071_);
  nand (_14001_, _12378_, _06071_);
  and (_00014_, _07342_, _06071_);
  and (_00186_, _08028_, _06071_);
  and (_00258_, t2ex_i, _06071_);
  and (_01709_, _09348_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand (_01710_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_01711_, _01710_, _09346_);
  nor (_01712_, _06609_, _06400_);
  or (_01713_, _01712_, _01711_);
  or (_01714_, _01713_, _01709_);
  and (_00264_, _01714_, _06071_);
  and (_00321_, _12076_, _06071_);
  and (_00359_, _07781_, _06071_);
  nor (_01715_, _12274_, _11403_);
  nor (_01717_, _01715_, _11795_);
  or (_01718_, _11876_, _11869_);
  or (_01720_, _01718_, _12268_);
  or (_01721_, _11845_, _11828_);
  or (_01722_, _11881_, _11865_);
  or (_01723_, _01722_, _01721_);
  or (_01724_, _01723_, _01720_);
  or (_01725_, _01724_, _11843_);
  and (_01726_, _01725_, _11421_);
  or (_01727_, _01726_, _01717_);
  and (_00388_, _01727_, _06071_);
  and (_01728_, _09228_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_01729_, _09239_, _09233_);
  nand (_01731_, _01729_, _01728_);
  nand (_01733_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_01735_, _01733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_01737_, _06840_, _06380_);
  nor (_01738_, _01737_, _10945_);
  or (_01740_, _01738_, _01735_);
  nand (_01741_, _01738_, _08799_);
  and (_01742_, _01741_, _01740_);
  nand (_01744_, _01742_, _09250_);
  nand (_01745_, _09249_, _09037_);
  and (_01746_, _01745_, _06071_);
  and (_00430_, _01746_, _01744_);
  nand (_01747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01748_, _01728_, _09240_);
  nor (_01749_, _01748_, _01747_);
  and (_01750_, _07105_, _06378_);
  nand (_01751_, _01750_, _06840_);
  or (_01752_, _01751_, _10945_);
  nand (_01753_, _01752_, _01749_);
  or (_01754_, _01752_, _06803_);
  and (_01755_, _01754_, _01753_);
  nand (_01757_, _01755_, _09250_);
  nand (_01758_, _09249_, _07945_);
  and (_01759_, _01758_, _06071_);
  and (_00433_, _01759_, _01757_);
  and (_01760_, _01609_, _06805_);
  or (_01761_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01762_, _01761_, _01623_);
  nand (_01764_, _01760_, _06803_);
  and (_01765_, _01764_, _01762_);
  nor (_01766_, _01623_, _06359_);
  or (_01767_, _01766_, _01765_);
  and (_00470_, _01767_, _06071_);
  and (_01768_, _01068_, _06805_);
  and (_01769_, _01768_, _06840_);
  and (_01770_, _01769_, _06803_);
  and (_01771_, _09238_, _09233_);
  nand (_01772_, _01771_, _09229_);
  nand (_01773_, _01772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_01774_, _01773_, _07876_);
  nor (_01775_, _01774_, _01769_);
  or (_01776_, _01775_, _01770_);
  nand (_01777_, _01776_, _09250_);
  nand (_01778_, _09249_, _06359_);
  and (_01779_, _01778_, _06071_);
  and (_00475_, _01779_, _01777_);
  and (_00531_, _11392_, _06071_);
  nor (_00563_, _11533_, rst);
  and (_00574_, _00646_, _06071_);
  and (_01780_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08003_);
  and (_01781_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01782_, _01781_, _01780_);
  and (_00592_, _01782_, _06071_);
  and (_01783_, _07824_, _06809_);
  nand (_01784_, _01783_, _06383_);
  or (_01785_, _01784_, _00593_);
  not (_01786_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_01787_, _01784_, _01786_);
  and (_01788_, _01787_, _06012_);
  and (_01789_, _01788_, _01785_);
  nor (_01790_, _06814_, _01786_);
  not (_01791_, _01783_);
  or (_01792_, _01791_, _10936_);
  and (_01793_, _01792_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_01794_, _10930_, _01786_);
  or (_01795_, _01794_, _10928_);
  and (_01796_, _01795_, _01783_);
  or (_01797_, _01796_, _01793_);
  and (_01798_, _01797_, _06815_);
  or (_01799_, _01798_, _01790_);
  or (_01800_, _01799_, _01789_);
  and (_00618_, _01800_, _06071_);
  or (_01801_, _01784_, _00612_);
  not (_01802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_01803_, _01784_, _01802_);
  and (_01804_, _01803_, _06012_);
  and (_01805_, _01804_, _01801_);
  nor (_01806_, _06814_, _01802_);
  and (_01807_, _01783_, _07105_);
  nand (_01808_, _01807_, _06803_);
  or (_01809_, _01807_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01810_, _01809_, _06815_);
  and (_01811_, _01810_, _01808_);
  or (_01812_, _01811_, _01806_);
  or (_01813_, _01812_, _01805_);
  and (_00621_, _01813_, _06071_);
  or (_01814_, _01784_, _07425_);
  not (_01815_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_01817_, _01784_, _01815_);
  and (_01818_, _01817_, _06012_);
  and (_01819_, _01818_, _01814_);
  nor (_01820_, _06814_, _01815_);
  and (_01821_, _01783_, _08801_);
  nand (_01822_, _01821_, _06803_);
  or (_01823_, _01821_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01824_, _01823_, _06815_);
  and (_01825_, _01824_, _01822_);
  or (_01826_, _01825_, _01820_);
  or (_01827_, _01826_, _01819_);
  and (_00641_, _01827_, _06071_);
  and (pc_log_change, _08705_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_01828_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_01830_, pc_log_change, _06086_);
  and (_01831_, _01830_, _06071_);
  and (_00725_, _01831_, _01828_);
  and (_01832_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08003_);
  and (_01833_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01834_, _01833_, _01832_);
  and (_00728_, _01834_, _06071_);
  and (_01836_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_01837_, _07945_, _06611_);
  or (_01838_, _01837_, _01836_);
  and (_00781_, _01838_, _06071_);
  and (_01839_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_01840_, _06611_, _06359_);
  or (_01841_, _01840_, _01839_);
  and (_00826_, _01841_, _06071_);
  nor (_00864_, _11965_, rst);
  nand (_01842_, _07977_, _07946_);
  or (_01843_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_01844_, _01843_, _01842_);
  and (_00872_, _01844_, _06071_);
  or (_01845_, _01784_, _00655_);
  not (_01846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_01847_, _01784_, _01846_);
  and (_01848_, _01847_, _06012_);
  and (_01849_, _01848_, _01845_);
  nor (_01850_, _06814_, _01846_);
  and (_01852_, _01783_, _06362_);
  nand (_01853_, _01852_, _06803_);
  or (_01854_, _01852_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01855_, _01854_, _06815_);
  and (_01856_, _01855_, _01853_);
  or (_01857_, _01856_, _01850_);
  or (_01858_, _01857_, _01849_);
  and (_00886_, _01858_, _06071_);
  or (_01859_, _01784_, _00660_);
  not (_01860_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_01861_, _01784_, _01860_);
  and (_01862_, _01861_, _06012_);
  and (_01863_, _01862_, _01859_);
  nor (_01864_, _06814_, _01860_);
  or (_01865_, _01784_, _08799_);
  and (_01866_, _01861_, _06815_);
  and (_01867_, _01866_, _01865_);
  or (_01868_, _01867_, _01864_);
  or (_01869_, _01868_, _01863_);
  and (_00897_, _01869_, _06071_);
  or (_01871_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not (_01872_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01873_, pc_log_change, _01872_);
  and (_01874_, _01873_, _06071_);
  and (_00999_, _01874_, _01871_);
  or (_01875_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_01876_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01877_, pc_log_change, _01876_);
  and (_01878_, _01877_, _06071_);
  and (_01002_, _01878_, _01875_);
  or (_01879_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_01880_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_01881_, pc_log_change, _01880_);
  and (_01882_, _01881_, _06071_);
  and (_01006_, _01882_, _01879_);
  and (_01883_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_01884_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_01885_, pc_log_change, _01884_);
  or (_01886_, _01885_, _01883_);
  and (_01009_, _01886_, _06071_);
  not (_01887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_01888_, _06062_, _01887_);
  or (_01889_, _01888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_01891_, _10947_, _09026_);
  or (_01892_, _01891_, _01889_);
  not (_01893_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_01894_, _08801_, _01893_);
  nand (_01895_, _01894_, _01891_);
  or (_01896_, _01895_, _08802_);
  and (_01897_, _01896_, _01892_);
  and (_01898_, _09248_, _05969_);
  or (_01899_, _01898_, _01897_);
  nand (_01900_, _01898_, _09341_);
  and (_01901_, _01900_, _06071_);
  and (_01013_, _01901_, _01899_);
  not (_01903_, _01898_);
  and (_01904_, _01891_, _06032_);
  or (_01905_, _01904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01906_, _01905_, _01903_);
  nand (_01907_, _01904_, _06803_);
  and (_01908_, _01907_, _01906_);
  nor (_01909_, _01903_, _06609_);
  or (_01910_, _01909_, _01908_);
  and (_01015_, _01910_, _06071_);
  not (_01911_, _01891_);
  or (_01912_, _01911_, _10936_);
  and (_01913_, _01912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_01915_, _01913_, _01898_);
  not (_01916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_01917_, _10930_, _01916_);
  or (_01918_, _01917_, _10928_);
  and (_01919_, _01918_, _01891_);
  or (_01920_, _01919_, _01915_);
  nand (_01921_, _01898_, _06993_);
  and (_01922_, _01921_, _06071_);
  and (_01019_, _01922_, _01920_);
  nor (_01923_, _01035_, rst);
  and (_01924_, _01034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and (_01925_, _01372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01926_, _01925_, _01358_);
  nand (_01927_, _01926_, _01234_);
  and (_01928_, _01927_, _01232_);
  or (_01929_, _01926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_01930_, _01929_, _01088_);
  nor (_01931_, _01930_, _01232_);
  nor (_01932_, _01931_, _01928_);
  nor (_01933_, _01932_, _01924_);
  nor (_01934_, _01933_, _01063_);
  and (_01024_, _01934_, _01923_);
  and (_01935_, _01373_, _01369_);
  or (_01936_, _01935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01937_, _01925_, _01397_);
  and (_01938_, _01937_, _01396_);
  and (_01939_, _01938_, _01936_);
  not (_01940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01941_, _01362_, _01940_);
  and (_01942_, _01941_, _01928_);
  and (_01943_, _01402_, _01372_);
  or (_01944_, _01943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01945_, _01925_, _01402_);
  not (_01946_, _01945_);
  and (_01947_, _01946_, _01404_);
  and (_01948_, _01947_, _01944_);
  or (_01949_, _01948_, _01942_);
  nor (_01950_, _01949_, _01939_);
  nor (_01951_, _01950_, _01035_);
  and (_01952_, _01035_, _06360_);
  or (_01953_, _01952_, _01951_);
  and (_01954_, _01953_, _01098_);
  and (_01955_, _01063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01956_, _01955_, _01954_);
  and (_01026_, _01956_, _06071_);
  nand (_01957_, _01063_, _06359_);
  and (_01958_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_01959_, _01958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_01960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01369_);
  nand (_01961_, _01960_, _01051_);
  nand (_01962_, _01961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_01963_, _01962_, _01256_);
  or (_01964_, _01963_, _01035_);
  and (_01965_, _01964_, _01959_);
  or (_01966_, _01965_, _01063_);
  and (_01967_, _01966_, _06071_);
  and (_01028_, _01967_, _01957_);
  and (_01968_, _01891_, _07105_);
  or (_01969_, _01968_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_01970_, _01969_, _01903_);
  nand (_01971_, _01968_, _06803_);
  and (_01972_, _01971_, _01970_);
  nor (_01973_, _01903_, _07945_);
  or (_01974_, _01973_, _01972_);
  and (_01036_, _01974_, _06071_);
  or (_01975_, _01581_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_01976_, _01975_, _06071_);
  nand (_01977_, _01581_, _06359_);
  and (_01039_, _01977_, _01976_);
  or (_01978_, _01911_, _01632_);
  and (_01979_, _01978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01980_, _01979_, _01898_);
  and (_01981_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_01982_, _01981_, _00275_);
  and (_01983_, _01982_, _01891_);
  or (_01984_, _01983_, _01980_);
  nand (_01985_, _01898_, _06434_);
  and (_01986_, _01985_, _06071_);
  and (_01042_, _01986_, _01984_);
  or (_01987_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01988_, pc_log_change, _06243_);
  and (_01989_, _01988_, _06071_);
  and (_01045_, _01989_, _01987_);
  not (_01990_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_01991_, _01378_, _01990_);
  or (_01992_, _01991_, _01945_);
  nand (_01993_, _01992_, _01404_);
  nor (_01994_, _01993_, _01063_);
  and (_01049_, _01994_, _01923_);
  and (_01995_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_01996_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_01997_, pc_log_change, _01996_);
  or (_01998_, _01997_, _01995_);
  and (_01052_, _01998_, _06071_);
  and (_01999_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_02000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_02001_, pc_log_change, _02000_);
  or (_02002_, _02001_, _01999_);
  and (_01056_, _02002_, _06071_);
  and (_02003_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_02004_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_02005_, pc_log_change, _02004_);
  or (_02006_, _02005_, _02003_);
  and (_01059_, _02006_, _06071_);
  and (_01067_, t0_i, _06071_);
  nand (_02007_, _00762_, _06359_);
  not (_02008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_02009_, _00790_, _02008_);
  or (_02010_, _00780_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_02011_, _00797_, _00787_);
  and (_02012_, _02011_, _02010_);
  and (_02013_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02014_, _02013_, _02012_);
  nor (_02015_, _02014_, _00789_);
  or (_02016_, _02015_, _02009_);
  or (_02017_, _02016_, _00762_);
  and (_02018_, _02017_, _06071_);
  and (_01071_, _02018_, _02007_);
  not (_02019_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_02020_, _00772_, _02019_);
  and (_02021_, _00772_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02022_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02023_, _00965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02024_, _02023_, _02022_);
  and (_02026_, _02024_, _02021_);
  or (_02027_, _02026_, _02020_);
  and (_02028_, _02027_, _00916_);
  and (_02029_, _02021_, _02023_);
  and (_02030_, _02029_, _00945_);
  or (_02031_, _02030_, _02020_);
  and (_02032_, _02031_, _00786_);
  nand (_02033_, _00772_, _00783_);
  and (_02034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02035_, _02034_, _02033_);
  or (_02036_, _02035_, _02032_);
  or (_02037_, _02036_, _00798_);
  or (_02038_, _02037_, _02028_);
  nand (_02039_, _02038_, _06071_);
  nor (_02040_, _02039_, _00860_);
  and (_01073_, _02040_, _01000_);
  nand (_02042_, _00789_, _06359_);
  nand (_02043_, _01220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02044_, _00916_, _00772_);
  and (_02045_, _02044_, _02023_);
  nand (_02046_, _02045_, _02022_);
  and (_02047_, _02046_, _02043_);
  nor (_02048_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_02049_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02050_, _02049_, _02048_);
  or (_02051_, _02050_, _00789_);
  and (_02052_, _02051_, _00914_);
  and (_02053_, _02052_, _02042_);
  and (_02054_, _00762_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02055_, _02054_, _02053_);
  and (_01075_, _02055_, _06071_);
  and (_01078_, t1_i, _06071_);
  and (_02056_, _01891_, _06362_);
  or (_02057_, _02056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_02058_, _02057_, _01903_);
  nand (_02059_, _02056_, _06803_);
  and (_02060_, _02059_, _02058_);
  nor (_02061_, _01903_, _09037_);
  or (_02062_, _02061_, _02060_);
  and (_01083_, _02062_, _06071_);
  and (_02063_, _01891_, _06383_);
  or (_02064_, _02063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_02065_, _02064_, _01903_);
  nand (_02066_, _02063_, _06803_);
  and (_02067_, _02066_, _02065_);
  and (_02068_, _01898_, _07978_);
  or (_02069_, _02068_, _02067_);
  and (_01086_, _02069_, _06071_);
  or (_02070_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_02071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_02072_, pc_log_change, _02071_);
  and (_02073_, _02072_, _06071_);
  and (_01135_, _02073_, _02070_);
  or (_02075_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not (_02076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_02077_, pc_log_change, _02076_);
  and (_02078_, _02077_, _06071_);
  and (_01138_, _02078_, _02075_);
  and (_02079_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_02081_, pc_log_change, _01872_);
  or (_02082_, _02081_, _02079_);
  and (_01145_, _02082_, _06071_);
  nand (_02083_, _09341_, _06035_);
  or (_02084_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_02085_, _06541_, _06065_);
  and (_02086_, _02085_, _02084_);
  or (_02087_, _06548_, _06065_);
  and (_02088_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_02089_, _02088_, _02086_);
  nand (_02090_, _02089_, _06036_);
  not (_02091_, _06029_);
  or (_02092_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_02093_, _02092_, _06071_);
  and (_02095_, _02093_, _02090_);
  and (_01149_, _02095_, _02083_);
  and (_02096_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_02097_, pc_log_change, _01880_);
  or (_02098_, _02097_, _02096_);
  and (_01152_, _02098_, _06071_);
  and (_02100_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not (_02101_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand (_02102_, _06065_, _02101_);
  not (_02103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_02105_, _06538_, _06045_);
  and (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_02107_, _02106_, _02103_);
  nor (_02108_, _02106_, _02103_);
  and (_02109_, _06548_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_02110_, _02109_, _06065_);
  or (_02111_, _02110_, _02108_);
  or (_02112_, _02111_, _02107_);
  and (_02113_, _02112_, _02102_);
  and (_02114_, _02113_, _06036_);
  or (_02115_, _02114_, _02100_);
  nor (_02116_, _06609_, _06555_);
  or (_02117_, _02116_, _02115_);
  and (_01154_, _02117_, _06071_);
  nand (_02118_, _06993_, _06035_);
  or (_02119_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_02120_, _02106_, _06065_);
  and (_02121_, _02120_, _02119_);
  and (_02122_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_02123_, _02122_, _02121_);
  nand (_02124_, _02123_, _06036_);
  or (_02125_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_02126_, _02125_, _06071_);
  and (_02127_, _02126_, _02124_);
  and (_01157_, _02127_, _02118_);
  and (_02128_, _06044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_02129_, _02128_, _06059_);
  and (_02130_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_02131_, _02130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_02132_, _02105_, _06065_);
  and (_02133_, _02132_, _02131_);
  and (_02134_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_02135_, _02134_, _02133_);
  nand (_02136_, _02135_, _06036_);
  nand (_02137_, _07945_, _06035_);
  or (_02138_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_02139_, _02138_, _06071_);
  and (_02140_, _02139_, _02137_);
  and (_01162_, _02140_, _02136_);
  and (_02141_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_02142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_02143_, pc_log_change, _02142_);
  or (_02144_, _02143_, _02141_);
  and (_01175_, _02144_, _06071_);
  and (_02145_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_02146_, pc_log_change, _02071_);
  or (_02147_, _02146_, _02145_);
  and (_01180_, _02147_, _06071_);
  and (_02148_, _11023_, _08864_);
  and (_02150_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_02151_, _02150_, _02148_);
  and (_01189_, _02151_, _06071_);
  nor (_02152_, _06538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_02153_, _02152_, _02130_);
  and (_02154_, _02153_, _06066_);
  and (_02155_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_02156_, _02155_, _02154_);
  nand (_02157_, _02156_, _06036_);
  nand (_02158_, _06434_, _06035_);
  or (_02159_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_02160_, _02159_, _06071_);
  and (_02161_, _02160_, _02158_);
  and (_01191_, _02161_, _02157_);
  and (_02162_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_02163_, _06537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_02164_, _06538_, _06065_);
  and (_02165_, _02164_, _02163_);
  nor (_02166_, _02165_, _02162_);
  nand (_02167_, _02166_, _06036_);
  nand (_02168_, _09037_, _06035_);
  or (_02169_, _02091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_02170_, _02169_, _06071_);
  and (_02171_, _02170_, _02168_);
  and (_01196_, _02171_, _02167_);
  or (_02172_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_02173_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_02174_, pc_log_change, _02173_);
  and (_02176_, _02174_, _06071_);
  and (_01199_, _02176_, _02172_);
  and (_02177_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_02178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_02179_, pc_log_change, _02178_);
  or (_02180_, _02179_, _02177_);
  and (_01202_, _02180_, _06071_);
  or (_02181_, _06066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_02182_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_02183_, _02182_, _06547_);
  and (_02184_, _06059_, _06043_);
  nor (_02185_, _02184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_02187_, _02185_, _06537_);
  or (_02188_, _02187_, _06065_);
  or (_02189_, _02188_, _02183_);
  and (_02190_, _02189_, _02181_);
  and (_02191_, _02190_, _06036_);
  and (_02192_, _06029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_02193_, _00788_, _05969_);
  and (_02194_, _07978_, _02193_);
  or (_02195_, _02194_, _02192_);
  or (_02196_, _02195_, _02191_);
  and (_01224_, _02196_, _06071_);
  nor (_02198_, _08865_, _06434_);
  and (_02199_, _01018_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_02200_, _02199_, _02198_);
  and (_01236_, _02200_, _06071_);
  and (_02201_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_02202_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  or (_02203_, _02202_, _02201_);
  and (_01247_, _02203_, _06071_);
  nor (_02204_, _06609_, _02091_);
  not (_02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_02206_, _06059_, _06040_);
  nor (_02207_, _02206_, _02205_);
  and (_02208_, _02206_, _02205_);
  or (_02209_, _02208_, _02207_);
  and (_02210_, _02209_, _06066_);
  and (_02211_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_02212_, _02211_, _02210_);
  and (_02213_, _02212_, _06036_);
  and (_02214_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_02215_, _02214_, _02213_);
  or (_02216_, _02215_, _02204_);
  and (_01275_, _02216_, _06071_);
  nor (_01278_, _11591_, rst);
  nor (_02217_, _09341_, _02091_);
  or (_02218_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_02219_, _06041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_02220_, _06059_, _06042_);
  and (_02221_, _02220_, _02219_);
  and (_02222_, _06547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_02223_, _02222_, _02221_);
  and (_02224_, _02223_, _02218_);
  or (_02225_, _02224_, _06065_);
  not (_02226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand (_02227_, _06065_, _02226_);
  and (_02228_, _02227_, _02225_);
  and (_02229_, _02228_, _06036_);
  and (_02230_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_02231_, _02230_, _02229_);
  or (_02232_, _02231_, _02217_);
  and (_01289_, _02232_, _06071_);
  nor (_02233_, _06993_, _02091_);
  and (_02234_, _06059_, _06039_);
  or (_02235_, _02234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_02236_, _02206_, _06065_);
  and (_02237_, _02236_, _02235_);
  and (_02238_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_02240_, _02238_, _02237_);
  and (_02241_, _02240_, _06036_);
  and (_02242_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_02243_, _02242_, _02241_);
  or (_02244_, _02243_, _02233_);
  and (_01292_, _02244_, _06071_);
  and (_01299_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06071_);
  and (_02245_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_01306_, _02245_, _08574_);
  nor (_02246_, _07344_, _06861_);
  and (_02247_, _06866_, _07344_);
  or (_02248_, _02247_, _02246_);
  and (_01317_, _02248_, _06071_);
  and (_02249_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_02250_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_02251_, _02250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_02252_, _06059_, _06037_);
  nor (_02253_, _02252_, _06065_);
  and (_02254_, _02253_, _02251_);
  or (_02256_, _02254_, _02249_);
  and (_02257_, _02256_, _06036_);
  nor (_02258_, _09037_, _02091_);
  and (_02259_, _06035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_02260_, _02259_, _02258_);
  or (_02262_, _02260_, _02257_);
  and (_01328_, _02262_, _06071_);
  nand (_02263_, _07945_, _06029_);
  and (_02264_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02265_, _06059_, _06038_);
  or (_02266_, _02265_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_02267_, _02234_, _06065_);
  and (_02268_, _02267_, _02266_);
  or (_02269_, _02268_, _02264_);
  or (_02270_, _02269_, _06029_);
  and (_02271_, _02270_, _02263_);
  or (_02272_, _02271_, _02193_);
  not (_02273_, _02193_);
  or (_02275_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_02276_, _02275_, _06071_);
  and (_01348_, _02276_, _02272_);
  nand (_02277_, _06434_, _06029_);
  and (_02278_, _02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_02279_, _02252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_02280_, _02265_, _06065_);
  and (_02281_, _02280_, _02279_);
  or (_02282_, _02281_, _02278_);
  or (_02283_, _02282_, _06029_);
  and (_02284_, _02283_, _02277_);
  or (_02285_, _02284_, _02193_);
  or (_02286_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_02287_, _02286_, _06071_);
  and (_01359_, _02287_, _02285_);
  or (_02288_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_02289_, _06547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_02290_, _02289_, _02250_);
  and (_02291_, _02290_, _02288_);
  or (_02292_, _02291_, _06065_);
  not (_02293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_02294_, _06065_, _02293_);
  and (_02295_, _02294_, _02292_);
  and (_02296_, _02295_, _06036_);
  and (_02297_, _07978_, _06029_);
  and (_02298_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_02299_, _02298_, _02297_);
  or (_02300_, _02299_, _02296_);
  and (_01367_, _02300_, _06071_);
  and (_02301_, _00437_, _08993_);
  nor (_02302_, _02301_, _07890_);
  and (_02303_, _07901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02304_, _02303_, _02302_);
  and (_02305_, _02304_, _07913_);
  nand (_02306_, _07898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_02307_, _02306_, _06560_);
  or (_01408_, _02307_, _02305_);
  nand (_02308_, _09341_, _07946_);
  or (_02309_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02310_, _02309_, _06071_);
  and (_01442_, _02310_, _02308_);
  nor (_01461_, _07874_, rst);
  and (_02311_, _00761_, _05969_);
  nand (_02312_, _02311_, _09341_);
  and (_02313_, _06545_, _06062_);
  not (_02314_, _02313_);
  and (_02315_, _01062_, _05969_);
  nor (_02316_, _02315_, _02314_);
  not (_02317_, _02316_);
  and (_02318_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_02319_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_02320_, _02319_, _02318_);
  or (_02321_, _02311_, _02320_);
  and (_02322_, _02321_, _06071_);
  and (_01464_, _02322_, _02312_);
  and (_02323_, _07105_, _06033_);
  or (_02324_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_02325_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_02326_, _02325_, _02324_);
  or (_02327_, _02326_, _02323_);
  nand (_02328_, _02311_, _09037_);
  and (_02329_, _02328_, _06071_);
  and (_01501_, _02329_, _02327_);
  nand (_02330_, _02311_, _06609_);
  nor (_02331_, _02316_, _02101_);
  and (_02332_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_02333_, _02332_, _02331_);
  or (_02334_, _02333_, _02311_);
  and (_02335_, _02334_, _06071_);
  and (_01505_, _02335_, _02330_);
  nand (_02336_, _02311_, _06993_);
  and (_02337_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_02338_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_02339_, _02338_, _02337_);
  or (_02340_, _02339_, _02311_);
  and (_02341_, _02340_, _06071_);
  and (_01512_, _02341_, _02336_);
  and (_02342_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_02343_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_02344_, _02343_, _02342_);
  or (_02345_, _02344_, _02311_);
  nand (_02346_, _02311_, _07945_);
  and (_02347_, _02346_, _06071_);
  and (_01515_, _02347_, _02345_);
  and (_02348_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_02349_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_02350_, _02349_, _02348_);
  or (_02351_, _02350_, _02311_);
  nand (_02352_, _02311_, _06434_);
  and (_02353_, _02352_, _06071_);
  and (_01517_, _02353_, _02351_);
  or (_02354_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_02355_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_02356_, _02355_, _02354_);
  or (_02357_, _02356_, _02323_);
  nand (_02358_, _02311_, _07977_);
  and (_02359_, _02358_, _06071_);
  and (_01520_, _02359_, _02357_);
  not (_02360_, _02315_);
  nor (_02361_, _02360_, _09341_);
  nor (_02362_, _02313_, _02226_);
  and (_02363_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_02364_, _02363_, _02362_);
  nor (_02365_, _02364_, _02315_);
  or (_02366_, _02365_, _02323_);
  or (_02367_, _02366_, _02361_);
  nand (_02368_, _02323_, _02226_);
  and (_02369_, _02368_, _06071_);
  and (_01572_, _02369_, _02367_);
  nand (_02370_, _02315_, _06609_);
  not (_02371_, _02311_);
  and (_02372_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_02373_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_02374_, _02373_, _02372_);
  or (_02375_, _02374_, _02315_);
  and (_02376_, _02375_, _02371_);
  and (_02377_, _02376_, _02370_);
  and (_02378_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_02379_, _02378_, _02377_);
  and (_01575_, _02379_, _06071_);
  nand (_02380_, _02315_, _06993_);
  and (_02381_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_02382_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_02383_, _02382_, _02381_);
  or (_02384_, _02383_, _02315_);
  and (_02385_, _02384_, _02371_);
  and (_02386_, _02385_, _02380_);
  and (_02387_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_02388_, _02387_, _02386_);
  and (_01580_, _02388_, _06071_);
  nand (_02389_, _02315_, _07945_);
  and (_02390_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02391_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_02392_, _02391_, _02390_);
  or (_02393_, _02392_, _02315_);
  and (_02394_, _02393_, _02371_);
  and (_02395_, _02394_, _02389_);
  and (_02396_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_02397_, _02396_, _02395_);
  and (_01616_, _02397_, _06071_);
  nand (_02399_, _02315_, _06434_);
  and (_02401_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02402_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_02403_, _02402_, _02401_);
  or (_02404_, _02403_, _02315_);
  and (_02405_, _02404_, _02371_);
  and (_02406_, _02405_, _02399_);
  and (_02407_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_02408_, _02407_, _02406_);
  and (_01618_, _02408_, _06071_);
  nand (_02409_, _02315_, _09037_);
  or (_02410_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02411_, _02314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_02412_, _02411_, _02410_);
  or (_02413_, _02412_, _02315_);
  and (_02414_, _02413_, _02371_);
  and (_02415_, _02414_, _02409_);
  and (_02416_, _02311_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02417_, _02416_, _02415_);
  and (_01620_, _02417_, _06071_);
  nor (_02418_, _02313_, _02293_);
  and (_02419_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_02420_, _02419_, _02418_);
  or (_02421_, _02420_, _02315_);
  nand (_02422_, _02315_, _07977_);
  and (_02423_, _02422_, _02421_);
  or (_02424_, _02423_, _02323_);
  nand (_02425_, _02311_, _02293_);
  and (_02426_, _02425_, _06071_);
  and (_01624_, _02426_, _02424_);
  and (_02428_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_02429_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_02430_, pc_log_change, _02429_);
  or (_02431_, _02430_, _02428_);
  and (_01642_, _02431_, _06071_);
  and (_02432_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_02433_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_02434_, pc_log_change, _02433_);
  or (_02435_, _02434_, _02432_);
  and (_01648_, _02435_, _06071_);
  and (_02436_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_02437_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_02438_, pc_log_change, _02437_);
  or (_02439_, _02438_, _02436_);
  and (_01651_, _02439_, _06071_);
  and (_02440_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_02441_, pc_log_change, _02076_);
  or (_02442_, _02441_, _02440_);
  and (_01658_, _02442_, _06071_);
  or (_02443_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_02444_, pc_log_change, _06210_);
  and (_02445_, _02444_, _06071_);
  and (_01663_, _02445_, _02443_);
  and (_02446_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_02447_, pc_log_change, _01876_);
  or (_02448_, _02447_, _02446_);
  and (_01673_, _02448_, _06071_);
  and (_02449_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02450_, pc_log_change, _02173_);
  or (_02451_, _02450_, _02449_);
  and (_01679_, _02451_, _06071_);
  and (_01705_, t2_i, _06071_);
  and (_02452_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_02453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_02454_, pc_log_change, _02453_);
  or (_02455_, _02454_, _02452_);
  and (_01716_, _02455_, _06071_);
  and (_02456_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_02457_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_02458_, pc_log_change, _02457_);
  or (_02459_, _02458_, _02456_);
  and (_01719_, _02459_, _06071_);
  and (_02460_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_02461_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_02462_, pc_log_change, _02461_);
  or (_02463_, _02462_, _02460_);
  and (_01730_, _02463_, _06071_);
  or (_02464_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand (_02465_, pc_log_change, _01996_);
  and (_02467_, _02465_, _06071_);
  and (_01732_, _02467_, _02464_);
  or (_02468_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand (_02469_, pc_log_change, _02437_);
  and (_02470_, _02469_, _06071_);
  and (_01734_, _02470_, _02468_);
  and (_02471_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  not (_02472_, pc_log_change);
  and (_02473_, _02472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or (_02474_, _02473_, _02471_);
  and (_01736_, _02474_, _06071_);
  nor (_02475_, _06359_, _02091_);
  not (_02476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_02477_, _06065_, _02476_);
  and (_02478_, _06059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_02479_, _02478_, _06547_);
  not (_02480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_02481_, _02220_, _02480_);
  nor (_02482_, _02481_, _02184_);
  or (_02483_, _02482_, _06065_);
  or (_02484_, _02483_, _02479_);
  and (_02485_, _02484_, _02477_);
  and (_02486_, _02485_, _06036_);
  and (_02487_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_02488_, _02487_, _02486_);
  or (_02489_, _02488_, _02475_);
  and (_01739_, _02489_, _06071_);
  and (_02491_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_02492_, _02472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or (_02493_, _02492_, _02491_);
  and (_01743_, _02493_, _06071_);
  and (_01763_, _07515_, _06071_);
  or (_02494_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_02495_, _06530_, _05754_);
  and (_02496_, _02495_, _06071_);
  and (_01816_, _02496_, _02494_);
  nor (_01829_, _11549_, rst);
  and (_02497_, _09349_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_02498_, _09341_, _06400_);
  and (_02500_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_02501_, _02500_, _09345_);
  or (_02502_, _02501_, _02498_);
  or (_02503_, _02502_, _02497_);
  and (_01835_, _02503_, _06071_);
  and (_01851_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and (_02504_, _09583_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02505_, _09003_, _09579_);
  and (_02507_, _02505_, _09005_);
  or (_02508_, _02507_, _02504_);
  and (_01870_, _02508_, _06071_);
  and (_02509_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_02510_, _11023_, _07979_);
  and (_02511_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_02512_, _02511_, _07983_);
  or (_02513_, _02512_, _02510_);
  or (_02514_, _02513_, _02509_);
  and (_01902_, _02514_, _06071_);
  and (_02515_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_02516_, _08865_, _06993_);
  or (_02517_, _02516_, _02515_);
  and (_01914_, _02517_, _06071_);
  nor (_02518_, _07011_, rst);
  or (_02519_, _06528_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_04199_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06071_);
  and (_02520_, _04199_, _02519_);
  or (_02025_, _02520_, _02518_);
  and (_02521_, _09576_, _06375_);
  nand (_02522_, _06375_, _06011_);
  and (_02523_, _02522_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_02524_, _02523_, _02521_);
  and (_02041_, _02524_, _06071_);
  nor (_02525_, _07945_, _06996_);
  and (_02526_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_02527_, _02526_, _06390_);
  or (_02528_, _02527_, _02525_);
  or (_02529_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_02530_, _02529_, _06071_);
  and (_02074_, _02530_, _02528_);
  and (_02531_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_02532_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_02533_, _02532_, _02531_);
  and (_02080_, _02533_, _06071_);
  nand (_02534_, _11791_, _07759_);
  or (_02535_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_02536_, _02535_, _06071_);
  and (_02094_, _02536_, _02534_);
  or (_02538_, _07757_, _07425_);
  or (_02539_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_02540_, _02539_, _06071_);
  and (_02099_, _02540_, _02538_);
  nor (_02541_, _11791_, _07107_);
  and (_02542_, _07107_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_02543_, _02542_, _07429_);
  or (_02544_, _02543_, _02541_);
  nand (_02546_, _12466_, _07429_);
  and (_02548_, _02546_, _06071_);
  and (_02104_, _02548_, _02544_);
  and (_02274_, _10978_, _06071_);
  and (_03772_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06071_);
  and (_02550_, _03772_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_02149_, _02550_, _02274_);
  and (_02552_, _08865_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_02553_, _08865_, _06359_);
  or (_02554_, _02553_, _02552_);
  and (_02175_, _02554_, _06071_);
  and (_02556_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_02197_, _02556_, _08597_);
  nor (_02239_, _11671_, rst);
  nand (_02557_, _07946_, _06993_);
  or (_02558_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_02560_, _02558_, _06071_);
  and (_02255_, _02560_, _02557_);
  not (_02562_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_02563_, _02562_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_02261_, _02563_, _06071_);
  and (_02564_, _13711_, _06032_);
  or (_02565_, _02564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_02566_, _02565_, _00557_);
  nand (_02567_, _02564_, _06803_);
  and (_02568_, _02567_, _02566_);
  nor (_02569_, _00557_, _06609_);
  or (_02570_, _02569_, _02568_);
  and (_02398_, _02570_, _06071_);
  and (_02571_, _13711_, _08801_);
  and (_02572_, _02571_, _06803_);
  nor (_02573_, _02571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_02574_, _02573_, _02572_);
  nand (_02575_, _02574_, _00557_);
  nand (_02576_, _13718_, _09341_);
  and (_02577_, _02576_, _06071_);
  and (_02400_, _02577_, _02575_);
  nand (_02578_, _11825_, _06071_);
  nor (_02427_, _02578_, _11933_);
  and (_02579_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_02466_, _02579_, _08588_);
  and (_02490_, _07848_, _06071_);
  and (_02580_, _06611_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02581_, _09576_, _06385_);
  or (_02582_, _02581_, _02580_);
  and (_02499_, _02582_, _06071_);
  and (_02506_, _07003_, _06508_);
  and (_02537_, _00268_, _06071_);
  nor (_02583_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_02584_, _11471_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02585_, _02584_, _02583_);
  nand (_02586_, _02585_, _00472_);
  nand (_02587_, _02586_, _06086_);
  or (_02588_, _02586_, _06086_);
  and (_02589_, _02588_, _02587_);
  and (_02590_, _02589_, _11751_);
  and (_02591_, _11827_, _07819_);
  and (_02592_, _11748_, _07870_);
  nor (_02593_, _00482_, _06086_);
  and (_02594_, _00482_, _06086_);
  or (_02595_, _02594_, _02593_);
  and (_02596_, _02595_, _12469_);
  and (_02597_, _12080_, _11424_);
  or (_02598_, _02597_, _02596_);
  and (_02599_, _12485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_02600_, _02599_, _02598_);
  nor (_02601_, _02600_, _02592_);
  nand (_02602_, _02601_, _12437_);
  or (_02603_, _02602_, _02591_);
  or (_02604_, _02603_, _02590_);
  and (_02605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_02606_, _02605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_02607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_02608_, _02607_, _12502_);
  and (_02609_, _02608_, _02606_);
  and (_02610_, _02609_, _12500_);
  or (_02611_, _02610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_02612_, _02610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_02613_, _02612_, _02611_);
  or (_02614_, _02613_, _12437_);
  and (_02615_, _02614_, _06071_);
  and (_02545_, _02615_, _02604_);
  and (_02616_, _05764_, _05722_);
  and (_02617_, _02616_, _05875_);
  nor (_02618_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_02619_, _02618_, _08705_);
  and (_02620_, _02619_, _05805_);
  and (_02621_, _05786_, _05743_);
  and (_02622_, _02621_, _02620_);
  and (_02623_, _05843_, _05825_);
  and (_02624_, _02623_, _02622_);
  and (_02547_, _02624_, _02617_);
  and (_02625_, _10959_, _06006_);
  or (_02626_, _02625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_02627_, _02626_, _09250_);
  nand (_02628_, _02625_, _06803_);
  and (_02629_, _02628_, _02627_);
  nor (_02630_, _09250_, _06993_);
  or (_02631_, _02630_, _02629_);
  and (_02549_, _02631_, _06071_);
  and (_02632_, _01609_, _06362_);
  or (_02633_, _02632_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_02634_, _02633_, _01623_);
  nand (_02635_, _02632_, _06803_);
  and (_02636_, _02635_, _02634_);
  nor (_02637_, _01623_, _09037_);
  or (_02638_, _02637_, _02636_);
  and (_02551_, _02638_, _06071_);
  and (_02639_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_02555_, _02639_, _07989_);
  and (_02640_, _10972_, rxd_i);
  not (_02641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nor (_02642_, _10972_, _02641_);
  or (_02643_, _02642_, _02640_);
  and (_02559_, _02643_, _06071_);
  or (_02644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_02645_, _02644_, _01891_);
  not (_02646_, _06805_);
  nor (_02647_, _02646_, _06803_);
  nand (_02648_, _02646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_02649_, _02648_, _01891_);
  or (_02650_, _02649_, _02647_);
  and (_02651_, _02650_, _02645_);
  or (_02652_, _02651_, _01898_);
  nand (_02653_, _01898_, _06359_);
  and (_02654_, _02653_, _06071_);
  and (_02561_, _02654_, _02652_);
  nand (_02655_, _13723_, _06359_);
  or (_02656_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_02657_, _02656_, _06071_);
  and (_02665_, _02657_, _02655_);
  and (_02658_, _13782_, _13731_);
  and (_02659_, _13784_, _13736_);
  and (_02660_, _02659_, _13780_);
  and (_02661_, _02660_, _13777_);
  nand (_02662_, _02661_, _13732_);
  nand (_02663_, _02662_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02664_, _02663_, _02658_);
  or (_02666_, _02664_, _13744_);
  and (_02673_, _02666_, _06071_);
  and (_02667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02668_, _07875_, _01916_);
  or (_02669_, _02668_, _07879_);
  nor (_02670_, _02669_, _02667_);
  or (_02671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_02672_, _02671_, _06071_);
  nor (_02674_, _02672_, _02670_);
  nor (_02688_, _11453_, rst);
  nor (_02675_, _13736_, _00436_);
  or (_02676_, _02675_, _02661_);
  and (_02677_, _02676_, _13733_);
  nand (_02678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_02679_, _02678_, _13732_);
  or (_02680_, _02679_, _02677_);
  and (_02681_, _02680_, _13765_);
  or (_02682_, _02681_, _02658_);
  and (_02707_, _02682_, _13798_);
  or (_02683_, _01691_, _01632_);
  and (_02684_, _02683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_02685_, _02684_, _10952_);
  and (_02686_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_02687_, _02686_, _00275_);
  and (_02689_, _02687_, _10948_);
  or (_02690_, _02689_, _02685_);
  nand (_02691_, _10952_, _06434_);
  and (_02692_, _02691_, _06071_);
  and (_02737_, _02692_, _02690_);
  and (_02693_, _01609_, _06383_);
  or (_02694_, _02693_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_02695_, _02694_, _01623_);
  nand (_02696_, _02693_, _06803_);
  and (_02697_, _02696_, _02695_);
  and (_02698_, _01608_, _07978_);
  or (_02699_, _02698_, _02697_);
  and (_02741_, _02699_, _06071_);
  and (_02700_, _01609_, _06032_);
  or (_02701_, _02700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_02702_, _02701_, _01623_);
  nand (_02703_, _02700_, _06803_);
  and (_02704_, _02703_, _02702_);
  nor (_02705_, _01623_, _06609_);
  or (_02706_, _02705_, _02704_);
  and (_02752_, _02706_, _06071_);
  nor (_02708_, _07912_, _07951_);
  or (_02709_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_02710_, _02709_, _07896_);
  or (_02711_, _02710_, _07887_);
  and (_02712_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_02713_, _02712_, rxd_i);
  and (_02714_, _02713_, _02711_);
  or (_02715_, _02714_, _02708_);
  nand (_02716_, _07887_, _09002_);
  and (_02717_, _02716_, _06560_);
  and (_02718_, _02717_, _02715_);
  and (_02719_, _06558_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02754_, _02719_, _02718_);
  and (_02720_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_02765_, _02720_, _07950_);
  nor (_02721_, _02670_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_02722_, _02721_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_02723_, _02721_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_02724_, _02723_, _06071_);
  and (_02769_, _02724_, _02722_);
  and (_02725_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02726_, _02725_, _13798_);
  and (_02727_, _13752_, _06071_);
  and (_02728_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02780_, _02728_, _02726_);
  nand (_02729_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_02730_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02731_, _02730_, _02729_);
  and (_02782_, _02731_, _13798_);
  and (_02732_, _13711_, _06805_);
  or (_02733_, _02732_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02734_, _02733_, _00557_);
  nand (_02735_, _02732_, _06803_);
  and (_02736_, _02735_, _02734_);
  nor (_02738_, _00557_, _06359_);
  or (_02739_, _02738_, _02736_);
  and (_02786_, _02739_, _06071_);
  and (_02740_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_02742_, _06530_, _05789_);
  or (_02743_, _02742_, _02740_);
  and (_02792_, _02743_, _06071_);
  nor (_02744_, _06496_, _06490_);
  or (_02745_, _06494_, _06483_);
  and (_02746_, _06481_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_02747_, _02746_, _02745_);
  and (_02748_, _02747_, _02744_);
  and (_02749_, _02748_, _01192_);
  or (_02750_, _06470_, _06457_);
  and (_02751_, _06468_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_02753_, _02751_, _02750_);
  and (_02755_, _02753_, _01176_);
  and (_02756_, _02755_, _01482_);
  or (_02757_, _02756_, _06508_);
  or (_02758_, _02757_, _02749_);
  or (_02759_, _06509_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_02760_, _02759_, _06071_);
  and (_02794_, _02760_, _02758_);
  nand (_02761_, _01192_, _06511_);
  and (_02762_, _06511_, _06474_);
  or (_02763_, _02762_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_02764_, _02763_, _06071_);
  and (_02810_, _02764_, _02761_);
  nand (_02766_, _00727_, _01192_);
  and (_02767_, _00727_, _06474_);
  or (_02768_, _02767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_02770_, _02768_, _06071_);
  and (_02813_, _02770_, _02766_);
  and (_02771_, _10959_, _07754_);
  or (_02772_, _02771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_02773_, _02772_, _09250_);
  nand (_02774_, _02771_, _06803_);
  and (_02775_, _02774_, _02773_);
  nor (_02776_, _09250_, _06434_);
  or (_02777_, _02776_, _02775_);
  and (_02825_, _02777_, _06071_);
  and (_02778_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_02779_, _06530_, _05773_);
  or (_02781_, _02779_, _02778_);
  and (_02874_, _02781_, _06071_);
  and (_02783_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_02784_, _06530_, _05835_);
  or (_02785_, _02784_, _02783_);
  and (_02895_, _02785_, _06071_);
  and (_02787_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_02788_, _06530_, _05817_);
  or (_02789_, _02788_, _02787_);
  and (_02908_, _02789_, _06071_);
  nor (_02980_, _11904_, rst);
  or (_02983_, _08776_, _08770_);
  and (_03013_, _08032_, _06071_);
  nor (_02790_, _13733_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02791_, _02790_, _13792_);
  and (_03057_, _02791_, _13798_);
  and (_02793_, _10943_, _06833_);
  and (_02795_, _02793_, _06032_);
  nand (_02796_, _02795_, _06803_);
  or (_02797_, _02795_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_02798_, _02797_, _06815_);
  and (_02799_, _02798_, _02796_);
  and (_02800_, _10951_, _06372_);
  not (_02801_, _02800_);
  nor (_02802_, _02801_, _06609_);
  not (_02803_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_02804_, _02800_, _02803_);
  or (_02805_, _02804_, _02802_);
  and (_02806_, _02805_, _06012_);
  nor (_02807_, _06814_, _02803_);
  or (_02808_, _02807_, rst);
  or (_02809_, _02808_, _02806_);
  or (_03119_, _02809_, _02799_);
  and (_02811_, _06810_, _08801_);
  nand (_02812_, _02811_, _06803_);
  or (_02814_, _02811_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02815_, _02814_, _06815_);
  and (_02816_, _02815_, _02812_);
  nand (_02817_, _09341_, _06822_);
  or (_02818_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02819_, _02818_, _06012_);
  and (_02820_, _02819_, _02817_);
  not (_02821_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_02822_, _06814_, _02821_);
  or (_02823_, _02822_, rst);
  or (_02824_, _02823_, _02820_);
  or (_03122_, _02824_, _02816_);
  and (_02826_, _06810_, _06362_);
  nand (_02827_, _02826_, _06803_);
  or (_02828_, _02826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02829_, _02828_, _06815_);
  and (_02830_, _02829_, _02827_);
  nand (_02831_, _09037_, _06822_);
  or (_02832_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02833_, _02832_, _06012_);
  and (_02834_, _02833_, _02831_);
  and (_02835_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_02836_, _02835_, rst);
  or (_02837_, _02836_, _02834_);
  or (_03124_, _02837_, _02830_);
  not (_02838_, _06834_);
  or (_02839_, _02838_, _01632_);
  and (_02840_, _02839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02841_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02842_, _02841_, _00275_);
  and (_02843_, _02842_, _06834_);
  or (_02844_, _02843_, _02840_);
  and (_02845_, _02844_, _06815_);
  nand (_02846_, _06841_, _06434_);
  or (_02847_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02848_, _02847_, _06012_);
  and (_02849_, _02848_, _02846_);
  and (_02850_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02851_, _02850_, rst);
  or (_02852_, _02851_, _02849_);
  or (_03127_, _02852_, _02845_);
  nor (_03136_, _11469_, rst);
  and (_02853_, _10943_, _06809_);
  and (_02854_, _02853_, _06006_);
  nand (_02855_, _02854_, _06803_);
  or (_02856_, _02854_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02857_, _02856_, _06815_);
  and (_02858_, _02857_, _02855_);
  and (_02859_, _01607_, _06372_);
  not (_02860_, _02859_);
  nor (_02861_, _02860_, _06993_);
  not (_02862_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_02863_, _02859_, _02862_);
  or (_02864_, _02863_, _02861_);
  and (_02865_, _02864_, _06012_);
  nor (_02866_, _06814_, _02862_);
  or (_02867_, _02866_, rst);
  or (_02868_, _02867_, _02865_);
  or (_03146_, _02868_, _02858_);
  and (_02869_, _02793_, _06006_);
  nand (_02870_, _02869_, _06803_);
  or (_02871_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_02872_, _02871_, _06815_);
  and (_02873_, _02872_, _02870_);
  nor (_02875_, _02801_, _06993_);
  not (_02876_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_02877_, _02800_, _02876_);
  or (_02878_, _02877_, _02875_);
  and (_02879_, _02878_, _06012_);
  nor (_02880_, _06814_, _02876_);
  or (_02881_, _02880_, rst);
  or (_02882_, _02881_, _02879_);
  or (_03148_, _02882_, _02873_);
  and (_02883_, _06810_, _06032_);
  nand (_02884_, _02883_, _06803_);
  or (_02885_, _02883_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02886_, _02885_, _06815_);
  and (_02887_, _02886_, _02884_);
  nand (_02888_, _06822_, _06609_);
  or (_02889_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02890_, _02889_, _06012_);
  and (_02891_, _02890_, _02888_);
  not (_02892_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_02893_, _06814_, _02892_);
  or (_02894_, _02893_, rst);
  or (_02896_, _02894_, _02891_);
  or (_03151_, _02896_, _02887_);
  and (_02897_, _06810_, _06383_);
  nand (_02898_, _02897_, _06803_);
  or (_02899_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_02900_, _02899_, _06815_);
  and (_02901_, _02900_, _02898_);
  nand (_02902_, _07977_, _06822_);
  and (_02903_, _02902_, _06012_);
  and (_02904_, _02903_, _02899_);
  nor (_02905_, _06814_, _00227_);
  or (_02906_, _02905_, rst);
  or (_02907_, _02906_, _02904_);
  or (_03153_, _02907_, _02901_);
  and (_02909_, _06810_, _07105_);
  nand (_02910_, _02909_, _06803_);
  or (_02911_, _02909_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02912_, _02911_, _06815_);
  and (_02913_, _02912_, _02910_);
  nand (_02914_, _07945_, _06822_);
  or (_02915_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02916_, _02915_, _06012_);
  and (_02917_, _02916_, _02914_);
  nor (_02918_, _06814_, _00003_);
  or (_02919_, _02918_, rst);
  or (_02920_, _02919_, _02917_);
  or (_03155_, _02920_, _02913_);
  and (_02921_, _06834_, _08801_);
  nand (_02922_, _02921_, _06803_);
  or (_02923_, _02921_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02924_, _02923_, _06815_);
  and (_02925_, _02924_, _02922_);
  nand (_02926_, _09341_, _06841_);
  or (_02927_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02928_, _02927_, _06012_);
  and (_02929_, _02928_, _02926_);
  not (_02930_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_02931_, _06814_, _02930_);
  or (_02932_, _02931_, rst);
  or (_02933_, _02932_, _02929_);
  or (_03157_, _02933_, _02925_);
  and (_02934_, _06840_, _06363_);
  nand (_02935_, _02934_, _06803_);
  or (_02936_, _02934_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02937_, _02936_, _06815_);
  and (_02938_, _02937_, _02935_);
  nand (_02939_, _09037_, _06841_);
  or (_02940_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02941_, _02940_, _06012_);
  and (_02942_, _02941_, _02939_);
  and (_02943_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_02944_, _02943_, rst);
  or (_02945_, _02944_, _02942_);
  or (_03159_, _02945_, _02938_);
  and (_02946_, _06834_, _06006_);
  nand (_02947_, _02946_, _06803_);
  or (_02948_, _02946_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02949_, _02948_, _06815_);
  and (_02950_, _02949_, _02947_);
  nand (_02951_, _06993_, _06841_);
  or (_02952_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02953_, _02952_, _06012_);
  and (_02954_, _02953_, _02951_);
  not (_02955_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_02956_, _06814_, _02955_);
  or (_02957_, _02956_, rst);
  or (_02958_, _02957_, _02954_);
  or (_03162_, _02958_, _02950_);
  and (_02959_, _02793_, _07105_);
  nand (_02960_, _02959_, _06803_);
  or (_02961_, _02959_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_02962_, _02961_, _06815_);
  and (_02963_, _02962_, _02960_);
  nor (_02964_, _02801_, _07945_);
  nor (_02965_, _02800_, _13994_);
  or (_02966_, _02965_, _02964_);
  and (_02967_, _02966_, _06012_);
  nor (_02968_, _06814_, _13994_);
  or (_02969_, _02968_, rst);
  or (_02970_, _02969_, _02967_);
  or (_03245_, _02970_, _02963_);
  and (_02971_, _02793_, _07754_);
  nand (_02972_, _02971_, _06803_);
  or (_02973_, _02971_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02974_, _02973_, _06815_);
  and (_02975_, _02974_, _02972_);
  nor (_02976_, _02801_, _06434_);
  and (_02977_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02978_, _02977_, _02976_);
  and (_02979_, _02978_, _06012_);
  and (_02981_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02982_, _02981_, rst);
  or (_02984_, _02982_, _02979_);
  or (_03246_, _02984_, _02975_);
  and (_02985_, _02793_, _06362_);
  nand (_02986_, _02985_, _06803_);
  or (_02987_, _02985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_02988_, _02987_, _06815_);
  and (_02989_, _02988_, _02986_);
  nor (_02990_, _02801_, _09037_);
  and (_02991_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02992_, _02991_, _02990_);
  and (_02993_, _02992_, _06012_);
  and (_02994_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_02995_, _02994_, rst);
  or (_02996_, _02995_, _02993_);
  or (_03261_, _02996_, _02989_);
  and (_02997_, _02853_, _07754_);
  nand (_02998_, _02997_, _06803_);
  or (_02999_, _02997_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_03000_, _02999_, _06815_);
  and (_03001_, _03000_, _02998_);
  nor (_03002_, _02860_, _06434_);
  and (_03003_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_03004_, _03003_, _03002_);
  and (_03005_, _03004_, _06012_);
  and (_03006_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_03007_, _03006_, rst);
  or (_03008_, _03007_, _03005_);
  or (_03263_, _03008_, _03001_);
  and (_03009_, _02853_, _06362_);
  nand (_03010_, _03009_, _06803_);
  or (_03011_, _03009_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_03012_, _03011_, _06815_);
  and (_03014_, _03012_, _03010_);
  nor (_03015_, _02860_, _09037_);
  and (_03016_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_03017_, _03016_, _03015_);
  and (_03018_, _03017_, _06012_);
  and (_03019_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_03020_, _03019_, rst);
  or (_03021_, _03020_, _03018_);
  or (_03264_, _03021_, _03014_);
  and (_03022_, _02853_, _08801_);
  nand (_03023_, _03022_, _06803_);
  or (_03024_, _03022_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03025_, _03024_, _06815_);
  and (_03026_, _03025_, _03023_);
  nor (_03027_, _02860_, _09341_);
  not (_03028_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_03029_, _02859_, _03028_);
  or (_03030_, _03029_, _03027_);
  and (_03031_, _03030_, _06012_);
  nor (_03032_, _06814_, _03028_);
  or (_03033_, _03032_, rst);
  or (_03034_, _03033_, _03031_);
  or (_03270_, _03034_, _03026_);
  and (_03035_, _06834_, _06383_);
  nand (_03036_, _03035_, _06803_);
  or (_03037_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_03038_, _03037_, _06815_);
  and (_03039_, _03038_, _03036_);
  nand (_03040_, _07977_, _06841_);
  and (_03041_, _03037_, _06012_);
  and (_03042_, _03041_, _03040_);
  nor (_03043_, _06814_, _00222_);
  or (_03044_, _03043_, rst);
  or (_03045_, _03044_, _03042_);
  or (_03285_, _03045_, _03039_);
  and (_03046_, _06834_, _06032_);
  nand (_03047_, _03046_, _06803_);
  or (_03048_, _03046_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03049_, _03048_, _06815_);
  and (_03050_, _03049_, _03047_);
  nand (_03051_, _06841_, _06609_);
  or (_03052_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03053_, _03052_, _06012_);
  and (_03054_, _03053_, _03051_);
  not (_03055_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_03056_, _06814_, _03055_);
  or (_03058_, _03056_, rst);
  or (_03059_, _03058_, _03054_);
  or (_03287_, _03059_, _03050_);
  and (_03060_, _06834_, _07105_);
  nand (_03061_, _03060_, _06803_);
  or (_03062_, _03060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03063_, _03062_, _06815_);
  and (_03064_, _03063_, _03061_);
  nand (_03065_, _07945_, _06841_);
  or (_03066_, _06841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03067_, _03066_, _06012_);
  and (_03068_, _03067_, _03065_);
  nor (_03069_, _06814_, _14003_);
  or (_03070_, _03069_, rst);
  or (_03071_, _03070_, _03068_);
  or (_03289_, _03071_, _03064_);
  and (_03072_, _02793_, _06383_);
  nand (_03073_, _03072_, _06803_);
  or (_03074_, _03072_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_03075_, _03074_, _06815_);
  and (_03076_, _03075_, _03073_);
  and (_03077_, _02800_, _07978_);
  nor (_03078_, _02800_, _00211_);
  or (_03079_, _03078_, _03077_);
  and (_03080_, _03079_, _06012_);
  nor (_03081_, _06814_, _00211_);
  or (_03082_, _03081_, rst);
  or (_03083_, _03082_, _03080_);
  or (_03291_, _03083_, _03076_);
  and (_03084_, _06810_, _06006_);
  nand (_03085_, _03084_, _06803_);
  or (_03086_, _03084_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03087_, _03086_, _06815_);
  and (_03088_, _03087_, _03085_);
  nand (_03089_, _06993_, _06822_);
  or (_03090_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03091_, _03090_, _06012_);
  and (_03092_, _03091_, _03089_);
  not (_03093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_03094_, _06814_, _03093_);
  or (_03095_, _03094_, rst);
  or (_03096_, _03095_, _03092_);
  or (_03294_, _03096_, _03088_);
  and (_03097_, _06810_, _07754_);
  nand (_03098_, _03097_, _06803_);
  or (_03099_, _03097_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03100_, _03099_, _06815_);
  and (_03101_, _03100_, _03098_);
  nand (_03102_, _06822_, _06434_);
  or (_03103_, _06822_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03104_, _03103_, _06012_);
  and (_03105_, _03104_, _03102_);
  and (_03106_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_03107_, _03106_, rst);
  or (_03108_, _03107_, _03105_);
  or (_03296_, _03108_, _03101_);
  nand (_03109_, _02859_, _06803_);
  or (_03110_, _02859_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_03111_, _03110_, _06815_);
  and (_03112_, _03111_, _03109_);
  nand (_03113_, _02859_, _07977_);
  and (_03114_, _03113_, _06012_);
  and (_03115_, _03114_, _03110_);
  nor (_03116_, _06814_, _00216_);
  or (_03117_, _03116_, rst);
  or (_03118_, _03117_, _03115_);
  or (_03298_, _03118_, _03112_);
  and (_03120_, _02793_, _08801_);
  nand (_03121_, _03120_, _06803_);
  or (_03123_, _03120_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_03125_, _03123_, _06815_);
  and (_03126_, _03125_, _03121_);
  nor (_03128_, _02801_, _09341_);
  not (_03129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_03130_, _02800_, _03129_);
  or (_03131_, _03130_, _03128_);
  and (_03132_, _03131_, _06012_);
  nor (_03133_, _06814_, _03129_);
  or (_03134_, _03133_, rst);
  or (_03135_, _03134_, _03132_);
  or (_03300_, _03135_, _03126_);
  and (_03137_, _02853_, _06032_);
  nand (_03138_, _03137_, _06803_);
  or (_03139_, _03137_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_03140_, _03139_, _06815_);
  and (_03141_, _03140_, _03138_);
  nor (_03142_, _02860_, _06609_);
  not (_03143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_03144_, _02859_, _03143_);
  or (_03145_, _03144_, _03142_);
  and (_03147_, _03145_, _06012_);
  nor (_03149_, _06814_, _03143_);
  or (_03150_, _03149_, rst);
  or (_03152_, _03150_, _03147_);
  or (_03303_, _03152_, _03141_);
  and (_03154_, _02853_, _07105_);
  nand (_03156_, _03154_, _06803_);
  or (_03158_, _03154_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03160_, _03158_, _06815_);
  and (_03161_, _03160_, _03156_);
  nor (_03163_, _02860_, _07945_);
  nor (_03164_, _02859_, _13986_);
  or (_03165_, _03164_, _03163_);
  and (_03166_, _03165_, _06012_);
  nor (_03167_, _06814_, _13986_);
  or (_03168_, _03167_, rst);
  or (_03169_, _03168_, _03166_);
  or (_03305_, _03169_, _03161_);
  nor (_03170_, _09037_, _06996_);
  and (_03171_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03172_, _03171_, _06390_);
  or (_03173_, _03172_, _03170_);
  or (_03174_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03175_, _03174_, _06071_);
  and (_03317_, _03175_, _03173_);
  or (_03176_, _08065_, _08032_);
  nor (_03177_, _03176_, _07103_);
  nand (_03178_, _03177_, _07751_);
  or (_03179_, _03178_, _07609_);
  or (_03180_, _03179_, _07365_);
  and (_03181_, _03180_, _07344_);
  or (_03182_, _06712_, _06710_);
  not (_03183_, _06618_);
  nand (_03184_, _06710_, _03183_);
  and (_03185_, _03184_, _06615_);
  and (_03186_, _03185_, _03182_);
  nand (_03187_, _06747_, _06717_);
  and (_03188_, _06748_, _06715_);
  and (_03189_, _03188_, _03187_);
  and (_03190_, _07454_, _07109_);
  and (_03191_, _03190_, _07449_);
  nand (_03192_, _03191_, _07108_);
  nand (_03193_, _03192_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_03194_, _03193_, _03189_);
  nor (_03195_, _03194_, _03186_);
  and (_03196_, _03195_, _07684_);
  nand (_03197_, _03196_, _07788_);
  or (_03198_, _03197_, _03181_);
  nor (_03199_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_03200_, _03199_, _10896_);
  and (_03201_, _03200_, _03198_);
  and (_03202_, _00274_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03203_, _03202_, _00275_);
  nand (_03204_, _03203_, _10896_);
  nand (_03205_, _03204_, _08985_);
  or (_03206_, _03205_, _03201_);
  nand (_03207_, _08988_, _06434_);
  and (_03208_, _03207_, _06071_);
  and (_03322_, _03208_, _03206_);
  nand (_03209_, _09037_, _07946_);
  or (_03210_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03211_, _03210_, _06071_);
  and (_03330_, _03211_, _03209_);
  nor (_03212_, _06967_, _06359_);
  and (_03213_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_03214_, _03213_, _03212_);
  and (_03344_, _03214_, _06071_);
  and (_03347_, _08065_, _06071_);
  and (_03215_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_03216_, _06530_, _05739_);
  or (_03217_, _03216_, _03215_);
  and (_03351_, _03217_, _06071_);
  and (_03218_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_03219_, _06530_, _05716_);
  or (_03220_, _03219_, _03218_);
  and (_03353_, _03220_, _06071_);
  or (_03221_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_03222_, _06530_, _05798_);
  and (_03223_, _03222_, _06071_);
  and (_03356_, _03223_, _03221_);
  and (_03224_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_03225_, _06530_, _05782_);
  or (_03226_, _03225_, _03224_);
  and (_03358_, _03226_, _06071_);
  nor (_03227_, _09341_, _06996_);
  and (_03228_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03229_, _03228_, _06390_);
  or (_03230_, _03229_, _03227_);
  or (_03231_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03232_, _03231_, _06071_);
  and (_03377_, _03232_, _03230_);
  and (_03233_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_03234_, _06530_, _05749_);
  or (_03235_, _03234_, _03233_);
  and (_03424_, _03235_, _06071_);
  or (_03236_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_03237_, _06530_, _05865_);
  and (_03238_, _03237_, _06071_);
  and (_03431_, _03238_, _03236_);
  and (_03239_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_03240_, _06530_, _05737_);
  or (_03241_, _03240_, _03239_);
  and (_03440_, _03241_, _06071_);
  or (_03242_, _09583_, _07893_);
  or (_03243_, _09005_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_03244_, _03243_, _06071_);
  and (_03444_, _03244_, _03242_);
  and (_03450_, _07741_, _06071_);
  and (_03247_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_03248_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_03249_, _03248_, _03247_);
  and (_03472_, _03249_, _06071_);
  and (_03250_, _11273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_03251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_03252_, _11290_, _03251_);
  and (_03253_, _11290_, _03251_);
  nor (_03254_, _03253_, _03252_);
  and (_03255_, _03254_, _11297_);
  nor (_03256_, _03254_, _11297_);
  or (_03257_, _03256_, _03255_);
  or (_03258_, _03257_, _09711_);
  or (_03259_, _09710_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03260_, _03259_, _11270_);
  and (_03262_, _03260_, _03258_);
  or (_03479_, _03262_, _03250_);
  nor (_03481_, _12052_, rst);
  nor (_03265_, _06530_, _06528_);
  nor (_03266_, _11370_, _11367_);
  nor (_03267_, _03266_, _06528_);
  and (_03268_, _03267_, _05694_);
  nor (_03269_, _03267_, _05694_);
  nor (_03271_, _03269_, _03268_);
  nor (_03272_, _03271_, _03265_);
  and (_03273_, _05699_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_03274_, _03273_, _03265_);
  nor (_03275_, _03274_, _11234_);
  or (_03276_, _03275_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_03277_, _03276_, _03272_);
  and (_03485_, _03277_, _06071_);
  or (_03278_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_03279_, _06530_, _05835_);
  and (_03280_, _03279_, _06071_);
  and (_03488_, _03280_, _03278_);
  and (_03499_, _07604_, _06071_);
  and (_03500_, _07680_, _06071_);
  nor (_03521_, _11763_, rst);
  or (_03281_, _01784_, _07564_);
  not (_03282_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_03283_, _01784_, _03282_);
  and (_03284_, _03283_, _06012_);
  and (_03286_, _03284_, _03281_);
  nor (_03288_, _06814_, _03282_);
  or (_03290_, _01791_, _01632_);
  and (_03292_, _03290_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_03293_, _06361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03295_, _03293_, _00275_);
  and (_03297_, _03295_, _01783_);
  or (_03299_, _03297_, _03292_);
  and (_03301_, _03299_, _06815_);
  or (_03302_, _03301_, _03288_);
  or (_03304_, _03302_, _03286_);
  and (_03554_, _03304_, _06071_);
  and (_03306_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_03307_, _06530_, _10690_);
  or (_03308_, _03307_, _03306_);
  and (_03563_, _03308_, _06071_);
  or (_03309_, _08535_, _05747_);
  or (_03310_, _06526_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_03311_, _03310_, _06071_);
  and (_03565_, _03311_, _03309_);
  and (_03312_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_03313_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nand (_03314_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_03315_, _03314_, _03313_);
  nand (_03316_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand (_03318_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_03319_, _03318_, _03316_);
  and (_03320_, _03319_, _03315_);
  nand (_03321_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand (_03323_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_03324_, _03323_, _03321_);
  nand (_03325_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand (_03326_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_03327_, _03326_, _03325_);
  and (_03328_, _03327_, _03324_);
  and (_03329_, _03328_, _03320_);
  nand (_03331_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand (_03332_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_03333_, _03332_, _03331_);
  nand (_03334_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_03335_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_03336_, _03335_, _03334_);
  and (_03337_, _03336_, _03333_);
  nand (_03338_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nand (_03339_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_03340_, _03339_, _03338_);
  nand (_03341_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_03342_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_03343_, _03342_, _03341_);
  and (_03345_, _03343_, _03340_);
  and (_03346_, _03345_, _03337_);
  and (_03348_, _03346_, _03329_);
  nand (_03349_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_03350_, _13897_, _12143_);
  and (_03352_, _03350_, _03349_);
  nand (_03354_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_03355_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_03357_, _03355_, _03354_);
  and (_03359_, _03357_, _03352_);
  nor (_03360_, _13983_, p1_in[5]);
  and (_03361_, _13983_, _02892_);
  nor (_03362_, _03361_, _03360_);
  nand (_03363_, _03362_, _14007_);
  nor (_03364_, _13983_, p0_in[5]);
  and (_03365_, _13983_, _03055_);
  nor (_03366_, _03365_, _03364_);
  nand (_03367_, _03366_, _14000_);
  and (_03368_, _03367_, _03363_);
  nor (_03369_, _13983_, p3_in[5]);
  and (_03370_, _13983_, _03143_);
  nor (_03371_, _03370_, _03369_);
  nand (_03372_, _03371_, _13966_);
  nor (_03373_, _13983_, p2_in[5]);
  and (_03374_, _13983_, _02803_);
  nor (_03375_, _03374_, _03373_);
  nand (_03376_, _03375_, _13991_);
  and (_03378_, _03376_, _03372_);
  and (_03379_, _03378_, _03368_);
  and (_03380_, _03379_, _03359_);
  nand (_03381_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_03382_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03383_, _03382_, _03381_);
  and (_03384_, _03383_, _03380_);
  nand (_03385_, _03384_, _03348_);
  nand (_03386_, _03385_, _13919_);
  nand (_03387_, _03386_, _13925_);
  or (_03388_, _03387_, _03312_);
  nand (_03389_, _13924_, _07643_);
  and (_03390_, _03389_, _06071_);
  and (_03570_, _03390_, _03388_);
  and (_03391_, _06967_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_03392_, _06967_, _06434_);
  or (_03393_, _03392_, _03391_);
  and (_03576_, _03393_, _06071_);
  or (_03394_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_03395_, _06530_, _05793_);
  and (_03396_, _03395_, _06071_);
  and (_03579_, _03396_, _03394_);
  and (_03585_, _07536_, _06071_);
  or (_03397_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_03398_, _06530_, _05732_);
  and (_03399_, _03398_, _06071_);
  and (_03587_, _03399_, _03397_);
  or (_03400_, _01784_, _00366_);
  not (_03401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_03402_, _01784_, _03401_);
  and (_03403_, _03402_, _06012_);
  and (_03404_, _03403_, _03400_);
  nor (_03405_, _06814_, _03401_);
  and (_03406_, _01783_, _06032_);
  nand (_03407_, _03406_, _06803_);
  or (_03408_, _03406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03409_, _03408_, _06815_);
  and (_03410_, _03409_, _03407_);
  or (_03411_, _03410_, _03405_);
  or (_03412_, _03411_, _03404_);
  and (_03592_, _03412_, _06071_);
  and (_03413_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_03414_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_03415_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_03416_, _03415_, _03414_);
  nand (_03417_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand (_03418_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_03419_, _03418_, _03417_);
  and (_03420_, _03419_, _03416_);
  nand (_03421_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand (_03422_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03423_, _03422_, _03421_);
  nand (_03425_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nand (_03426_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_03427_, _03426_, _03425_);
  and (_03428_, _03427_, _03423_);
  and (_03429_, _03428_, _03420_);
  nand (_03430_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand (_03432_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_03433_, _03432_, _03430_);
  nand (_03434_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_03435_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_03436_, _03435_, _03434_);
  and (_03437_, _03436_, _03433_);
  nand (_03438_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand (_03439_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_03441_, _03439_, _03438_);
  nand (_03442_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_03443_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_03445_, _03443_, _03442_);
  and (_03446_, _03445_, _03441_);
  and (_03447_, _03446_, _03437_);
  and (_03448_, _03447_, _03429_);
  nand (_03449_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_03451_, _13897_, _12100_);
  and (_03452_, _03451_, _03449_);
  nand (_03453_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand (_03454_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_03455_, _03454_, _03453_);
  and (_03456_, _03455_, _03452_);
  nor (_03457_, _13983_, p2_in[6]);
  and (_03458_, _13983_, _03129_);
  nor (_03459_, _03458_, _03457_);
  nand (_03460_, _03459_, _13991_);
  nor (_03461_, _13983_, p3_in[6]);
  and (_03462_, _13983_, _03028_);
  nor (_03463_, _03462_, _03461_);
  nand (_03464_, _03463_, _13966_);
  and (_03465_, _03464_, _03460_);
  nor (_03466_, _13983_, p0_in[6]);
  and (_03467_, _13983_, _02930_);
  nor (_03468_, _03467_, _03466_);
  nand (_03469_, _03468_, _14000_);
  nor (_03470_, _13983_, p1_in[6]);
  and (_03471_, _13983_, _02821_);
  nor (_03473_, _03471_, _03470_);
  nand (_03474_, _03473_, _14007_);
  and (_03475_, _03474_, _03469_);
  and (_03476_, _03475_, _03465_);
  and (_03477_, _03476_, _03456_);
  nand (_03478_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_03480_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_03482_, _03480_, _03478_);
  and (_03484_, _03482_, _03477_);
  nand (_03486_, _03484_, _03448_);
  nand (_03487_, _03486_, _13919_);
  nand (_03489_, _03487_, _13925_);
  or (_03490_, _03489_, _03413_);
  nand (_03491_, _13924_, _07426_);
  and (_03492_, _03491_, _06071_);
  and (_03614_, _03492_, _03490_);
  and (_03617_, _11935_, _06071_);
  or (_03493_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_03494_, _06530_, _05708_);
  and (_03495_, _03494_, _06071_);
  and (_03630_, _03495_, _03493_);
  and (_03639_, _08062_, _06071_);
  nor (_03645_, _12163_, rst);
  or (_03496_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_03497_, _06530_, _05791_);
  and (_03498_, _03497_, _06071_);
  and (_03650_, _03498_, _03496_);
  nor (_03652_, _12199_, rst);
  nor (_03669_, _12021_, rst);
  nand (_03671_, _12336_, _06071_);
  nor (_03678_, _12420_, rst);
  and (_03501_, _12524_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_03502_, _01721_, _11865_);
  and (_03503_, _11396_, _13379_);
  and (_03504_, _11874_, _11408_);
  and (_03505_, _11400_, _11396_);
  or (_03506_, _03505_, _03504_);
  or (_03507_, _03506_, _03503_);
  and (_03508_, _11404_, _11396_);
  or (_03509_, _03508_, _11859_);
  or (_03510_, _03509_, _03507_);
  or (_03511_, _03510_, _03502_);
  and (_03512_, _13639_, _11422_);
  or (_03513_, _03512_, _11837_);
  and (_03514_, _13379_, _08732_);
  and (_03515_, _03514_, _11412_);
  and (_03516_, _03514_, _11810_);
  or (_03517_, _03516_, _03515_);
  and (_03518_, _11401_, _08757_);
  and (_03519_, _11410_, _08757_);
  or (_03520_, _03519_, _03518_);
  or (_03522_, _03520_, _03517_);
  or (_03523_, _03522_, _03513_);
  and (_03524_, _11810_, _11410_);
  and (_03525_, _11415_, _11401_);
  or (_03526_, _03525_, _03524_);
  and (_03527_, _11404_, _08732_);
  and (_03528_, _03527_, _08757_);
  and (_03529_, _11414_, _08757_);
  or (_03530_, _03529_, _03528_);
  and (_03531_, _03514_, _11422_);
  and (_03532_, _11404_, _11391_);
  or (_03533_, _03532_, _03531_);
  or (_03534_, _03533_, _03530_);
  or (_03535_, _03534_, _03526_);
  or (_03536_, _11803_, _11413_);
  and (_03537_, _13632_, _11391_);
  and (_03538_, _11889_, _11408_);
  or (_03539_, _03538_, _13352_);
  or (_03540_, _03539_, _03537_);
  or (_03541_, _03540_, _03536_);
  and (_03542_, _11415_, _03527_);
  or (_03543_, _03542_, _03541_);
  or (_03544_, _03543_, _03535_);
  or (_03545_, _03544_, _03523_);
  or (_03546_, _03545_, _03511_);
  and (_03547_, _03546_, _08775_);
  or (_03682_, _03547_, _03501_);
  or (_03548_, _08535_, _05726_);
  or (_03549_, _06526_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_03550_, _03549_, _06071_);
  and (_03702_, _03550_, _03548_);
  and (_03551_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_03552_, _06530_, _06962_);
  or (_03553_, _03552_, _03551_);
  and (_03713_, _03553_, _06071_);
  and (_03555_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_03556_, _06530_, _06850_);
  or (_03557_, _03556_, _03555_);
  and (_03715_, _03557_, _06071_);
  and (_03558_, _06560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_03725_, _03558_, _08603_);
  and (_03559_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_03560_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_03561_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_03562_, _03561_, _03560_);
  nand (_03564_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand (_03566_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03567_, _03566_, _03564_);
  and (_03568_, _03567_, _03562_);
  nand (_03569_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_03571_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_03572_, _03571_, _03569_);
  nand (_03573_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_03574_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_03575_, _03574_, _03573_);
  and (_03577_, _03575_, _03572_);
  and (_03578_, _03577_, _03568_);
  nand (_03580_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand (_03581_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_03582_, _03581_, _03580_);
  nand (_03583_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand (_03584_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_03586_, _03584_, _03583_);
  and (_03588_, _03586_, _03582_);
  nand (_03589_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand (_03590_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_03591_, _03590_, _03589_);
  nand (_03593_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_03594_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_03595_, _03594_, _03593_);
  and (_03596_, _03595_, _03591_);
  and (_03597_, _03596_, _03588_);
  and (_03598_, _03597_, _03578_);
  nand (_03599_, _13897_, _12213_);
  nand (_03600_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03601_, _03600_, _03599_);
  nand (_03602_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_03603_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_03604_, _03603_, _03602_);
  and (_03605_, _03604_, _03601_);
  nor (_03606_, _13983_, p0_in[4]);
  and (_03607_, _13983_, _02955_);
  nor (_03608_, _03607_, _03606_);
  nand (_03609_, _03608_, _14000_);
  nor (_03610_, _13983_, p1_in[4]);
  and (_03611_, _13983_, _03093_);
  nor (_03612_, _03611_, _03610_);
  nand (_03613_, _03612_, _14007_);
  and (_03615_, _03613_, _03609_);
  nor (_03616_, _13983_, p3_in[4]);
  and (_03618_, _13983_, _02862_);
  nor (_03619_, _03618_, _03616_);
  nand (_03620_, _03619_, _13966_);
  nor (_03621_, _13983_, p2_in[4]);
  and (_03622_, _13983_, _02876_);
  nor (_03623_, _03622_, _03621_);
  nand (_03624_, _03623_, _13991_);
  and (_03625_, _03624_, _03620_);
  and (_03626_, _03625_, _03615_);
  and (_03627_, _03626_, _03605_);
  nand (_03628_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_03629_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03631_, _03629_, _03628_);
  and (_03632_, _03631_, _03627_);
  nand (_03633_, _03632_, _03598_);
  nand (_03634_, _03633_, _13919_);
  nand (_03635_, _03634_, _13925_);
  or (_03636_, _03635_, _03559_);
  nand (_03637_, _13924_, _07715_);
  and (_03638_, _03637_, _06071_);
  and (_03740_, _03638_, _03636_);
  or (_03640_, _13975_, _13625_);
  or (_03641_, _03640_, _01722_);
  not (_03642_, _11861_);
  and (_03643_, _08748_, _08732_);
  and (_03644_, _03643_, _11412_);
  or (_03646_, _03644_, _03642_);
  or (_03647_, _11885_, _11413_);
  or (_03648_, _11857_, _11847_);
  or (_03649_, _03648_, _03647_);
  or (_03651_, _03649_, _03646_);
  nand (_03653_, _11842_, _11835_);
  or (_03654_, _03653_, _03651_);
  or (_03655_, _03654_, _03641_);
  and (_03656_, _11889_, _08760_);
  or (_03657_, _03656_, _11917_);
  or (_03658_, _13627_, _11868_);
  or (_03659_, _03658_, _03657_);
  or (_03660_, _03659_, _03655_);
  and (_03661_, _03660_, _06527_);
  and (_03662_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03663_, _11403_, _11385_);
  or (_03664_, _03663_, _13643_);
  or (_03665_, _03664_, _03662_);
  or (_03666_, _03665_, _03661_);
  and (_03742_, _03666_, _06071_);
  and (_03667_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_03668_, _06530_, _06532_);
  or (_03670_, _03668_, _03667_);
  and (_03748_, _03670_, _06071_);
  and (_03672_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08003_);
  and (_03673_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03674_, _03673_, _03672_);
  and (_03752_, _03674_, _06071_);
  or (_03675_, _08535_, _05847_);
  or (_03676_, _06526_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_03677_, _03676_, _06071_);
  and (_03756_, _03677_, _03675_);
  nand (_03679_, _02311_, _06359_);
  and (_03680_, _02317_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_03681_, _02316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_03683_, _03681_, _03680_);
  or (_03684_, _03683_, _02311_);
  and (_03685_, _03684_, _06071_);
  and (_03780_, _03685_, _03679_);
  nand (_03686_, _07946_, _06609_);
  or (_03687_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03688_, _03687_, _06071_);
  and (_03813_, _03688_, _03686_);
  and (_03689_, _12524_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_03690_, _11840_, _08757_);
  or (_03691_, _03529_, _03524_);
  or (_03692_, _03691_, _03690_);
  and (_03693_, _11396_, _11388_);
  and (_03694_, _11391_, _11388_);
  or (_03695_, _03694_, _03693_);
  or (_03696_, _11876_, _03695_);
  or (_03697_, _03696_, _01721_);
  or (_03698_, _03697_, _03692_);
  and (_03699_, _13967_, _11387_);
  or (_03700_, _03699_, _11909_);
  or (_03701_, _03700_, _13360_);
  or (_03703_, _03701_, _13353_);
  or (_03704_, _11856_, _12548_);
  or (_03705_, _03528_, _03704_);
  or (_03706_, _03705_, _03703_);
  or (_03707_, _03706_, _03698_);
  or (_03708_, _03707_, _03523_);
  and (_03709_, _03708_, _08775_);
  or (_03822_, _03709_, _03689_);
  and (_03710_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03711_, _07979_, _12197_);
  and (_03712_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03714_, _03712_, _07983_);
  or (_03716_, _03714_, _03711_);
  or (_03717_, _03716_, _03710_);
  and (_03823_, _03717_, _06071_);
  and (_03718_, _13346_, _08732_);
  and (_03719_, _13360_, _08732_);
  or (_03720_, _13337_, _11811_);
  or (_03721_, _03720_, _08761_);
  or (_03722_, _03721_, _03719_);
  and (_03723_, _13360_, _08764_);
  or (_03724_, _12542_, _11908_);
  or (_03726_, _03724_, _13349_);
  or (_03727_, _03726_, _03723_);
  or (_03728_, _03727_, _03722_);
  or (_03729_, _03728_, _03718_);
  not (_03730_, _11836_);
  or (_03731_, _12533_, _03730_);
  and (_03732_, _11840_, _11415_);
  or (_03733_, _03524_, _11844_);
  nor (_03734_, _03733_, _03732_);
  nand (_03735_, _03734_, _11804_);
  or (_03736_, _11916_, _13978_);
  or (_03737_, _03736_, _03735_);
  or (_03738_, _03737_, _03731_);
  or (_03739_, _03738_, _03729_);
  and (_03741_, _03739_, _08775_);
  and (_03743_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_03744_, _11811_, _11744_);
  or (_03746_, _03744_, _03743_);
  and (_03747_, _03746_, _06071_);
  or (_03834_, _03747_, _03741_);
  and (_03749_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03750_, _07979_, _12019_);
  and (_03751_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03753_, _03751_, _07983_);
  or (_03754_, _03753_, _03750_);
  or (_03755_, _03754_, _03749_);
  and (_03837_, _03755_, _06071_);
  nand (_03757_, _07946_, _06359_);
  or (_03758_, _07946_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03759_, _03758_, _06071_);
  and (_03847_, _03759_, _03757_);
  and (_03760_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08003_);
  and (_03761_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03762_, _03761_, _03760_);
  and (_03853_, _03762_, _06071_);
  and (_03763_, _02793_, _06805_);
  nand (_03764_, _03763_, _06803_);
  or (_03765_, _03763_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03766_, _03765_, _06815_);
  and (_03767_, _03766_, _03764_);
  nor (_03768_, _02801_, _06359_);
  and (_03769_, _02801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_03770_, _03769_, _03768_);
  and (_03771_, _03770_, _06012_);
  and (_03773_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_03774_, _03773_, rst);
  or (_03775_, _03774_, _03771_);
  or (_03862_, _03775_, _03767_);
  and (_03776_, _02853_, _06805_);
  nand (_03777_, _03776_, _06803_);
  or (_03778_, _03776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03779_, _03778_, _06815_);
  and (_03781_, _03779_, _03777_);
  nor (_03782_, _02860_, _06359_);
  and (_03783_, _02860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_03784_, _03783_, _03782_);
  and (_03785_, _03784_, _06012_);
  and (_03786_, _06827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_03787_, _03786_, rst);
  or (_03788_, _03787_, _03785_);
  or (_03867_, _03788_, _03781_);
  and (_03880_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_03789_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  nand (_03790_, _06530_, _11005_);
  and (_03791_, _03790_, _06071_);
  and (_03889_, _03791_, _03789_);
  and (_03891_, _00283_, _06071_);
  and (_03792_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_03793_, _03792_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_03794_, _03792_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_03795_, _03794_, _03793_);
  and (_03897_, _03795_, _06071_);
  or (_03796_, _01784_, _07819_);
  not (_03797_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_03798_, _01784_, _03797_);
  and (_03799_, _03798_, _06012_);
  and (_03800_, _03799_, _03796_);
  nor (_03801_, _06814_, _03797_);
  and (_03802_, _01783_, _06805_);
  nand (_03803_, _03802_, _06803_);
  or (_03804_, _03802_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03805_, _03804_, _06815_);
  and (_03806_, _03805_, _03803_);
  or (_03807_, _03806_, _03801_);
  or (_03808_, _03807_, _03800_);
  and (_03903_, _03808_, _06071_);
  or (_03809_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_03810_, _06530_, _05817_);
  and (_03811_, _03810_, _06071_);
  and (_03907_, _03811_, _03809_);
  nor (_03812_, _02360_, _06359_);
  nor (_03814_, _02313_, _02476_);
  and (_03815_, _02313_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_03816_, _03815_, _03814_);
  nor (_03817_, _03816_, _02315_);
  or (_03818_, _03817_, _02323_);
  or (_03819_, _03818_, _03812_);
  nand (_03820_, _02323_, _02476_);
  and (_03821_, _03820_, _06071_);
  and (_03919_, _03821_, _03819_);
  nor (_03824_, _06996_, _06359_);
  and (_03825_, _06996_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03826_, _03825_, _06390_);
  or (_03827_, _03826_, _03824_);
  or (_03828_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03829_, _03828_, _06071_);
  and (_03924_, _03829_, _03827_);
  and (_03929_, _06071_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_03830_, _08535_, _05829_);
  or (_03831_, _06526_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_03832_, _03831_, _06071_);
  and (_03936_, _03832_, _03830_);
  and (_03833_, _07958_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03835_, _07979_, _12161_);
  and (_03836_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03838_, _03836_, _07983_);
  or (_03839_, _03838_, _03835_);
  or (_03840_, _03839_, _03833_);
  and (_03968_, _03840_, _06071_);
  or (_03841_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_03842_, _06530_, _05789_);
  and (_03843_, _03842_, _06071_);
  and (_04006_, _03843_, _03841_);
  and (_03844_, _06530_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_03845_, _12494_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_03846_, _03845_, _03844_);
  and (_04040_, _03846_, _06071_);
  or (_03848_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand (_03849_, _06530_, _09701_);
  and (_03850_, _03849_, _06071_);
  and (_04050_, _03850_, _03848_);
  and (_04054_, _00247_, _06071_);
  and (_03851_, _11097_, _05860_);
  and (_03852_, _11117_, _05849_);
  or (_03854_, _03852_, _11202_);
  or (_03855_, _03854_, _03851_);
  or (_03856_, _11178_, _05851_);
  or (_03857_, _03856_, _03855_);
  or (_03858_, _03857_, _11125_);
  nand (_03859_, _11138_, _11101_);
  nand (_03860_, _11231_, _03859_);
  and (_03861_, _11139_, _05850_);
  or (_03863_, _11117_, _11171_);
  and (_03864_, _03863_, _11101_);
  or (_03865_, _03864_, _03861_);
  or (_03866_, _03865_, _03860_);
  or (_03868_, _03866_, _05885_);
  nand (_03869_, _11136_, _11112_);
  or (_03870_, _03869_, _03868_);
  or (_03871_, _03870_, _03858_);
  and (_03872_, _03871_, _08705_);
  nor (_03873_, _05691_, _13383_);
  or (_03874_, _03873_, rst);
  or (_04056_, _03874_, _03872_);
  or (_03875_, _13340_, _11845_);
  and (_03876_, _11830_, _11391_);
  or (_03877_, _03876_, _13976_);
  or (_03878_, _03877_, _03875_);
  not (_03879_, _11910_);
  or (_03881_, _13344_, _03879_);
  or (_03882_, _03881_, _03878_);
  and (_03883_, _13354_, _11390_);
  or (_03884_, _03883_, _03732_);
  or (_03885_, _03884_, _12546_);
  or (_03886_, _03885_, _03882_);
  and (_03887_, _11884_, _11810_);
  or (_03888_, _03647_, _03887_);
  or (_03890_, _03888_, _03525_);
  or (_03892_, _12549_, _11416_);
  or (_03893_, _03892_, _03539_);
  and (_03894_, _11830_, _11396_);
  and (_03895_, _11414_, _08756_);
  or (_03896_, _03895_, _13335_);
  or (_03898_, _03896_, _03894_);
  nor (_03899_, _03898_, _03893_);
  nand (_03900_, _03899_, _13979_);
  or (_03901_, _03900_, _03890_);
  or (_03902_, _03901_, _03886_);
  and (_03904_, _03902_, _06527_);
  and (_03905_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03906_, _03905_, _11817_);
  or (_03908_, _03906_, _03904_);
  and (_04065_, _03908_, _06071_);
  nor (_04070_, _11823_, rst);
  and (_03909_, _11840_, _11810_);
  or (_03910_, _13349_, _13340_);
  or (_03911_, _03910_, _03909_);
  or (_03912_, _03911_, _13346_);
  or (_03913_, _12535_, _11868_);
  or (_03914_, _03913_, _03644_);
  or (_03915_, _11909_, _11811_);
  or (_03916_, _03915_, _11738_);
  or (_03917_, _03916_, _03914_);
  or (_03918_, _13353_, _03894_);
  and (_03920_, _11397_, _08749_);
  or (_03921_, _03920_, _03918_);
  or (_03922_, _03921_, _03917_);
  or (_03923_, _13335_, _11812_);
  or (_03925_, _03923_, _13355_);
  or (_03926_, _03925_, _03892_);
  or (_03927_, _11833_, _11806_);
  or (_03928_, _11880_, _11853_);
  or (_03930_, _03928_, _03927_);
  or (_03931_, _03930_, _03926_);
  or (_03932_, _03931_, _03922_);
  or (_03933_, _03932_, _03912_);
  and (_03934_, _03933_, _06527_);
  and (_03935_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03937_, _13641_, _11744_);
  or (_03938_, _13385_, _03937_);
  or (_03939_, _03938_, _03935_);
  or (_03940_, _03939_, _03934_);
  and (_04077_, _03940_, _06071_);
  or (_03941_, _13924_, rst);
  nor (_04086_, _03941_, _13919_);
  and (_04089_, _00427_, _06071_);
  or (_03942_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  nand (_03943_, _06530_, _10989_);
  and (_03944_, _03943_, _06071_);
  and (_04094_, _03944_, _03942_);
  nor (_04107_, _00294_, rst);
  and (_03945_, _11867_, _11422_);
  or (_03946_, _03723_, _13629_);
  or (_03947_, _03946_, _03945_);
  or (_03948_, _03947_, _03722_);
  or (_03949_, _03948_, _03926_);
  and (_03950_, _11391_, _08748_);
  or (_03951_, _03950_, _11909_);
  or (_03952_, _03951_, _11738_);
  or (_03953_, _13627_, _12533_);
  and (_03954_, _11412_, _08750_);
  and (_03955_, _11736_, _11810_);
  or (_03956_, _03955_, _03954_);
  or (_03957_, _03956_, _03953_);
  or (_03958_, _03957_, _03952_);
  or (_03959_, _03918_, _13625_);
  or (_03960_, _03959_, _03958_);
  or (_03961_, _03960_, _03912_);
  or (_03962_, _03961_, _03949_);
  and (_03963_, _03962_, _06527_);
  and (_03964_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03965_, _03964_, _03938_);
  or (_03966_, _03965_, _03963_);
  and (_04111_, _03966_, _06071_);
  and (_03967_, _13822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03969_, _13825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03970_, _03969_, _03967_);
  and (_03971_, _13830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_03972_, _13833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_03973_, _03972_, _03971_);
  or (_03974_, _03973_, _03970_);
  and (_03975_, _13840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03976_, _13844_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_03977_, _03976_, _03975_);
  and (_03978_, _13854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03979_, _13852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03980_, _03979_, _03978_);
  or (_03981_, _03980_, _03977_);
  or (_03982_, _03981_, _03974_);
  and (_03983_, _13860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03984_, _13863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03985_, _03984_, _03983_);
  and (_03986_, _13865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_03987_, _13866_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_03988_, _03987_, _03986_);
  or (_03989_, _03988_, _03985_);
  and (_03990_, _13876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03991_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03992_, _03991_, _03990_);
  and (_03993_, _13870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03994_, _13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03995_, _03994_, _03993_);
  or (_03996_, _03995_, _03992_);
  or (_03997_, _03996_, _03989_);
  or (_03998_, _03997_, _03982_);
  and (_03999_, _13899_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_04000_, _13897_, _12076_);
  or (_04001_, _04000_, _03999_);
  and (_04002_, _13893_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_04003_, _13895_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_04004_, _04003_, _04002_);
  or (_04005_, _04004_, _04001_);
  or (_04007_, _13983_, p2_in[7]);
  or (_04008_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_04009_, _04008_, _04007_);
  and (_04010_, _04009_, _13991_);
  or (_04011_, _13983_, p3_in[7]);
  or (_04012_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_04013_, _04012_, _04011_);
  and (_04014_, _04013_, _13966_);
  or (_04015_, _04014_, _04010_);
  or (_04016_, _13983_, p0_in[7]);
  or (_04017_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_04018_, _04017_, _04016_);
  and (_04019_, _04018_, _14000_);
  or (_04020_, _13983_, p1_in[7]);
  or (_04021_, _00064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_04022_, _04021_, _04020_);
  and (_04023_, _04022_, _14007_);
  or (_04024_, _04023_, _04019_);
  or (_04025_, _04024_, _04015_);
  or (_04026_, _04025_, _04005_);
  and (_04027_, _13889_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04028_, _13885_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_04029_, _04028_, _04027_);
  or (_04030_, _04029_, _04026_);
  or (_04031_, _04030_, _03998_);
  and (_04032_, _04031_, _13919_);
  and (_04033_, _13922_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_04034_, _04033_, _04032_);
  or (_04035_, _04034_, _13924_);
  or (_04036_, _13925_, _07819_);
  and (_04037_, _04036_, _06071_);
  and (_04114_, _04037_, _04035_);
  not (_04038_, _08774_);
  and (_04039_, _04038_, _08771_);
  or (_04041_, _08776_, _08761_);
  or (_04122_, _04041_, _04039_);
  or (_04042_, _08535_, _05768_);
  or (_04043_, _06526_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_04044_, _04043_, _06071_);
  and (_04144_, _04044_, _04042_);
  and (_04045_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_04046_, _12274_, _11735_);
  or (_04047_, _04046_, _03690_);
  and (_04048_, _11410_, _08756_);
  or (_04049_, _04048_, _12549_);
  or (_04051_, _04049_, _11841_);
  or (_04052_, _04051_, _12269_);
  or (_04053_, _04052_, _12532_);
  or (_04055_, _04053_, _04047_);
  and (_04057_, _04055_, _08775_);
  or (_04146_, _04057_, _04045_);
  or (_04058_, _03538_, _11908_);
  or (_04059_, _04058_, _03732_);
  or (_04060_, _12535_, _11803_);
  or (_04061_, _04060_, _04059_);
  and (_04062_, _04061_, _06527_);
  and (_04063_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04064_, _04063_, _04062_);
  or (_04066_, _04064_, _13642_);
  and (_04154_, _04066_, _06071_);
  and (_04067_, _12524_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_04068_, _03694_, _12548_);
  or (_04069_, _04068_, _12547_);
  or (_04071_, _03883_, _11912_);
  or (_04072_, _04071_, _04069_);
  or (_04073_, _04072_, _04060_);
  or (_04074_, _04073_, _03890_);
  and (_04075_, _04074_, _08775_);
  or (_04157_, _04075_, _04067_);
  and (_04076_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_04078_, _13639_, _11412_);
  and (_04079_, _04078_, _06527_);
  or (_04080_, _04079_, _04076_);
  or (_04081_, _04080_, _13642_);
  and (_04159_, _04081_, _06071_);
  or (_04083_, _13628_, _12532_);
  and (_04084_, _04083_, _11421_);
  or (_04085_, _04084_, _13385_);
  or (_04087_, _13638_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04088_, _04087_, _04085_);
  or (_04090_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05686_);
  and (_04091_, _04090_, _06071_);
  and (_04164_, _04091_, _04088_);
  and (_04092_, _12524_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_04093_, _03538_, _11859_);
  or (_04095_, _04093_, _03536_);
  or (_04096_, _04048_, _03537_);
  or (_04097_, _04096_, _03525_);
  or (_04098_, _11876_, _11839_);
  or (_04099_, _04098_, _03506_);
  or (_04100_, _04099_, _04097_);
  or (_04101_, _04100_, _04095_);
  and (_04102_, _04101_, _08775_);
  or (_04166_, _04102_, _04092_);
  and (_04103_, _12524_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  nor (_04104_, _13332_, _11837_);
  nand (_04105_, _04104_, _11846_);
  nor (_04106_, _04105_, _12543_);
  nand (_04108_, _04106_, _13977_);
  or (_04109_, _04108_, _03890_);
  or (_04110_, _13346_, _12528_);
  or (_04112_, _04110_, _03884_);
  or (_04113_, _04112_, _03731_);
  or (_04115_, _04113_, _04109_);
  and (_04116_, _04115_, _08775_);
  or (_04168_, _04116_, _04103_);
  or (_04117_, _06530_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_04118_, _06530_, _05773_);
  and (_04119_, _04118_, _06071_);
  and (_04184_, _04119_, _04117_);
  and (_04120_, _13884_, _12030_);
  or (_04121_, _00303_, _13849_);
  or (_04123_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_04124_, _04123_, _13818_);
  and (_04125_, _04124_, _04121_);
  and (_04126_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_04127_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_04128_, _04127_, _04126_);
  and (_04129_, _04128_, _13849_);
  nor (_04130_, _12426_, _10916_);
  and (_04131_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_04132_, _04131_, _04130_);
  and (_04133_, _04132_, _13828_);
  and (_04134_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_04135_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_04136_, _04135_, _04134_);
  and (_04137_, _04136_, _12426_);
  or (_04138_, _04137_, _04133_);
  or (_04139_, _04138_, _04129_);
  or (_04140_, _04139_, _04125_);
  and (_04141_, _04140_, _04120_);
  and (_04142_, _13847_, _12030_);
  and (_04143_, _13874_, _12030_);
  nor (_04145_, _04143_, _04142_);
  and (_04147_, _13887_, _12030_);
  and (_04148_, _04147_, _13816_);
  or (_04149_, _13838_, _13819_);
  and (_04150_, _04149_, _13837_);
  nor (_04151_, _04150_, _04148_);
  and (_04152_, _04151_, _04145_);
  not (_04153_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_04155_, _04120_, _04153_);
  and (_04156_, _13817_, _13819_);
  and (_04158_, _04147_, _13883_);
  nor (_04160_, _04158_, _04156_);
  and (_04161_, _04160_, _04155_);
  and (_04162_, _04161_, _04152_);
  and (_04163_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_04165_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_04167_, _04165_, _04163_);
  and (_04169_, _04167_, _13842_);
  or (_04170_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_04171_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_04172_, _04171_, _13831_);
  and (_04173_, _04172_, _04170_);
  nor (_04174_, _12426_, _01916_);
  and (_04175_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_04176_, _04175_, _04174_);
  and (_04177_, _04176_, _13818_);
  nand (_04178_, _12426_, _06056_);
  or (_04179_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04180_, _04179_, _13828_);
  and (_04181_, _04180_, _04178_);
  or (_04182_, _04181_, _04177_);
  or (_04183_, _04182_, _04173_);
  or (_04185_, _04183_, _04169_);
  and (_04187_, _04185_, _04156_);
  or (_04188_, _04187_, _04162_);
  and (_04189_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_04190_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_04191_, _04190_, _04189_);
  and (_04192_, _04191_, _13849_);
  nor (_04193_, _12426_, _01786_);
  and (_04195_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_04196_, _04195_, _04193_);
  and (_04198_, _04196_, _13818_);
  nor (_04200_, _12426_, _01815_);
  and (_04202_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_04203_, _04202_, _04200_);
  and (_04204_, _04203_, _13831_);
  or (_04205_, _04204_, _04198_);
  and (_04206_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_04207_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_04208_, _04207_, _04206_);
  and (_04209_, _04208_, _12426_);
  or (_04210_, _04209_, _04205_);
  or (_04211_, _04210_, _04192_);
  and (_04212_, _04211_, _04158_);
  and (_04213_, _00070_, _13831_);
  and (_04214_, _00229_, _13818_);
  or (_04215_, _04214_, _04213_);
  and (_04216_, _04215_, _12426_);
  or (_04217_, _00005_, _13849_);
  or (_04219_, _04022_, _12426_);
  and (_04220_, _04219_, _13842_);
  and (_04221_, _04220_, _04217_);
  or (_04222_, _00139_, _13849_);
  or (_04223_, _03362_, _12426_);
  and (_04224_, _04223_, _13828_);
  and (_04225_, _04224_, _04222_);
  or (_04226_, _04225_, _04221_);
  and (_04227_, _03473_, _13831_);
  and (_04228_, _03612_, _13818_);
  or (_04229_, _04228_, _04227_);
  and (_04230_, _04229_, _13849_);
  or (_04232_, _04230_, _04226_);
  or (_04233_, _04232_, _04216_);
  and (_04234_, _04233_, _04143_);
  or (_04235_, _04234_, _04212_);
  and (_04236_, _12432_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_04237_, _13839_, _12030_);
  and (_04238_, _03366_, _13828_);
  and (_04239_, _03608_, _13818_);
  or (_04240_, _04239_, _04238_);
  and (_04241_, _04240_, _13849_);
  and (_04242_, _00135_, _13828_);
  and (_04243_, _00224_, _13818_);
  or (_04244_, _04243_, _04242_);
  and (_04245_, _04244_, _12426_);
  or (_04246_, _14005_, _13849_);
  or (_04247_, _04018_, _12426_);
  and (_04248_, _04247_, _13842_);
  and (_04250_, _04248_, _04246_);
  or (_04251_, _00066_, _13849_);
  or (_04252_, _03468_, _12426_);
  and (_04253_, _04252_, _13831_);
  and (_04254_, _04253_, _04251_);
  or (_04255_, _04254_, _04250_);
  or (_04256_, _04255_, _04245_);
  or (_04257_, _04256_, _04241_);
  and (_04258_, _04257_, _04237_);
  or (_04259_, _04258_, _04236_);
  or (_04260_, _04259_, _04235_);
  or (_04261_, _04260_, _04188_);
  and (_04262_, _13988_, _13842_);
  and (_04263_, _00218_, _13818_);
  or (_04264_, _04263_, _04262_);
  and (_04265_, _00148_, _13828_);
  and (_04266_, _00075_, _13831_);
  or (_04267_, _04266_, _04265_);
  or (_04268_, _04267_, _04264_);
  and (_04269_, _04268_, _13846_);
  and (_04270_, _00144_, _13828_);
  and (_04271_, _00079_, _13831_);
  or (_04272_, _04271_, _04270_);
  and (_04273_, _13997_, _13842_);
  and (_04274_, _00213_, _13818_);
  or (_04275_, _04274_, _04273_);
  or (_04276_, _04275_, _04272_);
  and (_04277_, _04276_, _12221_);
  or (_04278_, _04277_, _04269_);
  and (_04279_, _04278_, _12426_);
  and (_04280_, _04009_, _13842_);
  and (_04281_, _03623_, _13818_);
  or (_04282_, _04281_, _04280_);
  and (_04283_, _03375_, _13828_);
  and (_04284_, _03459_, _13831_);
  or (_04285_, _04284_, _04283_);
  or (_04286_, _04285_, _04282_);
  and (_04287_, _04286_, _12221_);
  and (_04288_, _04013_, _13842_);
  and (_04289_, _03619_, _13818_);
  or (_04290_, _04289_, _04288_);
  and (_04291_, _03371_, _13828_);
  and (_04292_, _03463_, _13831_);
  or (_04293_, _04292_, _04291_);
  or (_04294_, _04293_, _04290_);
  and (_04295_, _04294_, _13846_);
  or (_04296_, _04295_, _04287_);
  and (_04297_, _04296_, _13849_);
  or (_04298_, _04297_, _04279_);
  and (_04299_, _04298_, _04142_);
  nor (_04300_, _12426_, _01030_);
  and (_04301_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_04302_, _04301_, _04300_);
  and (_04303_, _04302_, _13818_);
  or (_04304_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_04305_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_04306_, _04305_, _13828_);
  and (_04307_, _04306_, _04304_);
  or (_04308_, _04307_, _04303_);
  nor (_04309_, _12426_, _00764_);
  and (_04310_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_04311_, _04310_, _04309_);
  and (_04312_, _04311_, _13831_);
  or (_04313_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_04314_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_04315_, _04314_, _13842_);
  and (_04316_, _04315_, _04313_);
  or (_04317_, _04316_, _04312_);
  or (_04318_, _04317_, _04308_);
  and (_04319_, _04318_, _13839_);
  nor (_04320_, _12426_, _06464_);
  and (_04321_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_04322_, _04321_, _04320_);
  and (_04323_, _04322_, _13818_);
  or (_04324_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_04325_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_04326_, _04325_, _13828_);
  and (_04327_, _04326_, _04324_);
  or (_04328_, _04327_, _04323_);
  and (_04329_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04330_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_04331_, _04330_, _04329_);
  and (_04332_, _04331_, _13831_);
  or (_04333_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_04334_, _13849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04335_, _04334_, _13842_);
  and (_04336_, _04335_, _04333_);
  or (_04337_, _04336_, _04332_);
  or (_04338_, _04337_, _04328_);
  and (_04339_, _04338_, _13853_);
  or (_04340_, _04339_, _04319_);
  and (_04341_, _04340_, _13819_);
  and (_04342_, _13848_, _13819_);
  nand (_04343_, _12426_, _06495_);
  or (_04344_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_04345_, _04344_, _13828_);
  and (_04346_, _04345_, _04343_);
  nand (_04347_, _12426_, _06489_);
  or (_04348_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_04349_, _04348_, _13818_);
  and (_04350_, _04349_, _04347_);
  or (_04351_, _04350_, _04346_);
  or (_04352_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand (_04353_, _12426_, _06492_);
  and (_04354_, _04353_, _13831_);
  and (_04356_, _04354_, _04352_);
  or (_04357_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_04358_, _12426_, _06482_);
  and (_04359_, _04358_, _13842_);
  and (_04360_, _04359_, _04357_);
  or (_04362_, _04360_, _04356_);
  or (_04363_, _04362_, _04351_);
  and (_04364_, _04363_, _04342_);
  and (_04365_, _13874_, _13819_);
  nor (_04366_, _12426_, _13703_);
  and (_04367_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_04369_, _04367_, _04366_);
  and (_04370_, _04369_, _13828_);
  nand (_04372_, _12426_, _07907_);
  or (_04374_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_04375_, _04374_, _13818_);
  and (_04376_, _04375_, _04372_);
  or (_04377_, _04376_, _04370_);
  or (_04378_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand (_04379_, _12426_, _13746_);
  and (_04380_, _04379_, _13842_);
  and (_04381_, _04380_, _04378_);
  or (_04382_, _12426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand (_04383_, _12426_, _00435_);
  and (_04384_, _04383_, _13831_);
  and (_04385_, _04384_, _04382_);
  or (_04386_, _04385_, _04381_);
  or (_04387_, _04386_, _04377_);
  and (_04388_, _04387_, _04365_);
  and (_04389_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_04390_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_04391_, _04390_, _04389_);
  and (_04392_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04393_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_04394_, _04393_, _04392_);
  or (_04395_, _04394_, _04391_);
  and (_04396_, _04395_, _13849_);
  and (_04397_, _13842_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_04398_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_04399_, _04398_, _04397_);
  and (_04400_, _13831_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_04401_, _13828_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_04402_, _04401_, _04400_);
  or (_04403_, _04402_, _04399_);
  and (_04404_, _04403_, _12426_);
  or (_04405_, _04404_, _04396_);
  and (_04406_, _04405_, _04148_);
  or (_04407_, _04406_, _04388_);
  or (_04408_, _04407_, _04364_);
  or (_04409_, _04408_, _04341_);
  or (_04410_, _04409_, _04299_);
  or (_04411_, _04410_, _04261_);
  or (_04412_, _04411_, _04141_);
  and (_04413_, _04148_, _07766_);
  nor (_04414_, _04413_, _12231_);
  nand (_04415_, _04236_, _06803_);
  and (_04416_, _04415_, _04414_);
  and (_04417_, _04416_, _04412_);
  and (_04418_, _13842_, _06360_);
  and (_04419_, _13831_, _12120_);
  or (_04420_, _04419_, _04418_);
  and (_04421_, _04420_, _13849_);
  and (_04422_, _13842_, _12019_);
  and (_04423_, _13831_, _06435_);
  or (_04424_, _04423_, _04422_);
  and (_04425_, _04424_, _12426_);
  nor (_04426_, _12426_, _06609_);
  and (_04427_, _12426_, _11023_);
  or (_04428_, _04427_, _04426_);
  and (_04429_, _04428_, _13828_);
  nor (_04430_, _12426_, _06993_);
  and (_04431_, _12426_, _07978_);
  or (_04432_, _04431_, _04430_);
  and (_04433_, _04432_, _13818_);
  or (_04434_, _04433_, _04429_);
  or (_04435_, _04434_, _04425_);
  nor (_04436_, _04435_, _04421_);
  nor (_04438_, _04436_, _04414_);
  or (_04439_, _04438_, _04417_);
  and (_04186_, _04439_, _06071_);
  nor (_04440_, _00426_, rst);
  or (_04441_, _00425_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_04442_, _00425_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_04443_, _04442_, _04441_);
  and (_04194_, _04443_, _04440_);
  or (_04444_, _03703_, _13340_);
  and (_04445_, _04444_, _06527_);
  nand (_04446_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_04447_, _04446_, _11819_);
  or (_04448_, _04447_, _04445_);
  and (_04197_, _04448_, _06071_);
  and (_04449_, _11889_, _13378_);
  or (_04450_, _04449_, _03950_);
  or (_04451_, _04450_, _11917_);
  or (_04452_, _04451_, _03883_);
  or (_04453_, _04452_, _04058_);
  or (_04454_, _03658_, _13976_);
  or (_04455_, _04454_, _13630_);
  or (_04456_, _04455_, _04453_);
  or (_04457_, _04456_, _03655_);
  and (_04458_, _04457_, _06527_);
  and (_04459_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04460_, _04459_, _03664_);
  or (_04461_, _04460_, _04458_);
  and (_04201_, _04461_, _06071_);
  or (_04463_, _04093_, _03883_);
  or (_04465_, _04463_, _03898_);
  or (_04466_, _13337_, _11868_);
  or (_04467_, _13633_, _03876_);
  or (_04468_, _04467_, _04466_);
  or (_04469_, _03526_, _13345_);
  or (_04470_, _04469_, _04468_);
  or (_04471_, _11869_, _11837_);
  or (_04472_, _03888_, _04471_);
  or (_04473_, _04472_, _04470_);
  or (_04474_, _04473_, _04465_);
  and (_04475_, _04474_, _06527_);
  and (_04476_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04478_, _04476_, _11818_);
  or (_04479_, _04478_, _04475_);
  and (_04218_, _04479_, _06071_);
  or (_04481_, _07108_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_04482_, _03792_, rst);
  and (_04231_, _04482_, _04481_);
  nand (_04483_, _07759_, _07715_);
  or (_04484_, _07759_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_04485_, _04484_, _06071_);
  and (_04249_, _04485_, _04483_);
  nand (_04486_, _08988_, _06359_);
  and (_04487_, _04486_, _06071_);
  and (_04488_, _02646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_04489_, _04488_, _02647_);
  nand (_04490_, _04489_, _09028_);
  nor (_04491_, _12295_, _06803_);
  and (_04492_, _12295_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_04493_, _04492_, _04491_);
  or (_04494_, _04493_, _09028_);
  and (_04495_, _04494_, _04490_);
  or (_04496_, _04495_, _08988_);
  and (_04355_, _04496_, _04487_);
  nor (_04497_, _13738_, _13778_);
  and (_04498_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_04499_, _04498_, _04497_);
  and (_04500_, _04499_, _13798_);
  nand (_04501_, _07885_, _06359_);
  nand (_04502_, _09341_, _07902_);
  and (_04503_, _04502_, _02727_);
  and (_04504_, _04503_, _04501_);
  or (_04361_, _04504_, _04500_);
  and (_04505_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_04506_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_04507_, _04506_, _04505_);
  or (_04508_, _04507_, _13744_);
  and (_04509_, _04508_, _06071_);
  nand (_04510_, _13759_, _06359_);
  and (_04368_, _04510_, _04509_);
  and (_04511_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_04513_, pc_log_change, _04512_);
  or (_04514_, _04513_, _04511_);
  and (_04371_, _04514_, _06071_);
  nand (_04515_, _13723_, _07977_);
  or (_04516_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_04517_, _04516_, _06071_);
  and (_04373_, _04517_, _04515_);
  not (_04518_, _06054_);
  and (_04519_, _06059_, _04518_);
  and (_04520_, _04519_, _06036_);
  not (_04521_, _04520_);
  or (_04522_, _04521_, _06053_);
  or (_04523_, _04520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_04524_, _04523_, _06071_);
  and (_04437_, _04524_, _04522_);
  and (_04525_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_04526_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_04527_, _04526_, _04525_);
  and (_04528_, _04527_, _13798_);
  nand (_04529_, _09037_, _07885_);
  nand (_04530_, _07977_, _07902_);
  and (_04531_, _04530_, _02727_);
  and (_04532_, _04531_, _04529_);
  or (_04462_, _04532_, _04528_);
  and (_04533_, _13759_, _11023_);
  and (_04534_, _13740_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_04535_, _13738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_04536_, _04535_, _04534_);
  nor (_04537_, _04536_, _13744_);
  and (_04538_, _13753_, _06435_);
  or (_04539_, _04538_, _04537_);
  or (_04540_, _04539_, _04533_);
  and (_04464_, _04540_, _06071_);
  nand (_04541_, _13723_, _06609_);
  or (_04542_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_04543_, _04542_, _06071_);
  and (_04477_, _04543_, _04541_);
  nand (_04544_, _13723_, _06993_);
  or (_04545_, _13723_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_04546_, _04545_, _06071_);
  and (_04480_, _04546_, _04544_);
  and (_04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04548_, _04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04549_, _04548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_04550_, _04549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04551_, _04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_04552_, _04551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04553_, _04552_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04554_, _04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04555_, _04554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04556_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04557_, _04556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_04558_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04559_, _04558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04560_, _04558_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04561_, _04560_, _04559_);
  and (_04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04563_, _04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04564_, _04562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04565_, _04564_, _04563_);
  and (_04566_, _02453_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04567_, _04566_);
  nor (_04568_, _04563_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04569_, _04563_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04570_, _04569_, _04568_);
  nor (_04571_, _04570_, _08210_);
  and (_04572_, _04570_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04573_, _04572_, _04571_);
  or (_04574_, _04573_, _04567_);
  nor (_04575_, _04570_, _08176_);
  and (_04576_, _04570_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_04577_, _04576_, _04575_);
  nor (_04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04579_, _04578_);
  or (_04580_, _04579_, _04577_);
  and (_04581_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01884_);
  not (_04582_, _04581_);
  nor (_04583_, _04570_, _08240_);
  and (_04584_, _04570_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04585_, _04584_, _04583_);
  or (_04586_, _04585_, _04582_);
  and (_04587_, _04586_, _04580_);
  and (_04588_, _04587_, _04574_);
  or (_04589_, _04588_, _04565_);
  not (_04590_, _04563_);
  not (_04591_, _04570_);
  and (_04592_, _04591_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04593_, _04570_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04594_, _04593_, _04592_);
  or (_04595_, _04594_, _04590_);
  not (_04596_, _04565_);
  and (_04597_, _04570_, _08228_);
  or (_04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  nand (_04599_, _04598_, _04581_);
  or (_04600_, _04599_, _04597_);
  and (_04601_, _04570_, _08233_);
  or (_04602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_04603_, _04602_, _04562_);
  or (_04604_, _04603_, _04601_);
  and (_04605_, _04604_, _04600_);
  and (_04606_, _04570_, _08215_);
  or (_04607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nand (_04608_, _04607_, _04578_);
  or (_04609_, _04608_, _04606_);
  and (_04610_, _04570_, _08203_);
  or (_04611_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_04612_, _04611_, _04566_);
  or (_04613_, _04612_, _04610_);
  and (_04614_, _04613_, _04609_);
  and (_04615_, _04614_, _04605_);
  or (_04616_, _04615_, _04596_);
  and (_04617_, _04616_, _04595_);
  and (_04618_, _04617_, _04589_);
  and (_04619_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04620_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_04621_, _04620_, _04619_);
  and (_04622_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04623_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04624_, _04623_, _04622_);
  and (_04625_, _04624_, _04621_);
  and (_04626_, _04625_, _04596_);
  and (_04627_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04628_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04629_, _04628_, _04627_);
  and (_04630_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04631_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04632_, _04631_, _04630_);
  and (_04633_, _04632_, _04629_);
  and (_04634_, _04633_, _04565_);
  or (_04635_, _04634_, _04591_);
  nor (_04636_, _04635_, _04626_);
  and (_04637_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04638_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_04639_, _04638_, _04637_);
  and (_04640_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_04641_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04642_, _04641_, _04640_);
  and (_04643_, _04642_, _04639_);
  nor (_04644_, _04643_, _04565_);
  and (_04645_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04646_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04647_, _04646_, _04645_);
  and (_04648_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04649_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04650_, _04649_, _04648_);
  and (_04651_, _04650_, _04647_);
  nor (_04652_, _04651_, _04596_);
  or (_04653_, _04652_, _04644_);
  and (_04654_, _04653_, _04591_);
  nor (_04655_, _04654_, _04636_);
  nor (_04656_, _04655_, _04618_);
  nor (_04657_, _04556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04658_, _04657_, _04557_);
  and (_04659_, _04658_, _04656_);
  and (_04660_, _04659_, _02142_);
  nor (_04661_, _04557_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04662_, _04661_, _04558_);
  and (_04663_, _04662_, _04656_);
  nor (_04664_, _04662_, _04656_);
  nor (_04665_, _04664_, _04663_);
  nor (_04666_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04667_, _04666_, _04556_);
  and (_04668_, _04667_, _04656_);
  nor (_04669_, _04554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_04670_, _04669_, _04555_);
  and (_04671_, _04670_, _04656_);
  nor (_04672_, _04667_, _04656_);
  nor (_04673_, _04672_, _04668_);
  nor (_04674_, _04670_, _04656_);
  nor (_04675_, _04674_, _04671_);
  not (_04676_, _04675_);
  nor (_04677_, _04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_04678_, _04677_, _04554_);
  and (_04679_, _04678_, _04656_);
  nor (_04680_, _04552_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_04681_, _04680_, _04553_);
  and (_04682_, _04681_, _04656_);
  nor (_04683_, _04678_, _04656_);
  nor (_04684_, _04683_, _04679_);
  nor (_04685_, _04551_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_04686_, _04685_, _04552_);
  and (_04687_, _04686_, _04656_);
  nor (_04688_, _04686_, _04656_);
  and (_04689_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04690_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_04691_, _04690_, _04689_);
  and (_04692_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_04693_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04694_, _04693_, _04692_);
  and (_04695_, _04694_, _04691_);
  nor (_04696_, _04695_, _04565_);
  and (_04697_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04698_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04699_, _04698_, _04697_);
  and (_04700_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04701_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04702_, _04701_, _04700_);
  and (_04703_, _04702_, _04699_);
  nor (_04704_, _04703_, _04596_);
  or (_04705_, _04704_, _04696_);
  and (_04706_, _04705_, _04570_);
  and (_04707_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04708_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_04709_, _04708_, _04707_);
  and (_04710_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_04711_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04712_, _04711_, _04710_);
  and (_04713_, _04712_, _04709_);
  nor (_04714_, _04713_, _04565_);
  and (_04715_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04716_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04717_, _04716_, _04715_);
  and (_04718_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04719_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04720_, _04719_, _04718_);
  and (_04721_, _04720_, _04717_);
  nor (_04722_, _04721_, _04596_);
  or (_04723_, _04722_, _04714_);
  and (_04724_, _04723_, _04591_);
  nor (_04725_, _04724_, _04706_);
  nor (_04726_, _04725_, _04618_);
  nor (_04727_, _04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04728_, _04727_, _04551_);
  and (_04729_, _04728_, _04726_);
  nor (_04730_, _04728_, _04726_);
  nor (_04731_, _04730_, _04729_);
  not (_04732_, _04731_);
  and (_04733_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04734_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_04735_, _04734_, _04733_);
  and (_04736_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_04737_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04738_, _04737_, _04736_);
  and (_04739_, _04738_, _04735_);
  and (_04740_, _04739_, _04596_);
  and (_04741_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04742_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04743_, _04742_, _04741_);
  and (_04744_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04745_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04746_, _04745_, _04744_);
  and (_04747_, _04746_, _04743_);
  and (_04748_, _04747_, _04565_);
  or (_04749_, _04748_, _04591_);
  nor (_04750_, _04749_, _04740_);
  and (_04751_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_04752_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_04753_, _04752_, _04751_);
  and (_04754_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04755_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04756_, _04755_, _04754_);
  and (_04757_, _04756_, _04753_);
  nor (_04758_, _04757_, _04565_);
  and (_04759_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04760_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04761_, _04760_, _04759_);
  and (_04762_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04763_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04764_, _04763_, _04762_);
  and (_04765_, _04764_, _04761_);
  nor (_04766_, _04765_, _04596_);
  or (_04767_, _04766_, _04758_);
  and (_04768_, _04767_, _04591_);
  nor (_04769_, _04768_, _04750_);
  nor (_04770_, _04769_, _04618_);
  nor (_04771_, _04549_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_04772_, _04771_, _04550_);
  and (_04773_, _04772_, _04770_);
  nor (_04774_, _04772_, _04770_);
  nor (_04775_, _04774_, _04773_);
  not (_04776_, _04775_);
  and (_04777_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04778_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_04779_, _04778_, _04777_);
  and (_04780_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_04781_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04782_, _04781_, _04780_);
  and (_04783_, _04782_, _04779_);
  and (_04784_, _04783_, _04596_);
  and (_04785_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04786_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_04787_, _04786_, _04785_);
  and (_04788_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_04789_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04790_, _04789_, _04788_);
  and (_04791_, _04790_, _04787_);
  and (_04792_, _04791_, _04565_);
  or (_04793_, _04792_, _04570_);
  nor (_04794_, _04793_, _04784_);
  and (_04795_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04796_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_04797_, _04796_, _04795_);
  and (_04798_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_04799_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04800_, _04799_, _04798_);
  and (_04801_, _04800_, _04797_);
  and (_04802_, _04801_, _04596_);
  and (_04803_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04804_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04805_, _04804_, _04803_);
  and (_04806_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04807_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04808_, _04807_, _04806_);
  and (_04809_, _04808_, _04805_);
  and (_04810_, _04809_, _04565_);
  or (_04811_, _04810_, _04591_);
  nor (_04812_, _04811_, _04802_);
  nor (_04813_, _04812_, _04794_);
  nor (_04814_, _04813_, _04618_);
  nor (_04815_, _04548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04816_, _04815_, _04549_);
  and (_04817_, _04816_, _04814_);
  and (_04818_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04819_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_04820_, _04819_, _04818_);
  and (_04821_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_04822_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04823_, _04822_, _04821_);
  and (_04824_, _04823_, _04820_);
  and (_04825_, _04824_, _04596_);
  and (_04826_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04827_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_04828_, _04827_, _04826_);
  and (_04829_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_04830_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04831_, _04830_, _04829_);
  and (_04832_, _04831_, _04828_);
  and (_04833_, _04832_, _04565_);
  or (_04834_, _04833_, _04591_);
  nor (_04835_, _04834_, _04825_);
  and (_04836_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04837_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_04838_, _04837_, _04836_);
  and (_04839_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_04840_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04841_, _04840_, _04839_);
  and (_04842_, _04841_, _04838_);
  nor (_04843_, _04842_, _04565_);
  and (_04844_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04845_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04846_, _04845_, _04844_);
  and (_04847_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04848_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04849_, _04848_, _04847_);
  and (_04850_, _04849_, _04846_);
  nor (_04851_, _04850_, _04596_);
  or (_04852_, _04851_, _04843_);
  and (_04853_, _04852_, _04591_);
  nor (_04854_, _04853_, _04835_);
  nor (_04855_, _04854_, _04618_);
  nor (_04856_, _04547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04857_, _04856_, _04548_);
  and (_04858_, _04857_, _04855_);
  nor (_04859_, _04857_, _04855_);
  and (_04860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02461_);
  and (_04861_, _01884_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04862_, _04861_, _04860_);
  not (_04863_, _04862_);
  and (_04864_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04865_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_04866_, _04865_, _04864_);
  and (_04867_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_04868_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04869_, _04868_, _04867_);
  and (_04870_, _04869_, _04866_);
  nor (_04871_, _04870_, _04565_);
  and (_04872_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04873_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04874_, _04873_, _04872_);
  and (_04875_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04876_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04877_, _04876_, _04875_);
  and (_04878_, _04877_, _04874_);
  nor (_04879_, _04878_, _04596_);
  or (_04880_, _04879_, _04871_);
  and (_04881_, _04880_, _04570_);
  and (_04882_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04883_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_04884_, _04883_, _04882_);
  and (_04885_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_04886_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04887_, _04886_, _04885_);
  and (_04888_, _04887_, _04884_);
  nor (_04889_, _04888_, _04565_);
  and (_04890_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04891_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_04892_, _04891_, _04890_);
  and (_04893_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04894_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04895_, _04894_, _04893_);
  and (_04896_, _04895_, _04892_);
  nor (_04897_, _04896_, _04596_);
  or (_04898_, _04897_, _04889_);
  and (_04899_, _04898_, _04591_);
  nor (_04900_, _04899_, _04881_);
  nor (_04901_, _04900_, _04618_);
  and (_04902_, _04901_, _04863_);
  and (_04903_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_04904_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_04905_, _04904_, _04903_);
  and (_04906_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_04907_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_04908_, _04907_, _04906_);
  and (_04909_, _04908_, _04905_);
  nor (_04910_, _04909_, _04565_);
  and (_04911_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04912_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_04913_, _04912_, _04911_);
  and (_04914_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04915_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_04916_, _04915_, _04914_);
  and (_04917_, _04916_, _04913_);
  nor (_04918_, _04917_, _04596_);
  or (_04919_, _04918_, _04910_);
  and (_04920_, _04919_, _04591_);
  and (_04921_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04922_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_04923_, _04922_, _04921_);
  and (_04924_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04925_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_04926_, _04925_, _04924_);
  and (_04927_, _04926_, _04923_);
  nor (_04928_, _04927_, _04596_);
  and (_04929_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04930_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_04931_, _04930_, _04929_);
  and (_04932_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_04933_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_04934_, _04933_, _04932_);
  and (_04935_, _04934_, _04931_);
  nor (_04936_, _04935_, _04565_);
  nor (_04937_, _04936_, _04928_);
  nor (_04938_, _04937_, _04591_);
  nor (_04939_, _04938_, _04920_);
  nor (_04940_, _04939_, _04618_);
  and (_04941_, _04940_, _01884_);
  and (_04942_, _04566_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04943_, _04581_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_04944_, _04943_, _04942_);
  and (_04945_, _04578_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_04946_, _04562_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04947_, _04946_, _04945_);
  and (_04948_, _04947_, _04944_);
  and (_04949_, _04948_, _04596_);
  and (_04950_, _04581_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04951_, _04566_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_04952_, _04951_, _04950_);
  and (_04953_, _04578_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_04954_, _04562_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_04955_, _04954_, _04953_);
  and (_04956_, _04955_, _04952_);
  and (_04957_, _04956_, _04565_);
  or (_04958_, _04957_, _04570_);
  nor (_04959_, _04958_, _04949_);
  and (_04960_, _04581_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04961_, _04566_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_04962_, _04961_, _04960_);
  and (_04963_, _04578_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_04964_, _04562_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04965_, _04962_);
  nor (_04967_, _04966_, _04565_);
  and (_04968_, _04566_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04969_, _04562_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04970_, _04969_, _04968_);
  and (_04971_, _04581_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04972_, _04578_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04973_, _04972_, _04971_);
  and (_04974_, _04973_, _04970_);
  nor (_04975_, _04974_, _04596_);
  or (_04976_, _04975_, _04967_);
  and (_04977_, _04976_, _04570_);
  nor (_04978_, _04977_, _04959_);
  nor (_04979_, _04978_, _04618_);
  and (_04980_, _04979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04981_, _04940_, _01884_);
  nor (_04982_, _04981_, _04941_);
  and (_04983_, _04982_, _04980_);
  nor (_04984_, _04983_, _04941_);
  nor (_04985_, _04901_, _04863_);
  nor (_04986_, _04985_, _04902_);
  not (_04987_, _04986_);
  nor (_04988_, _04987_, _04984_);
  nor (_04989_, _04988_, _04902_);
  nor (_04990_, _04989_, _04859_);
  nor (_04991_, _04990_, _04858_);
  nor (_04992_, _04816_, _04814_);
  nor (_04993_, _04992_, _04817_);
  not (_04994_, _04993_);
  nor (_04995_, _04994_, _04991_);
  nor (_04996_, _04995_, _04817_);
  nor (_04997_, _04996_, _04776_);
  nor (_04998_, _04997_, _04773_);
  nor (_04999_, _04998_, _04732_);
  nor (_05000_, _04999_, _04729_);
  nor (_05001_, _05000_, _04688_);
  or (_05002_, _05001_, _04687_);
  nor (_05003_, _04681_, _04656_);
  nor (_05004_, _05003_, _04682_);
  and (_05005_, _05004_, _05002_);
  and (_05006_, _05005_, _04684_);
  or (_05007_, _05006_, _04682_);
  nor (_05008_, _05007_, _04679_);
  nor (_05009_, _05008_, _04676_);
  and (_05010_, _05009_, _04673_);
  or (_05011_, _05010_, _04671_);
  nor (_05012_, _05011_, _04668_);
  nor (_05013_, _04658_, _04656_);
  nor (_05014_, _05013_, _04659_);
  not (_05015_, _05014_);
  nor (_05016_, _05015_, _05012_);
  and (_05017_, _05016_, _04665_);
  or (_05018_, _05017_, _04663_);
  nor (_05019_, _05018_, _04660_);
  and (_05020_, _05019_, _04561_);
  not (_05021_, _05020_);
  not (_05022_, _04656_);
  nor (_05023_, _05019_, _05022_);
  nor (_05024_, _04656_, _04561_);
  nor (_05025_, _05024_, cy_reg);
  not (_05026_, _05025_);
  nor (_05027_, _05026_, _05023_);
  and (_05028_, _05027_, _05021_);
  nor (_05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_05030_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  or (_05031_, _05030_, _05029_);
  nand (_05032_, _05031_, _04559_);
  or (_05033_, _05031_, _04559_);
  and (_05034_, _05033_, _05032_);
  nor (_05035_, _05034_, _05028_);
  not (_05036_, cy_reg);
  nor (_05037_, _04662_, _05036_);
  nor (_05038_, _05016_, _04659_);
  nor (_05039_, _05038_, _04665_);
  and (_05040_, _05038_, _04665_);
  or (_05041_, _05040_, _05039_);
  nor (_05042_, _05041_, cy_reg);
  nor (_05043_, _05042_, _05037_);
  nor (_05044_, _05043_, _02178_);
  and (_05045_, _05034_, _05028_);
  or (_05046_, _05045_, _05044_);
  or (_05047_, _05046_, _05035_);
  and (_05048_, _04561_, cy_reg);
  and (_05049_, _04656_, _04561_);
  nor (_05050_, _05049_, _05024_);
  nor (_05051_, _05050_, _05019_);
  and (_05052_, _05050_, _05019_);
  or (_05053_, _05052_, _05051_);
  and (_05054_, _05053_, _05036_);
  nor (_05055_, _05054_, _05048_);
  and (_05056_, _05055_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_05057_, _05055_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_05058_, _05043_, _02178_);
  nor (_05059_, _04667_, _05036_);
  nor (_05060_, _05009_, _04671_);
  nor (_05061_, _05060_, _04673_);
  and (_05062_, _05060_, _04673_);
  or (_05063_, _05062_, _05061_);
  nor (_05064_, _05063_, cy_reg);
  nor (_05065_, _05064_, _05059_);
  and (_05066_, _05065_, _01872_);
  nor (_05067_, _05065_, _01872_);
  and (_05068_, _04678_, cy_reg);
  nor (_05069_, _05005_, _04682_);
  and (_05070_, _05069_, _04684_);
  nor (_05071_, _05069_, _04684_);
  nor (_05072_, _05071_, _05070_);
  nor (_05073_, _05072_, cy_reg);
  nor (_05074_, _05073_, _05068_);
  nor (_05075_, _05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_05076_, _05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_05077_, _04686_, cy_reg);
  nor (_05078_, _04687_, _04688_);
  and (_05079_, _05078_, _05000_);
  nor (_05080_, _05078_, _05000_);
  or (_05081_, _05080_, _05079_);
  and (_05082_, _05081_, _05036_);
  or (_05083_, _05082_, _05077_);
  and (_05084_, _05083_, _01996_);
  nor (_05085_, _05083_, _01996_);
  and (_05086_, _04998_, _04732_);
  nor (_05087_, _05086_, _04999_);
  nor (_05088_, _05087_, cy_reg);
  nor (_05089_, _04728_, _05036_);
  nor (_05090_, _05089_, _05088_);
  and (_05091_, _05090_, _02437_);
  nor (_05092_, _05090_, _02437_);
  and (_05093_, _04996_, _04776_);
  nor (_05094_, _05093_, _04997_);
  nor (_05095_, _05094_, cy_reg);
  nor (_05096_, _04772_, _05036_);
  nor (_05097_, _05096_, _05095_);
  and (_05098_, _05097_, _02076_);
  nor (_05099_, _05097_, _02076_);
  and (_05100_, _04816_, cy_reg);
  and (_05101_, _04994_, _04991_);
  nor (_05102_, _05101_, _04995_);
  and (_05103_, _05102_, _05036_);
  nor (_05104_, _05103_, _05100_);
  and (_05105_, _05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_05106_, _04857_, cy_reg);
  nor (_05107_, _04859_, _04858_);
  not (_05108_, _05107_);
  nor (_05109_, _05108_, _04989_);
  and (_05110_, _05108_, _04989_);
  nor (_05111_, _05110_, _05109_);
  and (_05112_, _05111_, _05036_);
  nor (_05113_, _05112_, _05106_);
  nor (_05114_, _05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05115_, _05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05116_, _04862_, _05036_);
  and (_05117_, _04987_, _04984_);
  nor (_05118_, _05117_, _04988_);
  and (_05119_, _05118_, _05036_);
  nor (_05120_, _05119_, _05116_);
  nor (_05121_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05122_, _04979_, _05036_);
  nor (_05123_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05124_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05125_, _05124_, _05123_);
  nand (_05126_, _05125_, _05122_);
  or (_05127_, _05125_, _05122_);
  and (_05128_, _05127_, _05126_);
  nor (_05129_, _04982_, _04980_);
  nor (_05130_, _05129_, _04983_);
  nor (_05131_, _05130_, cy_reg);
  and (_05132_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05133_, _05132_, _05131_);
  and (_05134_, _05133_, _02433_);
  nor (_05135_, _05133_, _02433_);
  or (_05136_, _05135_, _05134_);
  or (_05137_, _05136_, _05128_);
  and (_05138_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05139_, _05138_, _05137_);
  or (_05140_, _05139_, _05121_);
  or (_05141_, _05140_, _05115_);
  or (_05142_, _05141_, _05114_);
  nor (_05143_, _05104_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_05144_, _05143_, _05142_);
  or (_05145_, _05144_, _05105_);
  or (_05146_, _05145_, _05099_);
  or (_05147_, _05146_, _05098_);
  or (_05148_, _05147_, _05092_);
  or (_05149_, _05148_, _05091_);
  or (_05150_, _05149_, _05085_);
  or (_05151_, _05150_, _05084_);
  nor (_05152_, _05004_, _05002_);
  nor (_05153_, _05152_, _05005_);
  nor (_05154_, _05153_, cy_reg);
  nor (_05155_, _04681_, _05036_);
  nor (_05156_, _05155_, _05154_);
  nor (_05157_, _05156_, _01876_);
  and (_05158_, _05156_, _01876_);
  or (_05159_, _05158_, _05157_);
  or (_05160_, _05159_, _05151_);
  or (_05161_, _05160_, _05076_);
  or (_05162_, _05161_, _05075_);
  and (_05163_, _04670_, cy_reg);
  and (_05164_, _05008_, _04676_);
  nor (_05165_, _05164_, _05009_);
  and (_05166_, _05165_, _05036_);
  nor (_05167_, _05166_, _05163_);
  and (_05168_, _05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_05169_, _05167_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_05170_, _05169_, _05168_);
  or (_05171_, _05170_, _05162_);
  or (_05172_, _05171_, _05067_);
  or (_05173_, _05172_, _05066_);
  and (_05174_, _04658_, cy_reg);
  and (_05175_, _05015_, _05012_);
  nor (_05176_, _05175_, _05016_);
  and (_05177_, _05176_, _05036_);
  nor (_05178_, _05177_, _05174_);
  and (_05179_, _05178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_05180_, _05178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_05181_, _05180_, _05179_);
  or (_05182_, _05181_, _05173_);
  or (_05183_, _05182_, _05058_);
  or (_05184_, _05183_, _05057_);
  or (_05185_, _05184_, _05056_);
  or (_05186_, _05185_, _05047_);
  and (_05187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05188_, _05187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_05189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_05190_, _05189_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_05191_, _05190_, _05188_);
  not (_05192_, _05191_);
  nor (_05193_, _05188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05194_, _05188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05195_, _05194_, _05193_);
  or (_05196_, _05195_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_05197_, _05195_, _08925_);
  and (_05198_, _05197_, _05196_);
  and (_05199_, _05198_, _05192_);
  or (_05200_, _05195_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_05201_, _05195_, _08203_);
  and (_05202_, _05201_, _05191_);
  and (_05203_, _05202_, _05200_);
  or (_05204_, _05203_, _05199_);
  or (_05205_, _05204_, _02433_);
  or (_05206_, _02000_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05207_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05208_, _05207_, _05187_);
  and (_05209_, _05208_, _05206_);
  and (_05210_, _02429_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05211_, _02000_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05212_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_05213_, _05212_, _05211_);
  and (_05214_, _05213_, _05210_);
  or (_05215_, _05214_, _05209_);
  nor (_05216_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_05217_, _05216_, _02429_);
  nor (_05218_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05219_, _05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05220_, _05219_, _05218_);
  and (_05221_, _05220_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05222_, _05216_, _02429_);
  nor (_05223_, _05222_, _05217_);
  or (_05224_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _08819_);
  nand (_05225_, _05224_, _05223_);
  or (_05226_, _05225_, _05221_);
  and (_05227_, _05226_, _02433_);
  nor (_05228_, _05220_, _08210_);
  and (_05229_, _05220_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05230_, _05229_, _05228_);
  or (_05231_, _05230_, _05223_);
  and (_05232_, _05231_, _05227_);
  or (_05233_, _05232_, _05215_);
  and (_05234_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05235_, _02000_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05236_, _05235_, _05234_);
  and (_05237_, _05236_, _02429_);
  and (_05238_, _02000_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05239_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05240_, _05239_, _05238_);
  and (_05241_, _05240_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05242_, _05241_, _05237_);
  or (_05243_, _05242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05244_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05245_, _02000_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05246_, _05245_, _02429_);
  or (_05247_, _05246_, _05244_);
  or (_05248_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05249_, _02000_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05250_, _05249_, _05248_);
  or (_05251_, _05250_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05252_, _05251_, _05247_);
  or (_05253_, _05252_, _02433_);
  and (_05254_, _05253_, _02004_);
  and (_05255_, _05254_, _05243_);
  and (_05256_, _05210_, _05240_);
  or (_05257_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05258_, _02000_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05259_, _05258_, _05187_);
  and (_05260_, _05259_, _05257_);
  or (_05261_, _05260_, _05256_);
  and (_05262_, _05252_, _02433_);
  or (_05263_, _05262_, _05261_);
  and (_05264_, _05263_, _05255_);
  nor (_05265_, _05195_, _08176_);
  and (_05266_, _05195_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_05267_, _05266_, _05265_);
  and (_05268_, _05267_, _05192_);
  or (_05269_, _05195_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand (_05270_, _05195_, _08215_);
  and (_05271_, _05270_, _05191_);
  and (_05272_, _05271_, _05269_);
  or (_05273_, _05272_, _05268_);
  or (_05274_, _05273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05275_, _05274_, _05264_);
  and (_05276_, _05275_, _05233_);
  and (_05277_, _05276_, _05205_);
  or (_05278_, _02433_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05279_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_05280_, _05279_, _05278_);
  nand (_05281_, _05280_, _05220_);
  or (_05282_, _02433_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05283_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05284_, _05283_, _05282_);
  or (_05285_, _05284_, _05220_);
  and (_05286_, _05285_, _05281_);
  or (_05287_, _05286_, _05223_);
  or (_05288_, _05195_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_05289_, _05195_, _08246_);
  and (_05290_, _05289_, _05192_);
  and (_05291_, _05290_, _05288_);
  nand (_05292_, _05195_, _08233_);
  or (_05293_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05294_, _05293_, _05191_);
  and (_05295_, _05294_, _05292_);
  or (_05296_, _05295_, _02433_);
  or (_05297_, _05296_, _05291_);
  nand (_05298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_05299_, _05298_, _05224_);
  and (_05300_, _05299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05301_, _02000_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05302_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05303_, _05302_, _02429_);
  and (_05304_, _05303_, _05301_);
  or (_05305_, _05304_, _05300_);
  and (_05306_, _05305_, _05189_);
  and (_05307_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02433_);
  or (_05308_, _05213_, _02429_);
  or (_05309_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05310_, _02000_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05311_, _05310_, _05309_);
  or (_05312_, _05311_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05313_, _05312_, _05308_);
  and (_05314_, _05313_, _05307_);
  or (_05315_, _05314_, _05306_);
  and (_05316_, _05305_, _02433_);
  or (_05317_, _05316_, _05215_);
  and (_05318_, _05317_, _05315_);
  and (_05319_, _05318_, _05297_);
  and (_05320_, _05319_, _05287_);
  nand (_05321_, _05195_, _08228_);
  or (_05322_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05323_, _05322_, _05321_);
  or (_05324_, _05323_, _05192_);
  or (_05325_, _05195_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_05326_, _05195_, _08886_);
  and (_05327_, _05326_, _05325_);
  or (_05328_, _05327_, _05191_);
  and (_05329_, _05328_, _05324_);
  or (_05330_, _05329_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05331_, _05220_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_05332_, _05245_, _02433_);
  or (_05333_, _05332_, _05331_);
  and (_05334_, _05220_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05335_, _05238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_05336_, _05335_, _05334_);
  nand (_05337_, _05336_, _05333_);
  nand (_05338_, _05337_, _05223_);
  and (_05339_, _05338_, _05330_);
  and (_05340_, _05339_, _05320_);
  or (_05341_, _05340_, _05277_);
  nor (_05342_, _04578_, _02461_);
  nor (_05343_, _05342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_05344_, _05342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05345_, _05344_, _05343_);
  nand (_05346_, _05345_, _08233_);
  nor (_05347_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05348_, _05347_, _02453_);
  nor (_05349_, _05348_, _05342_);
  and (_05350_, _05349_, _04602_);
  and (_05351_, _05350_, _05346_);
  or (_05352_, _05345_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_05353_, _05349_);
  nand (_05354_, _05345_, _08246_);
  and (_05355_, _05354_, _05353_);
  and (_05356_, _05355_, _05352_);
  or (_05357_, _05356_, _05351_);
  and (_05358_, _05357_, _04581_);
  nand (_05359_, _05345_, _08215_);
  and (_05360_, _05349_, _04607_);
  and (_05361_, _05360_, _05359_);
  and (_05362_, _05345_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05363_, _05345_, _08176_);
  or (_05364_, _05363_, _05362_);
  and (_05365_, _05364_, _05353_);
  or (_05366_, _05365_, _05361_);
  and (_05367_, _05366_, _04566_);
  or (_05368_, _05367_, _05358_);
  nand (_05369_, _05345_, _08228_);
  and (_05370_, _05349_, _04598_);
  and (_05371_, _05370_, _05369_);
  and (_05372_, _05345_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05373_, _05345_, _08240_);
  or (_05374_, _05373_, _05372_);
  and (_05375_, _05374_, _05353_);
  or (_05376_, _05375_, _05371_);
  and (_05377_, _05376_, _04562_);
  nand (_05378_, _05345_, _08203_);
  and (_05379_, _05349_, _04611_);
  and (_05380_, _05379_, _05378_);
  and (_05381_, _05345_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05382_, _05345_, _08210_);
  or (_05383_, _05382_, _05381_);
  and (_05384_, _05383_, _05353_);
  or (_05385_, _05384_, _05380_);
  and (_05386_, _05385_, _04578_);
  or (_05387_, _05386_, _05377_);
  or (_05388_, _05387_, _05368_);
  nor (_05389_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_05390_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_05391_, _05390_, _05389_);
  or (_05392_, _05391_, _04579_);
  nor (_05393_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_05394_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nand (_05395_, _05394_, _05393_);
  nand (_05396_, _05395_, _04562_);
  and (_05397_, _05396_, _05392_);
  nor (_05398_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_05399_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_05400_, _05399_, _05398_);
  nand (_05401_, _05400_, _04566_);
  nor (_05402_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_05403_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_05404_, _05403_, _05402_);
  nand (_05405_, _05404_, _04581_);
  and (_05406_, _05405_, _05401_);
  and (_05407_, _05406_, _05397_);
  nand (_05408_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05409_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05410_, _05409_, _05408_);
  nand (_05411_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nand (_05412_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_05413_, _05412_, _05411_);
  and (_05414_, _05413_, _05410_);
  nand (_05415_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_05416_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_05417_, _05416_, _05415_);
  nand (_05418_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_05419_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_05420_, _05419_, _05418_);
  and (_05421_, _05420_, _05417_);
  and (_05422_, _05421_, _05414_);
  and (_05423_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_05424_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or (_05425_, _05424_, _05423_);
  and (_05426_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_05427_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or (_05428_, _05427_, _05426_);
  or (_05429_, _05428_, _05425_);
  and (_05430_, _04581_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_05431_, _04578_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or (_05432_, _05431_, _05430_);
  and (_05433_, _04562_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_05434_, _04566_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or (_05435_, _05434_, _05433_);
  or (_05436_, _05435_, _05432_);
  and (_05437_, _05436_, _05429_);
  and (_05438_, _05437_, _05422_);
  and (_05439_, _05438_, _05407_);
  or (_05440_, _05439_, _02461_);
  nor (_05441_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_05442_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_05443_, _05442_, _05441_);
  or (_05444_, _05443_, _04579_);
  or (_05445_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand (_05446_, _05445_, _04562_);
  or (_05447_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand (_05448_, _05447_, _04562_);
  and (_05449_, _05448_, _05446_);
  and (_05450_, _05449_, _05444_);
  nor (_05451_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_05452_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand (_05453_, _05452_, _05451_);
  nand (_05454_, _05453_, _04581_);
  nor (_05455_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_05456_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand (_05457_, _05456_, _05455_);
  nand (_05458_, _05457_, _04566_);
  and (_05459_, _05458_, _05454_);
  and (_05460_, _05459_, _05450_);
  nand (_05461_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05462_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05463_, _05462_, _05461_);
  nand (_05464_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_05465_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05466_, _05465_, _05464_);
  and (_05467_, _05466_, _05463_);
  nand (_05468_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nand (_05469_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_05470_, _05469_, _05468_);
  nand (_05471_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nand (_05472_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_05473_, _05472_, _05471_);
  and (_05474_, _05473_, _05470_);
  and (_05475_, _05474_, _05467_);
  and (_05476_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_05477_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or (_05478_, _05477_, _05476_);
  and (_05479_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_05480_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or (_05481_, _05480_, _05479_);
  or (_05482_, _05481_, _05478_);
  and (_05483_, _04562_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_05484_, _04581_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  or (_05485_, _05484_, _05483_);
  and (_05486_, _04566_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_05487_, _04578_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or (_05488_, _05487_, _05486_);
  or (_05489_, _05488_, _05485_);
  and (_05490_, _05489_, _05482_);
  and (_05491_, _05490_, _05475_);
  and (_05492_, _05491_, _05460_);
  or (_05493_, _05492_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05494_, _05493_, _05440_);
  or (_05495_, _05494_, _02457_);
  and (_05496_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_05497_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or (_05498_, _05497_, _05496_);
  and (_05499_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_05500_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or (_05501_, _05500_, _05499_);
  or (_05502_, _05501_, _05498_);
  and (_05503_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_05504_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or (_05505_, _05504_, _05503_);
  and (_05506_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_05507_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or (_05508_, _05507_, _05506_);
  or (_05509_, _05508_, _05505_);
  or (_05510_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_05511_, _05510_, _04578_);
  or (_05512_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_05513_, _05512_, _04562_);
  or (_05514_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_05515_, _05514_, _04581_);
  and (_05516_, _05515_, _05513_);
  and (_05517_, _05516_, _05511_);
  and (_05518_, _05517_, _05509_);
  and (_05519_, _05518_, _05502_);
  or (_05520_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_05521_, _05520_, _04562_);
  and (_05522_, _05521_, _02461_);
  nand (_05523_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or (_05524_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand (_05525_, _05524_, _04566_);
  and (_05526_, _05525_, _05523_);
  nand (_05527_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand (_05528_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_05529_, _05528_, _05527_);
  and (_05530_, _05529_, _05526_);
  and (_05531_, _05530_, _05522_);
  nand (_05532_, _04562_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_05533_, _04566_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05534_, _05533_, _05532_);
  nand (_05535_, _04578_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_05536_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_05537_, _05536_, _05535_);
  and (_05538_, _05537_, _05534_);
  nand (_05539_, _04581_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  or (_05540_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand (_05541_, _05540_, _04566_);
  and (_05542_, _05541_, _05539_);
  or (_05543_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_05544_, _05543_, _04581_);
  or (_05545_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand (_05546_, _05545_, _04578_);
  and (_05547_, _05546_, _05544_);
  and (_05548_, _05547_, _05542_);
  and (_05549_, _05548_, _05538_);
  and (_05550_, _05549_, _05531_);
  and (_05551_, _05550_, _05519_);
  and (_05552_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_05553_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or (_05554_, _05553_, _05552_);
  and (_05555_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_05556_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or (_05557_, _05556_, _05555_);
  or (_05558_, _05557_, _05554_);
  and (_05559_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_05560_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or (_05561_, _05560_, _05559_);
  and (_05562_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_05563_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or (_05564_, _05563_, _05562_);
  or (_05565_, _05564_, _05561_);
  or (_05566_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_05567_, _05566_, _04578_);
  or (_05568_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_05569_, _05568_, _04562_);
  or (_05570_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_05571_, _05570_, _04581_);
  and (_05572_, _05571_, _05569_);
  and (_05573_, _05572_, _05567_);
  and (_05574_, _05573_, _05565_);
  and (_05575_, _05574_, _05558_);
  nand (_05576_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05577_, _05576_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand (_05578_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05579_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05580_, _05579_, _05578_);
  or (_05581_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nand (_05582_, _05581_, _04562_);
  or (_05583_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_05584_, _05583_, _04581_);
  and (_05585_, _05584_, _05582_);
  and (_05586_, _05585_, _05580_);
  and (_05587_, _05586_, _05577_);
  nand (_05588_, _04562_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nand (_05589_, _04566_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_05590_, _05589_, _05588_);
  nand (_05591_, _04578_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  or (_05592_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_05593_, _05592_, _04578_);
  and (_05594_, _05593_, _05591_);
  and (_05595_, _05594_, _05590_);
  nand (_05596_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  or (_05597_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_05598_, _05597_, _04566_);
  and (_05599_, _05598_, _05596_);
  nand (_05600_, _04581_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  or (_05601_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_05602_, _05601_, _04566_);
  and (_05603_, _05602_, _05600_);
  and (_05604_, _05603_, _05599_);
  and (_05605_, _05604_, _05595_);
  and (_05606_, _05605_, _05587_);
  and (_05607_, _05606_, _05575_);
  or (_05608_, _05607_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05609_, _05608_, _05551_);
  or (_05610_, _02457_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05611_, _04611_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05612_, _05611_, _05610_);
  or (_05613_, _02457_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05614_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05615_, _05614_, _02461_);
  and (_05616_, _05615_, _05613_);
  or (_05617_, _05616_, _05612_);
  and (_05618_, _05617_, _01884_);
  or (_05619_, _02457_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_05620_, _05619_, _04607_);
  and (_05621_, _05620_, _04860_);
  or (_05622_, _02457_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05623_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05624_, _05623_, _04547_);
  and (_05625_, _05624_, _05622_);
  or (_05626_, _05625_, _05621_);
  or (_05627_, _05626_, _05618_);
  and (_05628_, _05627_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05629_, _02457_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05630_, _04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05631_, _05630_, _05629_);
  or (_05632_, _02457_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05634_, _05633_, _02461_);
  and (_05635_, _05634_, _05632_);
  or (_05636_, _05635_, _05631_);
  and (_05637_, _05636_, _04578_);
  and (_05638_, _04566_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or (_05639_, _02457_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05640_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05641_, _05640_, _05639_);
  and (_05642_, _05641_, _05638_);
  or (_05643_, _02457_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05644_, _05643_, _04602_);
  and (_05645_, _04860_, _02453_);
  and (_05646_, _05645_, _05644_);
  or (_05647_, _05646_, _05642_);
  or (_05648_, _05647_, _05637_);
  or (_05649_, _05648_, _05628_);
  and (_05650_, _05617_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05651_, _05620_, _04861_);
  or (_05652_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05653_, _02457_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05654_, _05653_, _05652_);
  and (_05655_, _05654_, _05347_);
  or (_05656_, _05655_, _02453_);
  or (_05657_, _05656_, _05651_);
  or (_05658_, _05657_, _05650_);
  and (_05659_, _05636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05660_, _05644_, _04861_);
  and (_05661_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05662_, _02457_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05663_, _05662_, _05661_);
  and (_05664_, _05663_, _05347_);
  or (_05665_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05666_, _05665_, _05660_);
  or (_05667_, _05666_, _05659_);
  nor (_05668_, _02472_, first_instr);
  and (_05669_, _05668_, _05667_);
  and (_05670_, _05669_, _05658_);
  and (_05671_, _05670_, _05649_);
  and (_05672_, _05671_, _05609_);
  nand (_05673_, _05672_, _05495_);
  nor (_05674_, _05673_, _04618_);
  and (_05675_, _05674_, _05388_);
  and (_05676_, _05675_, _05341_);
  and (property_invalid_jnc, _05676_, _05186_);
  or (_05677_, pc_log_change_r, _05036_);
  nand (_05678_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_00000_, _05678_, _05677_);
  and (_05679_, _02472_, first_instr);
  or (_00001_, _05679_, rst);
  dff (cy_reg, _00000_);
  dff (pc_log_change_r, pc_log_change);
  dff (first_instr, _00001_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _10170_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _10174_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _10176_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _10180_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _10184_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _10187_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _10190_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _14025_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _10077_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _10081_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _10086_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _10091_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _10094_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _10099_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _10104_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _10106_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _14024_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _09985_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _09989_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _09994_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _09996_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _10001_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _10005_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _10009_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _09885_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _09889_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _09892_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _09895_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _09898_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _09902_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _09905_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _09907_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _14016_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _14017_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _14018_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _14019_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _14020_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _14021_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _14022_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _14023_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _14008_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _14009_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _14010_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _14011_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _14012_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _14013_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _14014_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _14015_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _14046_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _14047_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _14048_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _14049_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _14050_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _14051_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _14052_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _14053_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _09547_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _09551_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _14040_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _14041_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _14042_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _14043_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _14044_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _14045_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _14032_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _14033_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _14034_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _14035_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _14036_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _14037_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _14038_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _14039_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _09356_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _09360_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _09363_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _09366_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _09371_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _09373_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _09376_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _09379_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _09253_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _09257_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _09261_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _09266_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _09270_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _09274_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _09278_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _09281_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _08846_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _08850_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _08855_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _08860_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _08863_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _08868_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _08872_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _08875_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _08738_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _08743_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _08747_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _08751_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _08755_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _08759_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _08763_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _08766_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _14027_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _09055_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _09058_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _09060_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _09065_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _09069_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _09074_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _09077_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _08960_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _08965_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _08969_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _08972_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _08976_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _14026_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _08981_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _08983_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _09161_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _09164_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _14028_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _14029_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _14030_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _14031_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _09176_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _09179_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _07408_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _07436_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _07476_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _07529_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _07582_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _07640_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _07708_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _07780_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _07842_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _07921_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _07995_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _08055_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _08149_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _08265_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _08385_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _07359_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13520_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11175_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _01851_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _13787_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03880_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _03929_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04231_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _03897_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _00186_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03639_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03585_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03521_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03500_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03499_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _00014_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00359_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07052_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _01317_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _06617_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _06606_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _06604_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _06589_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03450_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _05682_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _01763_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _02490_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _03013_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _03347_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _05974_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _06092_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _06074_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _06060_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _07066_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _07069_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _07072_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _07074_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _07077_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _07080_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _07082_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06950_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _12290_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _12300_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12907_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _02980_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _04070_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _02983_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _07649_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _04122_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _00393_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _04056_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _07568_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _07382_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _03936_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _03756_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _07485_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _03702_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _03565_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _04144_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _04146_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _11599_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04154_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _11499_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _04157_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03742_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _11988_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _04159_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _04111_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _04077_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04164_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03682_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _04166_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03834_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _04065_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _04218_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _04168_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03822_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _04197_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _04201_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _00388_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _00872_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _03330_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _08716_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _06658_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _02255_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03813_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _01442_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _03847_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _02041_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _03317_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _05935_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _02074_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _11489_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _07111_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _03377_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _03924_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _02499_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _13801_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _12048_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00781_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _06811_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _02186_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12624_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _00826_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _13436_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _01189_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _01236_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _07982_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _01914_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _11544_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _09983_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02175_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _06778_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _01902_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _12997_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _03837_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _03823_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _03968_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _11892_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _10178_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _13487_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _12018_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _13371_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _13605_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _11820_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _12012_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _13686_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _09300_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _11767_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _12099_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _03576_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _12101_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _05750_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _08866_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _08890_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _03344_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _09087_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _11072_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _08870_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _08894_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _09193_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _00264_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _01835_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _12917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _12170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _11443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _00531_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _00864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _08157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _01059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _01056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _01152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _01651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _01052_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _01673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _01663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _01045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _01145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _01202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _00725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _01716_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01009_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _01730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _01138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _01734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _01732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _01002_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _01743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _01736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _00999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _01135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _01175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _01199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _04371_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _03907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _03431_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _12214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _11720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _11898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _01247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _07987_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _13610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _11809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _11494_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _11285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _12254_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _12217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _10032_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _08447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _04050_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _12229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _11437_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _02080_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _04094_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _12261_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05683_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _13941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _12281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _11432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03678_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _03652_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _12287_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03481_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _02688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00574_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _01299_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _13110_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _13098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _13085_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _13056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _13034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12334_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _13281_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _13359_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _13328_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _13289_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12327_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _11409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _12526_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _12496_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _12490_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _02545_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _11941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _11832_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _12345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _12293_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _12089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _12220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _12175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _12141_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _12111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _12342_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11291_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _11181_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _11223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _11220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03479_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _11502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _02025_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _04199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _10459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _10449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10430_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12361_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _11034_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _10901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _11033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _12358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11393_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03485_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _11712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _11389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _11692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _11871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _09186_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _01829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _02239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _12367_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _11373_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _01278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _00563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _12179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _02547_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _06953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00728_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _07131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12392_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _03853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03772_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _07589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _07524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _07125_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03483_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _02874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _02792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _02908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _02895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11004_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _03353_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _03351_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _10999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _03358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _03356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _10996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11339_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _03440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _03424_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _10993_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _03579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _03563_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _10991_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _03630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _03587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _10986_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _03713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _03650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _10983_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11184_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _03748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _03715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _01816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _02261_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _02149_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _02274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _10909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11159_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _12694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _02427_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _04089_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _12448_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _12440_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12415_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04194_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _04186_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _04086_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _12265_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _12235_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _12232_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _12226_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03740_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03570_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03614_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04114_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _02537_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _04107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _04054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _07736_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _06199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _00897_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _03554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _00621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _03592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _00641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07260_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _06049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _02104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _06063_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _06052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _06034_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07234_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07238_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _06096_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _02094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _04249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _06130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _02099_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _09235_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _01461_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _13581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _13565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _13573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _13568_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _02794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _13601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _13596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _02506_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _13517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _01890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _00503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _13536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _13542_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _00316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _13478_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _13475_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _02813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _02810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _00433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _00430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08858_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _00475_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _13441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _02825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _10482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _13841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _13834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _02737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _13868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _13862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _13859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _13855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10480_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _02741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _02551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _13775_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _13773_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _13768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _02752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _13795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _00470_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _03285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _03159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _03289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _03287_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _05680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _03153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _03296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _03122_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _03745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _03261_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03246_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _03119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _03862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _03298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _03264_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _03305_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _03303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03867_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _08610_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _04355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _03671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _14001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _13965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _13995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _13992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _13989_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _13984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _00321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _01067_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _01078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _13388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _13392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _13369_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _13366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _13363_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _13374_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _13336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _01071_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _13413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _13433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13497_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _01075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _01073_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _01024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13439_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13464_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13461_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13508_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13502_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13505_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _01028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13571_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _01026_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _01049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13615_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13612_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _01039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _04082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _00258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _01624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _01618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _01616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _01580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _01575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _01572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _03919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _01520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _01501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _01517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _01515_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _01512_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _01505_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _01464_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _03780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _04437_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01367_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _01328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _01359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _01348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _01292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _01275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _01289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _01224_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _01196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _01191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _01157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _01154_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _01149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _05877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _01086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _01083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _01042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _01036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _01019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _01015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _01013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _02561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _07629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07472_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07522_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07513_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07510_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _06783_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _06379_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _06679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _06346_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _12554_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12396_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _01408_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _08216_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _08226_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _03444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _09148_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _10877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _03725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _02197_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _02466_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _02555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _06909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _02765_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02673_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _03057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _12211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _12373_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _12206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04462_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04464_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _12203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _12331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _12471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _12560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04361_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04368_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _12200_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _04373_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _12193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _12315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _12468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _04480_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _04477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _12190_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _12181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _12303_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _12461_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _12557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _12600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _02398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _02400_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02786_);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
